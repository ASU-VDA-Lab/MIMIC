module fake_netlist_6_3036_n_1782 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1782);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1782;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_127),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_30),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_21),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_62),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_35),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_51),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_149),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_25),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_53),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_19),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_110),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_97),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_69),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_119),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_77),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_31),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_157),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_26),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_39),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_40),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_115),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_14),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_86),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_13),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_0),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_31),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_57),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_99),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_128),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_105),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_76),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_121),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_83),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_1),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_67),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_85),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_50),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_154),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_29),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_98),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_44),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_89),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_55),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_146),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_21),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_88),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_159),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_161),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_148),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_92),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_66),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_3),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_3),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_96),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_151),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_15),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_7),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_114),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_112),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_109),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_116),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_91),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_45),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_170),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_7),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_165),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_52),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_14),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_5),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_124),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_137),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_108),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_64),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_52),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_11),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_73),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_35),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_81),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_17),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_37),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_74),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_33),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_6),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_102),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_164),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_145),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_103),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_141),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_68),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_61),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_156),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_90),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_29),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_155),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_41),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_24),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_123),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_54),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_129),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_33),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_142),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_169),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_126),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_168),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_56),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_44),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_166),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_65),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_134),
.Y(n_297)
);

HB1xp67_ASAP7_75t_SL g298 ( 
.A(n_48),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_133),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_41),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_143),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_160),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_8),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_117),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_27),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_9),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_106),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_46),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_13),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_60),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_152),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_30),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_135),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_153),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_51),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_43),
.Y(n_317)
);

BUFx10_ASAP7_75t_L g318 ( 
.A(n_132),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_70),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_4),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_144),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_34),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_36),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_24),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_59),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_28),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_100),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_136),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_9),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_147),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_101),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_45),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_15),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_80),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_140),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_16),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_47),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_78),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_11),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_5),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_167),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_95),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_203),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_207),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_192),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_192),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_192),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_208),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_298),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_192),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_192),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_175),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_221),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_221),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_211),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_196),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_214),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_225),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_229),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_230),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_297),
.B(n_2),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_232),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_342),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_R g365 ( 
.A(n_215),
.B(n_163),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_221),
.Y(n_366)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_177),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_172),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_221),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_174),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_233),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_172),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_253),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_234),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_253),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_199),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_253),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_212),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_290),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_253),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_253),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_183),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_238),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_191),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_193),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_202),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_226),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_242),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_247),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_219),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_206),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_263),
.B(n_2),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_269),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_258),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_250),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_281),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_254),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_255),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_340),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_256),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_R g403 ( 
.A(n_257),
.B(n_158),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_282),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_L g405 ( 
.A(n_180),
.B(n_6),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_260),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_294),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_262),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_174),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_309),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_R g411 ( 
.A(n_265),
.B(n_277),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_312),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_317),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_278),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_173),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_280),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_246),
.B(n_8),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_286),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_R g421 ( 
.A(n_289),
.B(n_104),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_295),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_299),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_209),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_301),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_182),
.B(n_10),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_339),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_302),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_424),
.B(n_209),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_344),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_345),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_348),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_355),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_359),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_347),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_347),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_370),
.B(n_204),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_350),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_351),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_353),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_360),
.B(n_210),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_353),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_354),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_354),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_400),
.B(n_307),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_356),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_352),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_366),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_361),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_369),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_363),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_369),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_373),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_357),
.B(n_376),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_371),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_377),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_377),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_374),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_349),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_R g472 ( 
.A(n_406),
.B(n_310),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_380),
.B(n_248),
.Y(n_473)
);

OA21x2_ASAP7_75t_L g474 ( 
.A1(n_426),
.A2(n_227),
.B(n_182),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_381),
.B(n_248),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_343),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_393),
.B(n_252),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_395),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_385),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_382),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_390),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_397),
.B(n_291),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_358),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_382),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_399),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_402),
.B(n_231),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_386),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_414),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_387),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_388),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_417),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_420),
.B(n_291),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_423),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_388),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_425),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_396),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_428),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_438),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_442),
.A2(n_362),
.B1(n_364),
.B2(n_419),
.Y(n_507)
);

INVx6_ASAP7_75t_L g508 ( 
.A(n_437),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_434),
.B(n_435),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_447),
.B(n_411),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_442),
.B(n_409),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_492),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_489),
.B(n_365),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_487),
.B(n_368),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

INVx4_ASAP7_75t_L g518 ( 
.A(n_440),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_494),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_445),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_471),
.A2(n_422),
.B1(n_408),
.B2(n_392),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_398),
.Y(n_522)
);

AND3x4_ASAP7_75t_L g523 ( 
.A(n_437),
.B(n_405),
.C(n_379),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_394),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_270),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_452),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_473),
.B(n_227),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_455),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_436),
.B(n_372),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_487),
.B(n_372),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_487),
.B(n_416),
.Y(n_532)
);

INVx6_ASAP7_75t_L g533 ( 
.A(n_473),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_473),
.B(n_276),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_473),
.B(n_288),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_457),
.B(n_383),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_440),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_475),
.B(n_311),
.Y(n_538)
);

NAND2xp33_ASAP7_75t_SL g539 ( 
.A(n_429),
.B(n_204),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_475),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_476),
.A2(n_267),
.B1(n_394),
.B2(n_279),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_494),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_475),
.B(n_237),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_477),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_477),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_475),
.B(n_237),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_432),
.B(n_268),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_431),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_499),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

BUFx4f_ASAP7_75t_L g552 ( 
.A(n_474),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_482),
.B(n_268),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_474),
.A2(n_315),
.B1(n_304),
.B2(n_292),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_482),
.B(n_292),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_482),
.B(n_205),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_474),
.A2(n_315),
.B1(n_304),
.B2(n_341),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_474),
.A2(n_341),
.B1(n_367),
.B2(n_272),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_433),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_448),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_448),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_456),
.Y(n_567)
);

INVx4_ASAP7_75t_SL g568 ( 
.A(n_431),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_440),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_482),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_485),
.A2(n_224),
.B1(n_285),
.B2(n_287),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_487),
.B(n_391),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_482),
.B(n_205),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_439),
.B(n_188),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_456),
.Y(n_576)
);

INVx4_ASAP7_75t_SL g577 ( 
.A(n_431),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_482),
.B(n_205),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_500),
.B(n_205),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_503),
.B(n_401),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_431),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_500),
.B(n_205),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_500),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_464),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_500),
.B(n_272),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_464),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_490),
.B(n_427),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_L g588 ( 
.A(n_500),
.B(n_272),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_472),
.B(n_272),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_490),
.B(n_427),
.Y(n_590)
);

AND2x2_ASAP7_75t_SL g591 ( 
.A(n_491),
.B(n_272),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_491),
.B(n_418),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_456),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_495),
.A2(n_410),
.B1(n_415),
.B2(n_413),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_441),
.Y(n_595)
);

CKINVDCx6p67_ASAP7_75t_R g596 ( 
.A(n_430),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_443),
.B(n_213),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_443),
.B(n_218),
.Y(n_598)
);

AND2x2_ASAP7_75t_SL g599 ( 
.A(n_480),
.B(n_223),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_463),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_480),
.B(n_391),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_444),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_480),
.A2(n_415),
.B1(n_413),
.B2(n_412),
.Y(n_603)
);

BUFx4f_ASAP7_75t_L g604 ( 
.A(n_463),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_444),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_446),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_463),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_463),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_430),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_449),
.B(n_404),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_463),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_449),
.B(n_241),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_467),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_459),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_467),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_451),
.B(n_404),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_451),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_466),
.B(n_469),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_467),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_453),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_481),
.B(n_378),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_453),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_454),
.B(n_243),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_479),
.B(n_407),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_454),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_458),
.B(n_245),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_483),
.B(n_271),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_458),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_467),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_488),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_460),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_467),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_460),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_461),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_461),
.B(n_407),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_462),
.B(n_273),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_462),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_467),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_478),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_493),
.A2(n_249),
.B1(n_244),
.B2(n_240),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_478),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_465),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_478),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_465),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_468),
.B(n_274),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_468),
.B(n_283),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_479),
.B(n_293),
.Y(n_649)
);

AND2x6_ASAP7_75t_L g650 ( 
.A(n_470),
.B(n_296),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_496),
.B(n_171),
.Y(n_651)
);

O2A1O1Ixp33_ASAP7_75t_L g652 ( 
.A1(n_516),
.A2(n_200),
.B(n_470),
.C(n_412),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_540),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_515),
.B(n_498),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_512),
.B(n_502),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_L g656 ( 
.A1(n_507),
.A2(n_504),
.B1(n_319),
.B2(n_321),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_562),
.B(n_450),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_525),
.B(n_450),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_540),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_651),
.B(n_430),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_526),
.B(n_430),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_531),
.Y(n_662)
);

OAI221xp5_ASAP7_75t_L g663 ( 
.A1(n_603),
.A2(n_325),
.B1(n_331),
.B2(n_410),
.C(n_217),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_531),
.B(n_450),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_587),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_532),
.B(n_478),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_513),
.B(n_479),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_592),
.Y(n_669)
);

O2A1O1Ixp5_ASAP7_75t_L g670 ( 
.A1(n_552),
.A2(n_479),
.B(n_421),
.C(n_403),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_513),
.B(n_266),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_522),
.B(n_171),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_629),
.B(n_178),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_514),
.B(n_178),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_602),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_508),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_552),
.B(n_179),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_552),
.B(n_179),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_580),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_629),
.B(n_184),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_590),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_555),
.B(n_478),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_606),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_561),
.B(n_478),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_526),
.Y(n_685)
);

INVxp67_ASAP7_75t_SL g686 ( 
.A(n_615),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_517),
.B(n_184),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_519),
.B(n_185),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_SL g689 ( 
.A1(n_510),
.A2(n_300),
.B1(n_324),
.B2(n_323),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_542),
.B(n_185),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_548),
.B(n_186),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_580),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_534),
.B(n_186),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_610),
.B(n_220),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_550),
.B(n_187),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_506),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_508),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_590),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_506),
.Y(n_699)
);

BUFx8_ASAP7_75t_L g700 ( 
.A(n_569),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_596),
.B(n_209),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_606),
.Y(n_702)
);

INVx2_ASAP7_75t_SL g703 ( 
.A(n_524),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_554),
.B(n_187),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_591),
.B(n_189),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_557),
.B(n_189),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_524),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_591),
.B(n_190),
.Y(n_708)
);

AO221x1_ASAP7_75t_L g709 ( 
.A1(n_541),
.A2(n_216),
.B1(n_222),
.B2(n_318),
.C(n_332),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_508),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_610),
.B(n_228),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_535),
.B(n_190),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_599),
.A2(n_173),
.B1(n_336),
.B2(n_333),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_533),
.A2(n_538),
.B1(n_524),
.B2(n_599),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_533),
.A2(n_338),
.B1(n_194),
.B2(n_335),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_546),
.B(n_194),
.Y(n_716)
);

BUFx8_ASAP7_75t_L g717 ( 
.A(n_528),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_642),
.B(n_201),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_620),
.B(n_201),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_611),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_573),
.A2(n_176),
.B1(n_336),
.B2(n_181),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_533),
.A2(n_338),
.B1(n_335),
.B2(n_334),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_630),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_524),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_573),
.B(n_314),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_SL g726 ( 
.A(n_596),
.B(n_216),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_536),
.B(n_314),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_630),
.B(n_327),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_644),
.B(n_327),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_544),
.B(n_545),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_644),
.B(n_646),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_560),
.B(n_328),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_612),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_527),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_563),
.B(n_328),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_530),
.B(n_275),
.C(n_235),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_521),
.B(n_236),
.Y(n_737)
);

NOR2xp67_ASAP7_75t_L g738 ( 
.A(n_616),
.B(n_632),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_616),
.B(n_239),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_564),
.B(n_330),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_623),
.Y(n_741)
);

BUFx12f_ASAP7_75t_SL g742 ( 
.A(n_612),
.Y(n_742)
);

NOR2x1p5_ASAP7_75t_L g743 ( 
.A(n_632),
.B(n_176),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_595),
.B(n_330),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_509),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_539),
.A2(n_334),
.B1(n_216),
.B2(n_222),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_618),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_572),
.B(n_303),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_618),
.B(n_305),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_539),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_618),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_637),
.Y(n_753)
);

NOR3xp33_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_284),
.C(n_251),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_528),
.Y(n_755)
);

INVx8_ASAP7_75t_L g756 ( 
.A(n_527),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_607),
.B(n_318),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_619),
.B(n_306),
.Y(n_758)
);

AND2x6_ASAP7_75t_SL g759 ( 
.A(n_586),
.B(n_333),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_527),
.B(n_264),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_622),
.B(n_222),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_624),
.B(n_308),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_627),
.B(n_313),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_633),
.B(n_318),
.Y(n_764)
);

NAND2x1_ASAP7_75t_L g765 ( 
.A(n_527),
.B(n_82),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_637),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_637),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_635),
.B(n_261),
.Y(n_768)
);

NAND2x1_ASAP7_75t_L g769 ( 
.A(n_527),
.B(n_511),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_527),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_636),
.B(n_259),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_509),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_639),
.B(n_332),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_601),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_589),
.B(n_543),
.Y(n_775)
);

INVx1_ASAP7_75t_SL g776 ( 
.A(n_589),
.Y(n_776)
);

BUFx8_ASAP7_75t_L g777 ( 
.A(n_601),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_626),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_543),
.B(n_326),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_626),
.B(n_326),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_571),
.B(n_322),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_594),
.B(n_322),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_571),
.B(n_71),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_523),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_649),
.B(n_320),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_650),
.B(n_320),
.Y(n_786)
);

INVx8_ASAP7_75t_L g787 ( 
.A(n_650),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_520),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_575),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_583),
.B(n_316),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_597),
.B(n_316),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_551),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_598),
.B(n_181),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_614),
.B(n_625),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_628),
.B(n_198),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_638),
.B(n_197),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_649),
.B(n_197),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_565),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_523),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_195),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_650),
.B(n_195),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_648),
.B(n_12),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_566),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_567),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_605),
.B(n_138),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_662),
.A2(n_553),
.B(n_556),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_657),
.A2(n_553),
.B(n_556),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_675),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_655),
.B(n_617),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_664),
.A2(n_576),
.B(n_593),
.Y(n_810)
);

INVx3_ASAP7_75t_L g811 ( 
.A(n_659),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_705),
.A2(n_547),
.B(n_585),
.C(n_578),
.Y(n_812)
);

OAI321xp33_ASAP7_75t_L g813 ( 
.A1(n_656),
.A2(n_578),
.A3(n_585),
.B1(n_574),
.B2(n_582),
.C(n_579),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_672),
.B(n_574),
.C(n_582),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_767),
.B(n_617),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_794),
.B(n_605),
.Y(n_816)
);

CKINVDCx6p67_ASAP7_75t_R g817 ( 
.A(n_784),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_667),
.A2(n_604),
.B(n_505),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_697),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_778),
.B(n_566),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_703),
.B(n_724),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_733),
.B(n_640),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_789),
.B(n_567),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_697),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_655),
.B(n_640),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_766),
.B(n_615),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_774),
.B(n_593),
.Y(n_827)
);

INVxp67_ASAP7_75t_SL g828 ( 
.A(n_659),
.Y(n_828)
);

BUFx4f_ASAP7_75t_L g829 ( 
.A(n_799),
.Y(n_829)
);

AOI21x1_ASAP7_75t_L g830 ( 
.A1(n_731),
.A2(n_579),
.B(n_576),
.Y(n_830)
);

AO21x1_ASAP7_75t_L g831 ( 
.A1(n_677),
.A2(n_588),
.B(n_558),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_673),
.A2(n_511),
.B(n_549),
.C(n_609),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_668),
.B(n_634),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_658),
.A2(n_600),
.B(n_570),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_672),
.B(n_654),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_772),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_744),
.B(n_645),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_766),
.B(n_615),
.Y(n_838)
);

AOI21x1_ASAP7_75t_L g839 ( 
.A1(n_731),
.A2(n_645),
.B(n_577),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_748),
.B(n_577),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_772),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_788),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_673),
.A2(n_511),
.B(n_549),
.C(n_634),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_721),
.A2(n_549),
.B1(n_634),
.B2(n_631),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_741),
.B(n_518),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_727),
.B(n_621),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_788),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_660),
.B(n_518),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_721),
.A2(n_609),
.B1(n_631),
.B2(n_621),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_752),
.B(n_568),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_660),
.B(n_518),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_669),
.B(n_631),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_680),
.A2(n_609),
.B(n_605),
.C(n_621),
.Y(n_853)
);

OAI22xp5_ASAP7_75t_L g854 ( 
.A1(n_680),
.A2(n_613),
.B1(n_559),
.B2(n_581),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_775),
.A2(n_714),
.B(n_756),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_756),
.A2(n_529),
.B(n_643),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_756),
.A2(n_529),
.B(n_643),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_727),
.B(n_613),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_730),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_755),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_686),
.A2(n_537),
.B(n_643),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_SL g862 ( 
.A(n_734),
.B(n_641),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_679),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_677),
.A2(n_650),
.B(n_558),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_676),
.A2(n_581),
.B(n_559),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_693),
.B(n_650),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_678),
.A2(n_652),
.B(n_705),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_753),
.A2(n_650),
.B1(n_641),
.B2(n_581),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_769),
.A2(n_581),
.B(n_559),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_678),
.A2(n_608),
.B(n_577),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_693),
.B(n_568),
.Y(n_871)
);

NAND3xp33_ASAP7_75t_L g872 ( 
.A(n_749),
.B(n_608),
.C(n_16),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_713),
.A2(n_608),
.B1(n_17),
.B2(n_18),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_708),
.A2(n_12),
.B(n_18),
.C(n_20),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_712),
.B(n_568),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_692),
.B(n_20),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_661),
.B(n_568),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_792),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_787),
.A2(n_608),
.B(n_130),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_710),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_787),
.A2(n_608),
.B(n_122),
.Y(n_881)
);

OAI22xp33_ASAP7_75t_L g882 ( 
.A1(n_665),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_718),
.B(n_22),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_685),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_798),
.Y(n_885)
);

CKINVDCx10_ASAP7_75t_R g886 ( 
.A(n_717),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_671),
.B(n_23),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_783),
.A2(n_111),
.B(n_107),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_776),
.B(n_94),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_783),
.A2(n_93),
.B(n_87),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_666),
.B(n_84),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_760),
.A2(n_75),
.B(n_72),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_694),
.Y(n_893)
);

AND2x4_ASAP7_75t_L g894 ( 
.A(n_710),
.B(n_58),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_681),
.B(n_28),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_683),
.A2(n_32),
.B(n_34),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_702),
.A2(n_32),
.B(n_36),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_698),
.B(n_702),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_700),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_720),
.B(n_42),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_798),
.Y(n_901)
);

AOI33xp33_ASAP7_75t_L g902 ( 
.A1(n_689),
.A2(n_46),
.A3(n_48),
.B1(n_49),
.B2(n_50),
.B3(n_54),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_723),
.A2(n_49),
.B(n_55),
.Y(n_903)
);

BUFx4f_ASAP7_75t_L g904 ( 
.A(n_674),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_708),
.A2(n_725),
.B(n_670),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_781),
.A2(n_790),
.B(n_805),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_653),
.A2(n_699),
.B(n_696),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_804),
.A2(n_734),
.B(n_803),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_795),
.B(n_780),
.Y(n_909)
);

BUFx8_ASAP7_75t_L g910 ( 
.A(n_784),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_739),
.B(n_711),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_712),
.B(n_791),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_734),
.A2(n_716),
.B(n_725),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_791),
.B(n_800),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_758),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_763),
.Y(n_916)
);

O2A1O1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_802),
.A2(n_716),
.B(n_728),
.C(n_729),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_771),
.A2(n_706),
.B(n_732),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_687),
.A2(n_704),
.B(n_735),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_796),
.B(n_800),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_796),
.B(n_719),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_765),
.Y(n_922)
);

AO21x1_ASAP7_75t_L g923 ( 
.A1(n_802),
.A2(n_749),
.B(n_718),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_779),
.A2(n_768),
.B(n_773),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_688),
.A2(n_690),
.B(n_691),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_701),
.B(n_726),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_742),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_768),
.A2(n_729),
.B(n_728),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_674),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_750),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_695),
.A2(n_740),
.B(n_801),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_751),
.A2(n_762),
.B1(n_736),
.B2(n_745),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_762),
.A2(n_745),
.B(n_786),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_782),
.B(n_793),
.Y(n_934)
);

BUFx3_ASAP7_75t_L g935 ( 
.A(n_777),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_785),
.A2(n_797),
.B(n_663),
.Y(n_936)
);

AO21x1_ASAP7_75t_L g937 ( 
.A1(n_797),
.A2(n_785),
.B(n_764),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_713),
.A2(n_707),
.B1(n_747),
.B2(n_722),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_770),
.A2(n_757),
.B(n_761),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_757),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_761),
.A2(n_764),
.B(n_737),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_715),
.A2(n_743),
.B1(n_754),
.B2(n_709),
.Y(n_942)
);

INVx4_ASAP7_75t_L g943 ( 
.A(n_770),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_770),
.A2(n_777),
.B(n_700),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_759),
.B(n_717),
.Y(n_945)
);

BUFx2_ASAP7_75t_L g946 ( 
.A(n_770),
.Y(n_946)
);

NAND2x1p5_ASAP7_75t_L g947 ( 
.A(n_770),
.B(n_734),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_948)
);

OAI21xp33_ASAP7_75t_L g949 ( 
.A1(n_727),
.A2(n_672),
.B(n_713),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_655),
.B(n_741),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_794),
.B(n_662),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_746),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_675),
.Y(n_956)
);

BUFx12f_ASAP7_75t_L g957 ( 
.A(n_700),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_662),
.A2(n_562),
.B1(n_555),
.B2(n_561),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_669),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_794),
.B(n_662),
.Y(n_961)
);

AO21x1_ASAP7_75t_L g962 ( 
.A1(n_677),
.A2(n_678),
.B(n_672),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_662),
.A2(n_552),
.B(n_657),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_746),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_655),
.B(n_741),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_669),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_682),
.A2(n_684),
.B(n_667),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_738),
.B(n_703),
.Y(n_969)
);

AO31x2_ASAP7_75t_L g970 ( 
.A1(n_962),
.A2(n_923),
.A3(n_831),
.B(n_853),
.Y(n_970)
);

AO31x2_ASAP7_75t_L g971 ( 
.A1(n_832),
.A2(n_843),
.A3(n_937),
.B(n_958),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_929),
.B(n_821),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_953),
.B(n_961),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_949),
.A2(n_920),
.B(n_914),
.C(n_912),
.Y(n_974)
);

BUFx2_ASAP7_75t_L g975 ( 
.A(n_860),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_835),
.B(n_912),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_951),
.A2(n_959),
.B(n_955),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_952),
.B(n_966),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_859),
.B(n_915),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_916),
.B(n_909),
.Y(n_980)
);

OAI21x1_ASAP7_75t_SL g981 ( 
.A1(n_939),
.A2(n_913),
.B(n_890),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_862),
.B(n_840),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_963),
.A2(n_968),
.B(n_964),
.Y(n_983)
);

BUFx8_ASAP7_75t_L g984 ( 
.A(n_957),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_943),
.A2(n_958),
.B(n_855),
.Y(n_985)
);

AOI21x1_ASAP7_75t_L g986 ( 
.A1(n_871),
.A2(n_875),
.B(n_858),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_883),
.A2(n_844),
.A3(n_849),
.B(n_854),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_918),
.B(n_816),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_863),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_873),
.A2(n_932),
.B1(n_936),
.B2(n_933),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_906),
.A2(n_866),
.B(n_857),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_934),
.B(n_911),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_887),
.B(n_893),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_819),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_929),
.B(n_821),
.Y(n_995)
);

AO31x2_ASAP7_75t_L g996 ( 
.A1(n_844),
.A2(n_849),
.A3(n_854),
.B(n_846),
.Y(n_996)
);

AND3x2_ASAP7_75t_L g997 ( 
.A(n_899),
.B(n_945),
.C(n_936),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_819),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_921),
.A2(n_851),
.B(n_848),
.C(n_933),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_930),
.B(n_960),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_SL g1001 ( 
.A1(n_947),
.A2(n_963),
.B(n_864),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_905),
.A2(n_867),
.B(n_870),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_917),
.A2(n_928),
.B(n_867),
.C(n_924),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_919),
.B(n_809),
.Y(n_1004)
);

AO31x2_ASAP7_75t_L g1005 ( 
.A1(n_900),
.A2(n_873),
.A3(n_818),
.B(n_825),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_967),
.B(n_940),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_898),
.B(n_823),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_905),
.A2(n_807),
.B(n_806),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_810),
.A2(n_834),
.B(n_869),
.Y(n_1009)
);

AOI221xp5_ASAP7_75t_SL g1010 ( 
.A1(n_938),
.A2(n_895),
.B1(n_882),
.B2(n_942),
.C(n_928),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_898),
.B(n_823),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_924),
.B(n_820),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_856),
.A2(n_931),
.B(n_833),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_884),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_812),
.A2(n_891),
.B(n_925),
.C(n_904),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_908),
.A2(n_807),
.B(n_861),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_865),
.A2(n_806),
.B(n_907),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_820),
.B(n_827),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_947),
.A2(n_864),
.B(n_870),
.Y(n_1019)
);

OA21x2_ASAP7_75t_L g1020 ( 
.A1(n_814),
.A2(n_813),
.B(n_891),
.Y(n_1020)
);

AOI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_938),
.A2(n_874),
.B(n_895),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_946),
.A2(n_828),
.B(n_838),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_826),
.A2(n_811),
.B(n_845),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_900),
.A2(n_956),
.B(n_872),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_840),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_SL g1026 ( 
.A1(n_888),
.A2(n_941),
.B(n_892),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_811),
.B(n_885),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_815),
.A2(n_837),
.B(n_822),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_836),
.B(n_847),
.Y(n_1029)
);

AO21x1_ASAP7_75t_L g1030 ( 
.A1(n_889),
.A2(n_877),
.B(n_942),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_815),
.A2(n_837),
.B(n_822),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_841),
.B(n_954),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_868),
.A2(n_922),
.B(n_904),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_850),
.Y(n_1034)
);

OAI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_842),
.A2(n_878),
.B(n_965),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_901),
.A2(n_879),
.B(n_881),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_922),
.A2(n_850),
.B(n_894),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_852),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_819),
.B(n_824),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_824),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_894),
.B(n_824),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_880),
.B(n_902),
.Y(n_1042)
);

NOR2x1_ASAP7_75t_SL g1043 ( 
.A(n_969),
.B(n_922),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_876),
.B(n_817),
.Y(n_1044)
);

OA21x2_ASAP7_75t_L g1045 ( 
.A1(n_896),
.A2(n_903),
.B(n_897),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_927),
.A2(n_926),
.B(n_880),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_829),
.A2(n_969),
.B(n_935),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_969),
.A2(n_829),
.A3(n_880),
.B(n_910),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_910),
.A2(n_839),
.B(n_830),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_886),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_859),
.B(n_730),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_952),
.B(n_966),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_948),
.A2(n_951),
.B(n_950),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_949),
.A2(n_914),
.B(n_920),
.C(n_912),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_963),
.A2(n_950),
.B(n_948),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_819),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_L g1057 ( 
.A1(n_923),
.A2(n_920),
.B(n_914),
.C(n_912),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_943),
.A2(n_552),
.B(n_756),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_943),
.A2(n_552),
.B(n_756),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_860),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_934),
.B(n_909),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_808),
.Y(n_1062)
);

O2A1O1Ixp5_ASAP7_75t_L g1063 ( 
.A1(n_923),
.A2(n_920),
.B(n_914),
.C(n_912),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_949),
.A2(n_920),
.B1(n_914),
.B2(n_912),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_949),
.A2(n_966),
.B1(n_952),
.B2(n_914),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_SL g1066 ( 
.A1(n_939),
.A2(n_937),
.B(n_913),
.Y(n_1066)
);

AOI221xp5_ASAP7_75t_SL g1067 ( 
.A1(n_949),
.A2(n_883),
.B1(n_873),
.B2(n_656),
.C(n_914),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_949),
.A2(n_914),
.B(n_920),
.C(n_912),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_943),
.A2(n_552),
.B(n_756),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_819),
.Y(n_1070)
);

BUFx2_ASAP7_75t_SL g1071 ( 
.A(n_935),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_963),
.A2(n_950),
.B(n_948),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_952),
.B(n_966),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_840),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_963),
.A2(n_950),
.B(n_948),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_934),
.B(n_909),
.Y(n_1076)
);

NAND3xp33_ASAP7_75t_L g1077 ( 
.A(n_949),
.B(n_920),
.C(n_914),
.Y(n_1077)
);

NAND2x1_ASAP7_75t_L g1078 ( 
.A(n_862),
.B(n_943),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_943),
.A2(n_552),
.B(n_756),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_953),
.B(n_961),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_884),
.B(n_610),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_953),
.B(n_961),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_808),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_953),
.B(n_961),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_859),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_SL g1086 ( 
.A1(n_939),
.A2(n_937),
.B(n_913),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_948),
.A2(n_951),
.B(n_950),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_949),
.A2(n_914),
.B(n_920),
.C(n_912),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_948),
.A2(n_951),
.B(n_950),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_952),
.B(n_966),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_963),
.A2(n_950),
.B(n_948),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_962),
.A2(n_923),
.A3(n_831),
.B(n_853),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_920),
.B1(n_914),
.B2(n_912),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_934),
.B(n_909),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_960),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_808),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_934),
.B(n_909),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_957),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_840),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_953),
.B(n_961),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_943),
.A2(n_552),
.B(n_756),
.Y(n_1101)
);

AND2x2_ASAP7_75t_SL g1102 ( 
.A(n_883),
.B(n_660),
.Y(n_1102)
);

NOR2x1_ASAP7_75t_L g1103 ( 
.A(n_926),
.B(n_738),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_953),
.B(n_961),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_840),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_950),
.B(n_948),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_953),
.B(n_961),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_808),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1065),
.A2(n_976),
.B1(n_1102),
.B2(n_1090),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_SL g1110 ( 
.A(n_990),
.B(n_1052),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_976),
.B(n_973),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1039),
.B(n_972),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_973),
.B(n_1080),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1004),
.A2(n_1053),
.B(n_977),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_975),
.Y(n_1115)
);

OR2x6_ASAP7_75t_L g1116 ( 
.A(n_1071),
.B(n_1037),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_992),
.A2(n_979),
.B1(n_1107),
.B2(n_1082),
.Y(n_1117)
);

OR2x6_ASAP7_75t_SL g1118 ( 
.A(n_1051),
.B(n_1041),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_1060),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1039),
.B(n_972),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_1061),
.B(n_1076),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_995),
.B(n_1041),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1094),
.B(n_1097),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_1085),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_989),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_998),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1074),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1080),
.B(n_1082),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_995),
.B(n_1043),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_1074),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_980),
.B(n_978),
.Y(n_1131)
);

BUFx4f_ASAP7_75t_L g1132 ( 
.A(n_1098),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1087),
.A2(n_1089),
.B(n_988),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1062),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_978),
.A2(n_1084),
.B1(n_1107),
.B2(n_1100),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_1074),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1087),
.A2(n_1089),
.B(n_1106),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_1095),
.Y(n_1138)
);

BUFx6f_ASAP7_75t_L g1139 ( 
.A(n_998),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1084),
.B(n_1100),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_990),
.A2(n_1003),
.B(n_1057),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1014),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1074),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1083),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1104),
.B(n_1064),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1013),
.A2(n_1072),
.B(n_1106),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_998),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1077),
.A2(n_1064),
.B1(n_1093),
.B2(n_1021),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1093),
.A2(n_1021),
.B1(n_1073),
.B2(n_1104),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_993),
.B(n_1000),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_974),
.B(n_1054),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1048),
.B(n_1047),
.Y(n_1152)
);

INVx1_ASAP7_75t_SL g1153 ( 
.A(n_980),
.Y(n_1153)
);

INVx3_ASAP7_75t_SL g1154 ( 
.A(n_1040),
.Y(n_1154)
);

AOI21xp33_ASAP7_75t_L g1155 ( 
.A1(n_1067),
.A2(n_1010),
.B(n_1063),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_984),
.Y(n_1156)
);

O2A1O1Ixp5_ASAP7_75t_SL g1157 ( 
.A1(n_983),
.A2(n_1091),
.B(n_1055),
.C(n_1075),
.Y(n_1157)
);

BUFx12f_ASAP7_75t_L g1158 ( 
.A(n_984),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_983),
.A2(n_1055),
.B(n_1072),
.Y(n_1159)
);

OR2x6_ASAP7_75t_L g1160 ( 
.A(n_1047),
.B(n_1033),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1028),
.B(n_1031),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1068),
.A2(n_1088),
.B(n_999),
.C(n_1024),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1096),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_1015),
.A2(n_1012),
.B(n_1011),
.C(n_1007),
.Y(n_1164)
);

OR2x2_ASAP7_75t_SL g1165 ( 
.A(n_1050),
.B(n_1042),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1038),
.B(n_1042),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1108),
.Y(n_1167)
);

OAI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1081),
.A2(n_1007),
.B1(n_1011),
.B2(n_1018),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1030),
.A2(n_1006),
.B1(n_1103),
.B2(n_1044),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1029),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1018),
.B(n_1012),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1029),
.B(n_1032),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1032),
.B(n_987),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_982),
.A2(n_1001),
.B1(n_1008),
.B2(n_1078),
.Y(n_1174)
);

BUFx12f_ASAP7_75t_L g1175 ( 
.A(n_1040),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1056),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1056),
.B(n_1070),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_987),
.B(n_1027),
.Y(n_1178)
);

BUFx4f_ASAP7_75t_SL g1179 ( 
.A(n_1070),
.Y(n_1179)
);

AO21x2_ASAP7_75t_L g1180 ( 
.A1(n_1075),
.A2(n_1091),
.B(n_1066),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1048),
.B(n_1070),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_994),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1048),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1025),
.Y(n_1184)
);

INVxp67_ASAP7_75t_SL g1185 ( 
.A(n_982),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1105),
.B(n_1034),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_1099),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1099),
.B(n_1105),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_985),
.A2(n_1008),
.B(n_1026),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1046),
.B(n_1049),
.Y(n_1190)
);

AND2x6_ASAP7_75t_L g1191 ( 
.A(n_970),
.B(n_1092),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_997),
.B(n_1024),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_987),
.B(n_996),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1035),
.B(n_970),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1035),
.B(n_970),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_996),
.B(n_1005),
.Y(n_1196)
);

AND2x4_ASAP7_75t_L g1197 ( 
.A(n_1036),
.B(n_1022),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1086),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1020),
.A2(n_1023),
.B1(n_1045),
.B2(n_1101),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1092),
.B(n_1005),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_981),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_1002),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_L g1203 ( 
.A1(n_1020),
.A2(n_1002),
.B(n_1079),
.C(n_1069),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1092),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1019),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_971),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1017),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_971),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_996),
.B(n_986),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1016),
.Y(n_1210)
);

INVx2_ASAP7_75t_SL g1211 ( 
.A(n_1009),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1058),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1059),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1039),
.B(n_972),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1004),
.A2(n_988),
.B(n_943),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_976),
.B(n_973),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1051),
.B(n_730),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_979),
.B(n_738),
.Y(n_1218)
);

AOI222xp33_ASAP7_75t_L g1219 ( 
.A1(n_1052),
.A2(n_949),
.B1(n_1090),
.B2(n_1102),
.C1(n_920),
.C2(n_914),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1004),
.A2(n_988),
.B(n_943),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_998),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1074),
.B(n_1039),
.Y(n_1222)
);

INVx3_ASAP7_75t_L g1223 ( 
.A(n_1074),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1004),
.A2(n_988),
.B(n_943),
.Y(n_1224)
);

AND2x6_ASAP7_75t_L g1225 ( 
.A(n_1025),
.B(n_1034),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1102),
.A2(n_949),
.B1(n_923),
.B2(n_883),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1004),
.A2(n_991),
.B(n_977),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1039),
.B(n_972),
.Y(n_1228)
);

AO32x1_ASAP7_75t_L g1229 ( 
.A1(n_990),
.A2(n_873),
.A3(n_1093),
.B1(n_1064),
.B2(n_656),
.Y(n_1229)
);

BUFx3_ASAP7_75t_L g1230 ( 
.A(n_975),
.Y(n_1230)
);

CKINVDCx14_ASAP7_75t_R g1231 ( 
.A(n_1050),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1065),
.A2(n_976),
.B1(n_1102),
.B2(n_1090),
.Y(n_1232)
);

BUFx2_ASAP7_75t_SL g1233 ( 
.A(n_1014),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_976),
.B(n_973),
.Y(n_1234)
);

INVx5_ASAP7_75t_L g1235 ( 
.A(n_998),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1085),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_998),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_998),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1061),
.B(n_1076),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1004),
.A2(n_991),
.B(n_977),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1071),
.B(n_944),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1004),
.A2(n_991),
.B(n_977),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1085),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1051),
.B(n_730),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1039),
.B(n_972),
.Y(n_1245)
);

OAI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1110),
.A2(n_1117),
.B1(n_1113),
.B2(n_1128),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1122),
.B(n_1129),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1219),
.A2(n_1110),
.B1(n_1109),
.B2(n_1232),
.Y(n_1248)
);

CKINVDCx11_ASAP7_75t_R g1249 ( 
.A(n_1158),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_1231),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1142),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1219),
.A2(n_1226),
.B(n_1109),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1232),
.A2(n_1148),
.B1(n_1149),
.B2(n_1135),
.Y(n_1253)
);

AOI222xp33_ASAP7_75t_L g1254 ( 
.A1(n_1121),
.A2(n_1239),
.B1(n_1123),
.B2(n_1131),
.C1(n_1153),
.C2(n_1135),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1170),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_SL g1256 ( 
.A1(n_1192),
.A2(n_1160),
.B1(n_1233),
.B2(n_1153),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1134),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1235),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1163),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1167),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1145),
.A2(n_1140),
.B1(n_1128),
.B2(n_1113),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1140),
.B(n_1111),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1230),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1166),
.Y(n_1264)
);

BUFx2_ASAP7_75t_R g1265 ( 
.A(n_1156),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1168),
.A2(n_1218),
.B(n_1162),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1184),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1187),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1172),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1179),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1122),
.B(n_1129),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1145),
.A2(n_1151),
.B1(n_1141),
.B2(n_1111),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1172),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1204),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1151),
.A2(n_1141),
.B1(n_1234),
.B2(n_1216),
.Y(n_1275)
);

BUFx2_ASAP7_75t_SL g1276 ( 
.A(n_1115),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1125),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1216),
.A2(n_1234),
.B1(n_1160),
.B2(n_1155),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1225),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1160),
.A2(n_1155),
.B1(n_1159),
.B2(n_1169),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1150),
.B(n_1217),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1225),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1177),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1181),
.Y(n_1284)
);

NAND2x1p5_ASAP7_75t_L g1285 ( 
.A(n_1235),
.B(n_1127),
.Y(n_1285)
);

BUFx4f_ASAP7_75t_SL g1286 ( 
.A(n_1175),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1118),
.A2(n_1244),
.B1(n_1119),
.B2(n_1116),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1235),
.Y(n_1288)
);

BUFx8_ASAP7_75t_L g1289 ( 
.A(n_1138),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1235),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1152),
.A2(n_1202),
.B1(n_1171),
.B2(n_1180),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1171),
.B(n_1124),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1178),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1178),
.Y(n_1294)
);

AOI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1215),
.A2(n_1220),
.B(n_1224),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1227),
.A2(n_1242),
.B(n_1240),
.Y(n_1296)
);

AO21x2_ASAP7_75t_L g1297 ( 
.A1(n_1137),
.A2(n_1114),
.B(n_1133),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_SL g1298 ( 
.A(n_1176),
.Y(n_1298)
);

CKINVDCx11_ASAP7_75t_R g1299 ( 
.A(n_1154),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_1236),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1182),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1152),
.A2(n_1180),
.B1(n_1198),
.B2(n_1243),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1165),
.A2(n_1116),
.B1(n_1183),
.B2(n_1185),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1112),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1112),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1157),
.A2(n_1146),
.B(n_1189),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1225),
.Y(n_1307)
);

CKINVDCx11_ASAP7_75t_R g1308 ( 
.A(n_1139),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1245),
.B(n_1120),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1173),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1214),
.B(n_1245),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1214),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1173),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1228),
.B(n_1186),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1206),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1228),
.B(n_1188),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1208),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1193),
.A2(n_1161),
.B1(n_1191),
.B2(n_1241),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1147),
.Y(n_1319)
);

OAI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1189),
.A2(n_1114),
.B(n_1133),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1222),
.B(n_1139),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1182),
.Y(n_1322)
);

OAI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1196),
.A2(n_1193),
.B(n_1209),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1221),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1242),
.A2(n_1137),
.B(n_1203),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1182),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1130),
.B(n_1136),
.Y(n_1327)
);

BUFx8_ASAP7_75t_L g1328 ( 
.A(n_1221),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_1164),
.B(n_1174),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1237),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1225),
.B(n_1195),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1237),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1191),
.A2(n_1200),
.B1(n_1196),
.B2(n_1194),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1237),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1199),
.A2(n_1213),
.B(n_1197),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1238),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1238),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1222),
.B(n_1238),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1136),
.B(n_1223),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1132),
.Y(n_1340)
);

BUFx12f_ASAP7_75t_L g1341 ( 
.A(n_1126),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_1174),
.A2(n_1132),
.B1(n_1143),
.B2(n_1223),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1210),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1191),
.A2(n_1229),
.B1(n_1197),
.B2(n_1207),
.Y(n_1344)
);

OAI22x1_ASAP7_75t_L g1345 ( 
.A1(n_1190),
.A2(n_1205),
.B1(n_1201),
.B2(n_1229),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1126),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1191),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1229),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1207),
.Y(n_1349)
);

AO21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1201),
.A2(n_1212),
.B(n_1211),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1110),
.A2(n_914),
.B1(n_920),
.B2(n_912),
.Y(n_1351)
);

NAND2x1p5_ASAP7_75t_L g1352 ( 
.A(n_1235),
.B(n_1127),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1144),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1235),
.Y(n_1354)
);

CKINVDCx6p67_ASAP7_75t_R g1355 ( 
.A(n_1158),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1110),
.A2(n_1102),
.B1(n_660),
.B2(n_883),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1219),
.A2(n_949),
.B1(n_1110),
.B2(n_1102),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1122),
.B(n_1129),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1219),
.A2(n_949),
.B1(n_1110),
.B2(n_1102),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1293),
.B(n_1294),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1284),
.B(n_1333),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1277),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1350),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1274),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1262),
.B(n_1292),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1333),
.B(n_1310),
.Y(n_1366)
);

AO21x1_ASAP7_75t_SL g1367 ( 
.A1(n_1248),
.A2(n_1253),
.B(n_1266),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1300),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1264),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1267),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1313),
.B(n_1291),
.Y(n_1371)
);

AO21x2_ASAP7_75t_L g1372 ( 
.A1(n_1320),
.A2(n_1306),
.B(n_1325),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1291),
.B(n_1248),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1325),
.A2(n_1252),
.B(n_1295),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1343),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1323),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1315),
.Y(n_1377)
);

OR2x6_ASAP7_75t_L g1378 ( 
.A(n_1296),
.B(n_1329),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1255),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1278),
.B(n_1343),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1269),
.B(n_1273),
.Y(n_1381)
);

NOR2x1_ASAP7_75t_R g1382 ( 
.A(n_1249),
.B(n_1299),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1349),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1255),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1317),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1329),
.B(n_1347),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1297),
.Y(n_1387)
);

OR2x2_ASAP7_75t_L g1388 ( 
.A(n_1278),
.B(n_1331),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1280),
.B(n_1260),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1260),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1335),
.A2(n_1348),
.B(n_1351),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1303),
.B(n_1345),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1280),
.B(n_1253),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1250),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1318),
.A2(n_1344),
.B(n_1279),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1257),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1259),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1353),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1302),
.B(n_1272),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1344),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1328),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1281),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1246),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1302),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1272),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1275),
.Y(n_1406)
);

BUFx2_ASAP7_75t_L g1407 ( 
.A(n_1342),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1261),
.B(n_1359),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1283),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1282),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1327),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1307),
.A2(n_1275),
.B(n_1261),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1339),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1254),
.B(n_1356),
.Y(n_1414)
);

INVxp33_ASAP7_75t_L g1415 ( 
.A(n_1263),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1287),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1328),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1357),
.B(n_1359),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1357),
.B(n_1316),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1327),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1256),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1316),
.B(n_1247),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1285),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1352),
.A2(n_1314),
.B(n_1346),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1352),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1271),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1364),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1368),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1364),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1365),
.B(n_1358),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1386),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1404),
.B(n_1276),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1402),
.B(n_1362),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1410),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1404),
.B(n_1391),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1386),
.B(n_1321),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1386),
.B(n_1338),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1366),
.B(n_1336),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1366),
.B(n_1324),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1394),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1371),
.B(n_1332),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1371),
.B(n_1337),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1369),
.B(n_1312),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1361),
.B(n_1330),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1375),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1391),
.B(n_1305),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_1415),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1375),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_1378),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1361),
.B(n_1309),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1390),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1370),
.Y(n_1452)
);

NOR4xp25_ASAP7_75t_SL g1453 ( 
.A(n_1407),
.B(n_1403),
.C(n_1421),
.D(n_1376),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1393),
.A2(n_1340),
.B1(n_1268),
.B2(n_1250),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1391),
.B(n_1304),
.Y(n_1455)
);

INVx1_ASAP7_75t_SL g1456 ( 
.A(n_1411),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1379),
.Y(n_1457)
);

BUFx2_ASAP7_75t_SL g1458 ( 
.A(n_1363),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1396),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1403),
.B(n_1289),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1384),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1381),
.B(n_1289),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1409),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1367),
.A2(n_1268),
.B1(n_1355),
.B2(n_1311),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1393),
.B(n_1289),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1391),
.B(n_1251),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1380),
.B(n_1334),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1422),
.B(n_1298),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1380),
.B(n_1334),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1363),
.B(n_1424),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1378),
.B(n_1319),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1378),
.B(n_1319),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1378),
.B(n_1290),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1378),
.B(n_1326),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1414),
.A2(n_1270),
.B1(n_1326),
.B2(n_1258),
.C(n_1301),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1427),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1428),
.B(n_1389),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1431),
.B(n_1392),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1431),
.B(n_1392),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1464),
.A2(n_1407),
.B(n_1373),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1392),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1466),
.B(n_1416),
.C(n_1421),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1463),
.B(n_1389),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1433),
.B(n_1376),
.Y(n_1484)
);

AND2x2_ASAP7_75t_SL g1485 ( 
.A(n_1449),
.B(n_1399),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1452),
.B(n_1441),
.Y(n_1486)
);

NAND3xp33_ASAP7_75t_L g1487 ( 
.A(n_1466),
.B(n_1416),
.C(n_1388),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1442),
.B(n_1388),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1442),
.B(n_1392),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1427),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1454),
.A2(n_1418),
.B1(n_1408),
.B2(n_1373),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1475),
.A2(n_1367),
.B1(n_1418),
.B2(n_1408),
.Y(n_1492)
);

NAND3xp33_ASAP7_75t_L g1493 ( 
.A(n_1453),
.B(n_1406),
.C(n_1405),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1465),
.A2(n_1405),
.B1(n_1401),
.B2(n_1406),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1460),
.A2(n_1401),
.B1(n_1417),
.B2(n_1399),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1451),
.B(n_1383),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1438),
.B(n_1392),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1438),
.B(n_1395),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1457),
.B(n_1383),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1462),
.B(n_1382),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1430),
.A2(n_1401),
.B1(n_1417),
.B2(n_1400),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1439),
.B(n_1395),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1435),
.B(n_1420),
.C(n_1426),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1439),
.B(n_1372),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1461),
.B(n_1385),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1444),
.B(n_1385),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1467),
.B(n_1372),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1432),
.B(n_1426),
.C(n_1425),
.Y(n_1508)
);

NAND2x1_ASAP7_75t_L g1509 ( 
.A(n_1473),
.B(n_1363),
.Y(n_1509)
);

OAI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1432),
.A2(n_1424),
.B(n_1412),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1436),
.B(n_1363),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_SL g1512 ( 
.A(n_1440),
.B(n_1382),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1443),
.B(n_1397),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1456),
.B(n_1448),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1455),
.B(n_1425),
.C(n_1423),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1467),
.B(n_1377),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1447),
.B(n_1413),
.C(n_1423),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1469),
.B(n_1372),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1377),
.Y(n_1519)
);

OR2x2_ASAP7_75t_SL g1520 ( 
.A(n_1471),
.B(n_1472),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1450),
.B(n_1398),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1436),
.B(n_1363),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1468),
.B(n_1422),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1459),
.B(n_1374),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1429),
.Y(n_1525)
);

OAI21xp33_ASAP7_75t_L g1526 ( 
.A1(n_1455),
.A2(n_1419),
.B(n_1360),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1524),
.B(n_1473),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1498),
.B(n_1502),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1476),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1476),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1482),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1490),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.B(n_1507),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1490),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1507),
.B(n_1518),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1518),
.B(n_1473),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1504),
.B(n_1473),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1520),
.B(n_1446),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1504),
.B(n_1481),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1488),
.B(n_1446),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1481),
.B(n_1374),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1525),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1520),
.B(n_1445),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1487),
.B(n_1445),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1489),
.B(n_1374),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1489),
.B(n_1374),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1483),
.B(n_1387),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1525),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1509),
.B(n_1434),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1509),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1511),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1514),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1496),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1511),
.B(n_1522),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1484),
.B(n_1521),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1499),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1513),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1478),
.B(n_1470),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1505),
.Y(n_1560)
);

BUFx3_ASAP7_75t_L g1561 ( 
.A(n_1479),
.Y(n_1561)
);

BUFx2_ASAP7_75t_L g1562 ( 
.A(n_1479),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1485),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1560),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1551),
.B(n_1555),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1532),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1549),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1532),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1551),
.B(n_1458),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_SL g1571 ( 
.A1(n_1531),
.A2(n_1491),
.B(n_1480),
.C(n_1500),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1553),
.B(n_1516),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1553),
.B(n_1512),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1542),
.Y(n_1574)
);

OA211x2_ASAP7_75t_L g1575 ( 
.A1(n_1531),
.A2(n_1510),
.B(n_1526),
.C(n_1493),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1533),
.B(n_1485),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1540),
.B(n_1519),
.Y(n_1577)
);

OAI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1538),
.A2(n_1492),
.B(n_1477),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1529),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1560),
.B(n_1506),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1533),
.B(n_1486),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1508),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1558),
.B(n_1517),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1549),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1530),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_L g1588 ( 
.A(n_1554),
.B(n_1495),
.C(n_1494),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1530),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1549),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1556),
.B(n_1440),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1528),
.B(n_1470),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1540),
.B(n_1515),
.Y(n_1593)
);

INVxp67_ASAP7_75t_L g1594 ( 
.A(n_1554),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1530),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1549),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1534),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1543),
.B(n_1265),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1534),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1534),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1563),
.B(n_1555),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1566),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1588),
.B(n_1558),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1563),
.B(n_1555),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1577),
.B(n_1556),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1568),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1565),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1571),
.A2(n_1544),
.B(n_1543),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1574),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1576),
.B(n_1555),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1567),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1564),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1593),
.B(n_1544),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1593),
.B(n_1544),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1569),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1567),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1569),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1555),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1577),
.B(n_1538),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1594),
.B(n_1538),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1582),
.B(n_1543),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_L g1624 ( 
.A(n_1571),
.B(n_1363),
.Y(n_1624)
);

AOI211xp5_ASAP7_75t_L g1625 ( 
.A1(n_1573),
.A2(n_1501),
.B(n_1555),
.C(n_1554),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1591),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1587),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1575),
.A2(n_1536),
.B1(n_1527),
.B2(n_1559),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1587),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1572),
.B(n_1548),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1599),
.Y(n_1631)
);

NAND5xp2_ASAP7_75t_L g1632 ( 
.A(n_1598),
.B(n_1523),
.C(n_1536),
.D(n_1537),
.E(n_1546),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1578),
.B(n_1557),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1557),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1565),
.B(n_1539),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1599),
.Y(n_1636)
);

NAND2x1p5_ASAP7_75t_L g1637 ( 
.A(n_1584),
.B(n_1552),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1586),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1580),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1581),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1584),
.B(n_1557),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1589),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1565),
.B(n_1539),
.Y(n_1643)
);

BUFx3_ASAP7_75t_L g1644 ( 
.A(n_1614),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1615),
.B(n_1595),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1603),
.B(n_1583),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1617),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1619),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1633),
.B(n_1539),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1627),
.Y(n_1650)
);

NAND2xp33_ASAP7_75t_SL g1651 ( 
.A(n_1624),
.B(n_1340),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1635),
.B(n_1584),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1637),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1607),
.B(n_1570),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1629),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1626),
.B(n_1355),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1635),
.B(n_1643),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1631),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1637),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1607),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1643),
.B(n_1592),
.Y(n_1661)
);

BUFx2_ASAP7_75t_SL g1662 ( 
.A(n_1601),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1601),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1604),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1615),
.B(n_1597),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1604),
.B(n_1592),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1616),
.B(n_1600),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1609),
.B(n_1249),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1633),
.B(n_1528),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1636),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1639),
.Y(n_1671)
);

AND2x4_ASAP7_75t_L g1672 ( 
.A(n_1611),
.B(n_1570),
.Y(n_1672)
);

AOI22xp33_ASAP7_75t_L g1673 ( 
.A1(n_1624),
.A2(n_1527),
.B1(n_1437),
.B2(n_1436),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1616),
.B(n_1586),
.Y(n_1674)
);

INVxp67_ASAP7_75t_SL g1675 ( 
.A(n_1608),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1625),
.Y(n_1676)
);

CKINVDCx16_ASAP7_75t_R g1677 ( 
.A(n_1628),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1611),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1641),
.B(n_1528),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1632),
.A2(n_1620),
.B1(n_1623),
.B2(n_1605),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1668),
.B(n_1620),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1675),
.A2(n_1602),
.B1(n_1606),
.B2(n_1610),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1660),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1644),
.Y(n_1685)
);

NAND2xp33_ASAP7_75t_L g1686 ( 
.A(n_1676),
.B(n_1622),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1660),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1644),
.B(n_1634),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1646),
.B(n_1680),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1663),
.B(n_1613),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1651),
.A2(n_1622),
.B(n_1570),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1677),
.A2(n_1640),
.B1(n_1642),
.B2(n_1570),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1678),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1662),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1417),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1647),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1621),
.Y(n_1697)
);

AOI322xp5_ASAP7_75t_L g1698 ( 
.A1(n_1669),
.A2(n_1535),
.A3(n_1552),
.B1(n_1562),
.B2(n_1541),
.C1(n_1545),
.C2(n_1546),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1648),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1663),
.B(n_1621),
.Y(n_1700)
);

AOI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1653),
.A2(n_1618),
.B(n_1612),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1679),
.B(n_1630),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1657),
.B(n_1547),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1657),
.B(n_1547),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1648),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1650),
.Y(n_1706)
);

INVx1_ASAP7_75t_SL g1707 ( 
.A(n_1694),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1695),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1684),
.B(n_1687),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1684),
.Y(n_1710)
);

INVx3_ASAP7_75t_SL g1711 ( 
.A(n_1687),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1681),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1686),
.A2(n_1656),
.B(n_1653),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1696),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1695),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1685),
.B(n_1664),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1685),
.B(n_1664),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1682),
.B(n_1659),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1695),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1686),
.B(n_1678),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1699),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1700),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1693),
.B(n_1678),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1693),
.B(n_1652),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1688),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1689),
.B(n_1666),
.Y(n_1726)
);

OAI221xp5_ASAP7_75t_SL g1727 ( 
.A1(n_1707),
.A2(n_1683),
.B1(n_1692),
.B2(n_1698),
.C(n_1705),
.Y(n_1727)
);

NOR3x1_ASAP7_75t_L g1728 ( 
.A(n_1716),
.B(n_1690),
.C(n_1706),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1711),
.B(n_1682),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1718),
.A2(n_1726),
.B1(n_1722),
.B2(n_1691),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1713),
.A2(n_1720),
.B(n_1710),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1725),
.A2(n_1672),
.B1(n_1697),
.B2(n_1702),
.Y(n_1732)
);

AOI211xp5_ASAP7_75t_L g1733 ( 
.A1(n_1711),
.A2(n_1659),
.B(n_1671),
.C(n_1672),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1709),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1715),
.A2(n_1671),
.B1(n_1652),
.B2(n_1650),
.C(n_1655),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1723),
.Y(n_1736)
);

OAI21xp5_ASAP7_75t_SL g1737 ( 
.A1(n_1719),
.A2(n_1673),
.B(n_1672),
.Y(n_1737)
);

AO22x1_ASAP7_75t_L g1738 ( 
.A1(n_1723),
.A2(n_1654),
.B1(n_1658),
.B2(n_1670),
.Y(n_1738)
);

NOR4xp25_ASAP7_75t_L g1739 ( 
.A(n_1727),
.B(n_1709),
.C(n_1717),
.D(n_1721),
.Y(n_1739)
);

OAI21xp33_ASAP7_75t_L g1740 ( 
.A1(n_1727),
.A2(n_1724),
.B(n_1708),
.Y(n_1740)
);

NAND3xp33_ASAP7_75t_SL g1741 ( 
.A(n_1731),
.B(n_1724),
.C(n_1714),
.Y(n_1741)
);

AND3x1_ASAP7_75t_L g1742 ( 
.A(n_1733),
.B(n_1708),
.C(n_1712),
.Y(n_1742)
);

NAND3xp33_ASAP7_75t_SL g1743 ( 
.A(n_1730),
.B(n_1714),
.C(n_1712),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1736),
.B(n_1734),
.Y(n_1744)
);

NAND3xp33_ASAP7_75t_SL g1745 ( 
.A(n_1729),
.B(n_1721),
.C(n_1665),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1732),
.B(n_1728),
.Y(n_1746)
);

AOI22xp5_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1735),
.B1(n_1738),
.B2(n_1654),
.Y(n_1747)
);

NAND2x1p5_ASAP7_75t_L g1748 ( 
.A(n_1736),
.B(n_1270),
.Y(n_1748)
);

NOR3xp33_ASAP7_75t_L g1749 ( 
.A(n_1740),
.B(n_1299),
.C(n_1701),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_SL g1750 ( 
.A(n_1741),
.B(n_1658),
.C(n_1655),
.Y(n_1750)
);

AOI222xp33_ASAP7_75t_L g1751 ( 
.A1(n_1746),
.A2(n_1670),
.B1(n_1654),
.B2(n_1703),
.C1(n_1704),
.C2(n_1666),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1739),
.A2(n_1674),
.B1(n_1667),
.B2(n_1665),
.C(n_1645),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1747),
.A2(n_1674),
.B(n_1645),
.C(n_1667),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1742),
.A2(n_1661),
.B(n_1618),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_SL g1755 ( 
.A(n_1743),
.B(n_1286),
.C(n_1503),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1750),
.A2(n_1748),
.B1(n_1744),
.B2(n_1661),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1754),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1751),
.Y(n_1758)
);

NOR2x1_ASAP7_75t_L g1759 ( 
.A(n_1753),
.B(n_1745),
.Y(n_1759)
);

AOI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1749),
.A2(n_1638),
.B1(n_1612),
.B2(n_1552),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1752),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1755),
.B(n_1638),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_SL g1763 ( 
.A(n_1759),
.B(n_1341),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1757),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1756),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_SL g1766 ( 
.A(n_1758),
.B(n_1341),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1760),
.Y(n_1767)
);

XNOR2xp5_ASAP7_75t_L g1768 ( 
.A(n_1765),
.B(n_1761),
.Y(n_1768)
);

XNOR2x1_ASAP7_75t_L g1769 ( 
.A(n_1767),
.B(n_1762),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1764),
.Y(n_1770)
);

XNOR2x1_ASAP7_75t_L g1771 ( 
.A(n_1768),
.B(n_1766),
.Y(n_1771)
);

OAI22x1_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1770),
.B1(n_1763),
.B2(n_1769),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1772),
.B(n_1763),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1772),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1596),
.B1(n_1590),
.B2(n_1401),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1773),
.B(n_1308),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1596),
.B(n_1590),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1775),
.Y(n_1778)
);

OAI21xp33_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1561),
.B(n_1550),
.Y(n_1779)
);

AOI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1777),
.B1(n_1308),
.B2(n_1328),
.C1(n_1322),
.C2(n_1562),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_R g1781 ( 
.A1(n_1780),
.A2(n_1401),
.B1(n_1562),
.B2(n_1550),
.C(n_1561),
.Y(n_1781)
);

AOI211xp5_ASAP7_75t_L g1782 ( 
.A1(n_1781),
.A2(n_1288),
.B(n_1354),
.C(n_1258),
.Y(n_1782)
);


endmodule