module fake_jpeg_31608_n_506 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_506);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_506;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx13_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_53),
.B(n_62),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_21),
.B(n_1),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_2),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_42),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_65),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_2),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_66),
.B(n_90),
.Y(n_136)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g168 ( 
.A(n_78),
.Y(n_168)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx2_ASAP7_75t_SL g123 ( 
.A(n_80),
.Y(n_123)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_4),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_97),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_16),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_102),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_17),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_103),
.Y(n_155)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_104),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_106),
.Y(n_154)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

AOI21xp33_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_51),
.B(n_20),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_116),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_27),
.B1(n_47),
.B2(n_43),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_110),
.A2(n_118),
.B1(n_43),
.B2(n_39),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_26),
.B1(n_47),
.B2(n_23),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_112),
.A2(n_141),
.B1(n_152),
.B2(n_39),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_166),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_57),
.A2(n_63),
.B1(n_69),
.B2(n_65),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_54),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_147),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_59),
.A2(n_17),
.B1(n_24),
.B2(n_37),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_133),
.A2(n_45),
.B1(n_85),
.B2(n_101),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_17),
.B1(n_30),
.B2(n_41),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_94),
.C(n_95),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_83),
.A2(n_41),
.B1(n_51),
.B2(n_31),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g158 ( 
.A(n_80),
.Y(n_158)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_98),
.B(n_26),
.Y(n_166)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_173),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_139),
.Y(n_174)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_138),
.B1(n_20),
.B2(n_36),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_178),
.A2(n_182),
.B1(n_191),
.B2(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_179),
.B(n_186),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_159),
.A2(n_36),
.B1(n_35),
.B2(n_32),
.Y(n_182)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

INVx11_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_37),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_45),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_135),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_188),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_189),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_163),
.Y(n_190)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_166),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_196),
.Y(n_232)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_131),
.Y(n_195)
);

INVx13_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_199),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_198),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_134),
.B(n_42),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_216),
.Y(n_238)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_202),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_117),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_212),
.B1(n_155),
.B2(n_144),
.Y(n_237)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_148),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_204),
.B(n_205),
.Y(n_252)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

BUFx6f_ASAP7_75t_SL g227 ( 
.A(n_206),
.Y(n_227)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_207),
.Y(n_253)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_124),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_118),
.A2(n_102),
.B1(n_88),
.B2(n_87),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_214),
.B1(n_115),
.B2(n_128),
.Y(n_245)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_119),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_130),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_213),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_41),
.B1(n_38),
.B2(n_15),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_134),
.B(n_15),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_38),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_137),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_137),
.B(n_38),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_218),
.A2(n_152),
.B(n_133),
.C(n_141),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_228),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_157),
.B1(n_150),
.B2(n_165),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_144),
.B(n_154),
.C(n_155),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_239),
.A2(n_172),
.B(n_183),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_154),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_242),
.Y(n_258)
);

NAND3xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_243),
.C(n_232),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_181),
.B(n_149),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_113),
.B1(n_142),
.B2(n_145),
.Y(n_277)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_209),
.A2(n_122),
.B1(n_126),
.B2(n_125),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_212),
.Y(n_268)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_256),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_185),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_257),
.B(n_260),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_229),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_259),
.B(n_262),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_175),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_221),
.B(n_184),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_187),
.C(n_176),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_263),
.B(n_264),
.C(n_271),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_221),
.B(n_194),
.C(n_192),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_188),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_267),
.B(n_269),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_233),
.Y(n_270)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_270),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_200),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_238),
.B(n_216),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_238),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_279),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_220),
.B1(n_246),
.B2(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_233),
.Y(n_275)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_280),
.B1(n_281),
.B2(n_286),
.Y(n_289)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_223),
.Y(n_278)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

O2A1O1Ixp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_196),
.B(n_195),
.C(n_198),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_169),
.B1(n_207),
.B2(n_217),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_237),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_213),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_282),
.B(n_246),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_239),
.B(n_251),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_223),
.Y(n_285)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_285),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_228),
.A2(n_189),
.B1(n_168),
.B2(n_211),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_288),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_226),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_290),
.B(n_297),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_293),
.A2(n_315),
.B1(n_251),
.B2(n_231),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_262),
.B(n_252),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_256),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_299),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_252),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_229),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_300),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_236),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_301),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_272),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_307),
.Y(n_329)
);

AO22x2_ASAP7_75t_L g307 ( 
.A1(n_276),
.A2(n_228),
.B1(n_246),
.B2(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_272),
.Y(n_310)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_258),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_313),
.A2(n_282),
.B(n_274),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_268),
.A2(n_246),
.B1(n_239),
.B2(n_220),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_296),
.A2(n_276),
.B(n_283),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_320),
.B(n_321),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_292),
.B(n_258),
.Y(n_319)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_319),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_296),
.A2(n_313),
.B(n_310),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_269),
.B(n_273),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_322),
.B(n_332),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_268),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_312),
.A2(n_286),
.B(n_279),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_326),
.Y(n_368)
);

XNOR2x1_ASAP7_75t_SL g328 ( 
.A(n_314),
.B(n_260),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_328),
.B(n_292),
.Y(n_346)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_287),
.B(n_281),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_342),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_335),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_302),
.A2(n_285),
.B(n_278),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_311),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_289),
.A2(n_277),
.B1(n_280),
.B2(n_261),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_337),
.A2(n_341),
.B1(n_294),
.B2(n_311),
.Y(n_350)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_284),
.B(n_275),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_338),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_339),
.A2(n_326),
.B1(n_323),
.B2(n_325),
.Y(n_355)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_294),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_309),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_289),
.A2(n_270),
.B1(n_224),
.B2(n_247),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_250),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_295),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_343),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_332),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_306),
.B1(n_293),
.B2(n_308),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_350),
.A2(n_325),
.B1(n_337),
.B2(n_341),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_354),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_304),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_353),
.C(n_366),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_304),
.C(n_308),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_355),
.A2(n_362),
.B1(n_367),
.B2(n_254),
.Y(n_396)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_357),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_319),
.B(n_309),
.Y(n_359)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_359),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_339),
.A2(n_307),
.B1(n_303),
.B2(n_295),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_335),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_365),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_318),
.B(n_303),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_307),
.C(n_250),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_323),
.A2(n_307),
.B1(n_305),
.B2(n_265),
.Y(n_367)
);

AO22x1_ASAP7_75t_SL g369 ( 
.A1(n_329),
.A2(n_307),
.B1(n_224),
.B2(n_230),
.Y(n_369)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_369),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_253),
.Y(n_371)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

BUFx12_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_368),
.A2(n_329),
.B(n_316),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_384),
.Y(n_406)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_356),
.Y(n_378)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_378),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_371),
.B(n_324),
.Y(n_380)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_343),
.Y(n_381)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_383),
.A2(n_358),
.B1(n_369),
.B2(n_219),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_368),
.A2(n_320),
.B(n_336),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_345),
.B(n_330),
.C(n_327),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_388),
.C(n_360),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_340),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_391),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_345),
.B(n_330),
.C(n_327),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_361),
.B(n_333),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_394),
.B1(n_399),
.B2(n_230),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_321),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_328),
.B1(n_224),
.B2(n_253),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_393),
.A2(n_396),
.B1(n_219),
.B2(n_227),
.Y(n_415)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_370),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_344),
.B(n_254),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_395),
.B(n_355),
.Y(n_400)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_372),
.Y(n_399)
);

XOR2x2_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_376),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_398),
.A2(n_350),
.B1(n_346),
.B2(n_349),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_401),
.B(n_402),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_352),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_408),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_366),
.C(n_353),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_405),
.C(n_414),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_388),
.C(n_373),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_390),
.A2(n_358),
.B(n_362),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_407),
.B(n_419),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_393),
.B(n_360),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_410),
.A2(n_377),
.B1(n_394),
.B2(n_399),
.Y(n_431)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_412),
.Y(n_422)
);

NOR2xp67_ASAP7_75t_SL g413 ( 
.A(n_379),
.B(n_369),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_413),
.B(n_375),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_384),
.C(n_392),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_415),
.A2(n_382),
.B1(n_387),
.B2(n_395),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_227),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_390),
.A2(n_234),
.B1(n_244),
.B2(n_170),
.Y(n_420)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_420),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_383),
.A2(n_244),
.B1(n_234),
.B2(n_122),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_421),
.B(n_378),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_409),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_435),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_396),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_436),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_417),
.A2(n_392),
.B1(n_382),
.B2(n_387),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_427),
.A2(n_431),
.B1(n_438),
.B2(n_415),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_428),
.A2(n_422),
.B1(n_439),
.B2(n_434),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_414),
.A2(n_381),
.B(n_391),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_429),
.A2(n_406),
.B(n_418),
.Y(n_443)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_432),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_386),
.C(n_389),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_437),
.C(n_402),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_409),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_376),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_440),
.B(n_448),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_441),
.B(n_444),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_442),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_443),
.A2(n_423),
.B(n_248),
.Y(n_459)
);

FAx1_ASAP7_75t_SL g444 ( 
.A(n_433),
.B(n_405),
.CI(n_407),
.CON(n_444),
.SN(n_444)
);

XOR2x2_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_400),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_445),
.B(n_248),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_437),
.B(n_411),
.C(n_419),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_449),
.C(n_456),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_424),
.B(n_429),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_416),
.C(n_376),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_451),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_439),
.B(n_378),
.Y(n_451)
);

OAI321xp33_ASAP7_75t_L g453 ( 
.A1(n_428),
.A2(n_234),
.A3(n_248),
.B1(n_126),
.B2(n_10),
.C(n_11),
.Y(n_453)
);

BUFx24_ASAP7_75t_SL g458 ( 
.A(n_453),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_4),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_455),
.B(n_4),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_423),
.B(n_151),
.C(n_143),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_454),
.A2(n_430),
.B(n_436),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_457),
.A2(n_6),
.B(n_9),
.Y(n_480)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_459),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_461),
.B(n_465),
.Y(n_482)
);

INVx11_ASAP7_75t_L g463 ( 
.A(n_451),
.Y(n_463)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_464),
.B(n_469),
.Y(n_472)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_442),
.A2(n_447),
.B1(n_445),
.B2(n_452),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_471),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_449),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_447),
.B(n_115),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_462),
.B(n_446),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_474),
.B(n_475),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_468),
.B(n_456),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_15),
.C(n_9),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_476),
.B(n_481),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_478),
.A2(n_470),
.B1(n_463),
.B2(n_466),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_480),
.A2(n_6),
.B1(n_10),
.B2(n_12),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_15),
.C(n_180),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_458),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_483),
.B(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_486),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_482),
.B(n_466),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_487),
.B(n_488),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_472),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_15),
.C(n_12),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_490),
.A2(n_10),
.B(n_12),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_180),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_491),
.A2(n_473),
.B(n_481),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_493),
.B(n_496),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_12),
.Y(n_499)
);

OAI21x1_ASAP7_75t_L g497 ( 
.A1(n_492),
.A2(n_491),
.B(n_479),
.Y(n_497)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_497),
.A2(n_499),
.B(n_495),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_500),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_484),
.C(n_485),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_502),
.B(n_501),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_503),
.A2(n_38),
.B(n_13),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_14),
.Y(n_505)
);

O2A1O1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_505),
.A2(n_14),
.B(n_504),
.C(n_482),
.Y(n_506)
);


endmodule