module fake_netlist_5_503_n_3727 (n_137, n_924, n_676, n_294, n_431, n_318, n_380, n_419, n_977, n_653, n_611, n_444, n_642, n_469, n_615, n_851, n_82, n_194, n_316, n_785, n_389, n_843, n_855, n_549, n_684, n_850, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_865, n_61, n_913, n_678, n_664, n_376, n_697, n_503, n_967, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_928, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_916, n_452, n_885, n_397, n_493, n_111, n_525, n_880, n_703, n_698, n_980, n_483, n_544, n_683, n_1007, n_155, n_780, n_649, n_552, n_547, n_43, n_721, n_998, n_116, n_841, n_956, n_22, n_467, n_564, n_802, n_423, n_840, n_284, n_46, n_245, n_21, n_501, n_823, n_725, n_983, n_139, n_38, n_105, n_280, n_744, n_590, n_629, n_672, n_4, n_873, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_898, n_254, n_690, n_33, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_526, n_915, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_859, n_864, n_951, n_821, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_909, n_625, n_854, n_949, n_621, n_753, n_997, n_100, n_455, n_674, n_1008, n_932, n_417, n_946, n_612, n_1001, n_212, n_385, n_498, n_516, n_933, n_788, n_507, n_119, n_497, n_689, n_738, n_912, n_606, n_559, n_275, n_640, n_968, n_252, n_624, n_825, n_26, n_295, n_133, n_1010, n_330, n_877, n_508, n_739, n_506, n_2, n_737, n_610, n_972, n_692, n_986, n_755, n_6, n_509, n_568, n_936, n_39, n_147, n_373, n_820, n_757, n_947, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_758, n_999, n_668, n_733, n_991, n_375, n_301, n_828, n_779, n_576, n_941, n_929, n_981, n_68, n_804, n_93, n_867, n_186, n_537, n_134, n_902, n_191, n_587, n_945, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_878, n_524, n_943, n_399, n_341, n_204, n_394, n_250, n_579, n_992, n_938, n_741, n_548, n_543, n_260, n_812, n_842, n_298, n_650, n_984, n_320, n_694, n_518, n_505, n_286, n_883, n_122, n_282, n_752, n_331, n_10, n_905, n_906, n_24, n_406, n_519, n_470, n_908, n_782, n_919, n_325, n_449, n_132, n_862, n_90, n_900, n_724, n_856, n_546, n_101, n_760, n_658, n_281, n_918, n_240, n_942, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_959, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_940, n_896, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_920, n_894, n_271, n_934, n_94, n_831, n_826, n_335, n_123, n_886, n_978, n_964, n_654, n_370, n_167, n_976, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_833, n_297, n_156, n_5, n_853, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_988, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_1009, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_961, n_995, n_955, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_882, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_897, n_215, n_350, n_196, n_798, n_662, n_459, n_646, n_211, n_218, n_400, n_930, n_181, n_436, n_962, n_3, n_290, n_580, n_221, n_178, n_622, n_723, n_386, n_578, n_994, n_926, n_287, n_344, n_848, n_555, n_783, n_473, n_422, n_475, n_777, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_496, n_355, n_958, n_849, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_922, n_145, n_48, n_521, n_614, n_663, n_845, n_50, n_337, n_430, n_313, n_631, n_673, n_837, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_974, n_395, n_164, n_432, n_553, n_727, n_839, n_901, n_311, n_813, n_957, n_830, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_888, n_296, n_613, n_871, n_241, n_637, n_357, n_875, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_829, n_144, n_858, n_114, n_96, n_923, n_772, n_691, n_881, n_717, n_165, n_468, n_499, n_939, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_866, n_969, n_236, n_388, n_761, n_1012, n_1, n_249, n_903, n_1006, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_889, n_80, n_973, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_836, n_990, n_84, n_462, n_975, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_907, n_722, n_458, n_288, n_770, n_188, n_190, n_844, n_201, n_263, n_471, n_609, n_852, n_989, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_711, n_781, n_834, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_892, n_893, n_1000, n_891, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_979, n_1002, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_846, n_874, n_465, n_838, n_76, n_358, n_362, n_876, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_953, n_601, n_279, n_917, n_966, n_70, n_987, n_253, n_261, n_174, n_289, n_745, n_963, n_954, n_627, n_767, n_172, n_206, n_217, n_993, n_440, n_726, n_478, n_793, n_545, n_982, n_441, n_860, n_450, n_648, n_312, n_476, n_818, n_429, n_861, n_534, n_948, n_884, n_899, n_345, n_210, n_944, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_176, n_970, n_911, n_557, n_182, n_143, n_83, n_1005, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_832, n_180, n_857, n_560, n_656, n_340, n_207, n_561, n_37, n_346, n_937, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_879, n_16, n_720, n_0, n_58, n_623, n_405, n_824, n_18, n_359, n_863, n_910, n_971, n_490, n_805, n_117, n_326, n_794, n_768, n_921, n_996, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_847, n_815, n_246, n_596, n_179, n_125, n_410, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_822, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_895, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_887, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_870, n_931, n_159, n_334, n_599, n_766, n_811, n_952, n_541, n_807, n_391, n_701, n_434, n_645, n_539, n_835, n_175, n_538, n_666, n_262, n_803, n_868, n_238, n_639, n_799, n_914, n_99, n_687, n_715, n_411, n_414, n_319, n_364, n_965, n_927, n_20, n_536, n_531, n_935, n_1004, n_121, n_242, n_817, n_872, n_360, n_36, n_594, n_764, n_200, n_890, n_162, n_960, n_64, n_759, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_1011, n_904, n_985, n_869, n_324, n_810, n_634, n_416, n_199, n_827, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_925, n_424, n_1003, n_7, n_706, n_746, n_256, n_305, n_533, n_950, n_747, n_52, n_278, n_784, n_110, n_3727);

input n_137;
input n_924;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_977;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_851;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_843;
input n_855;
input n_549;
input n_684;
input n_850;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_865;
input n_61;
input n_913;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_967;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_928;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_916;
input n_452;
input n_885;
input n_397;
input n_493;
input n_111;
input n_525;
input n_880;
input n_703;
input n_698;
input n_980;
input n_483;
input n_544;
input n_683;
input n_1007;
input n_155;
input n_780;
input n_649;
input n_552;
input n_547;
input n_43;
input n_721;
input n_998;
input n_116;
input n_841;
input n_956;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_840;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_823;
input n_725;
input n_983;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_590;
input n_629;
input n_672;
input n_4;
input n_873;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_898;
input n_254;
input n_690;
input n_33;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_526;
input n_915;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_859;
input n_864;
input n_951;
input n_821;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_909;
input n_625;
input n_854;
input n_949;
input n_621;
input n_753;
input n_997;
input n_100;
input n_455;
input n_674;
input n_1008;
input n_932;
input n_417;
input n_946;
input n_612;
input n_1001;
input n_212;
input n_385;
input n_498;
input n_516;
input n_933;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_912;
input n_606;
input n_559;
input n_275;
input n_640;
input n_968;
input n_252;
input n_624;
input n_825;
input n_26;
input n_295;
input n_133;
input n_1010;
input n_330;
input n_877;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_972;
input n_692;
input n_986;
input n_755;
input n_6;
input n_509;
input n_568;
input n_936;
input n_39;
input n_147;
input n_373;
input n_820;
input n_757;
input n_947;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_999;
input n_668;
input n_733;
input n_991;
input n_375;
input n_301;
input n_828;
input n_779;
input n_576;
input n_941;
input n_929;
input n_981;
input n_68;
input n_804;
input n_93;
input n_867;
input n_186;
input n_537;
input n_134;
input n_902;
input n_191;
input n_587;
input n_945;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_878;
input n_524;
input n_943;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_992;
input n_938;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_842;
input n_298;
input n_650;
input n_984;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_883;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_905;
input n_906;
input n_24;
input n_406;
input n_519;
input n_470;
input n_908;
input n_782;
input n_919;
input n_325;
input n_449;
input n_132;
input n_862;
input n_90;
input n_900;
input n_724;
input n_856;
input n_546;
input n_101;
input n_760;
input n_658;
input n_281;
input n_918;
input n_240;
input n_942;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_959;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_940;
input n_896;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_920;
input n_894;
input n_271;
input n_934;
input n_94;
input n_831;
input n_826;
input n_335;
input n_123;
input n_886;
input n_978;
input n_964;
input n_654;
input n_370;
input n_167;
input n_976;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_833;
input n_297;
input n_156;
input n_5;
input n_853;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_988;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_1009;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_961;
input n_995;
input n_955;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_882;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_646;
input n_211;
input n_218;
input n_400;
input n_930;
input n_181;
input n_436;
input n_962;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_723;
input n_386;
input n_578;
input n_994;
input n_926;
input n_287;
input n_344;
input n_848;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_958;
input n_849;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_922;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_845;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_837;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_974;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_839;
input n_901;
input n_311;
input n_813;
input n_957;
input n_830;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_888;
input n_296;
input n_613;
input n_871;
input n_241;
input n_637;
input n_357;
input n_875;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_829;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_772;
input n_691;
input n_881;
input n_717;
input n_165;
input n_468;
input n_499;
input n_939;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_866;
input n_969;
input n_236;
input n_388;
input n_761;
input n_1012;
input n_1;
input n_249;
input n_903;
input n_1006;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_889;
input n_80;
input n_973;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_836;
input n_990;
input n_84;
input n_462;
input n_975;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_907;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_844;
input n_201;
input n_263;
input n_471;
input n_609;
input n_852;
input n_989;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_711;
input n_781;
input n_834;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_892;
input n_893;
input n_1000;
input n_891;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_979;
input n_1002;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_846;
input n_874;
input n_465;
input n_838;
input n_76;
input n_358;
input n_362;
input n_876;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_953;
input n_601;
input n_279;
input n_917;
input n_966;
input n_70;
input n_987;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_963;
input n_954;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_993;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_982;
input n_441;
input n_860;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_861;
input n_534;
input n_948;
input n_884;
input n_899;
input n_345;
input n_210;
input n_944;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_176;
input n_970;
input n_911;
input n_557;
input n_182;
input n_143;
input n_83;
input n_1005;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_832;
input n_180;
input n_857;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_937;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_879;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_824;
input n_18;
input n_359;
input n_863;
input n_910;
input n_971;
input n_490;
input n_805;
input n_117;
input n_326;
input n_794;
input n_768;
input n_921;
input n_996;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_847;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_822;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_895;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_887;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_870;
input n_931;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_952;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_645;
input n_539;
input n_835;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_868;
input n_238;
input n_639;
input n_799;
input n_914;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_319;
input n_364;
input n_965;
input n_927;
input n_20;
input n_536;
input n_531;
input n_935;
input n_1004;
input n_121;
input n_242;
input n_817;
input n_872;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_890;
input n_162;
input n_960;
input n_64;
input n_759;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_1011;
input n_904;
input n_985;
input n_869;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_827;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_925;
input n_424;
input n_1003;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_950;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_3727;

wire n_1263;
wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_1488;
wire n_2955;
wire n_2899;
wire n_3619;
wire n_1055;
wire n_3541;
wire n_3622;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_3086;
wire n_3297;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_3641;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_1545;
wire n_2374;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_1285;
wire n_3710;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_3036;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1705;
wire n_1294;
wire n_1104;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_3650;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_2091;
wire n_1517;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_3631;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_3490;
wire n_3656;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_2099;
wire n_2408;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_3702;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_1547;
wire n_1070;
wire n_2089;
wire n_3420;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_1034;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_2235;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_2432;
wire n_3668;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_1880;
wire n_2769;
wire n_3542;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3550;
wire n_2615;
wire n_1556;
wire n_1384;
wire n_1863;
wire n_1064;
wire n_2079;
wire n_2238;
wire n_2118;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_2358;
wire n_3716;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_3593;
wire n_3193;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_3496;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_3714;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_3071;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_1058;
wire n_3359;
wire n_2784;
wire n_3718;
wire n_2919;
wire n_3092;
wire n_1053;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_1014;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_3598;
wire n_1052;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_1754;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_3433;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_2305;
wire n_3392;
wire n_3430;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1027;
wire n_1156;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_2837;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_3655;
wire n_2808;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_3640;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1847;
wire n_1199;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_3602;
wire n_1038;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_2454;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_1876;
wire n_1743;
wire n_3491;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_3643;
wire n_2222;
wire n_1892;
wire n_3510;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_1189;
wire n_2690;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_3150;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_1537;
wire n_2227;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_3416;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_3469;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_2539;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1539;
wire n_2736;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1744;
wire n_1380;
wire n_2623;
wire n_1617;
wire n_1994;
wire n_1231;
wire n_1406;
wire n_1279;
wire n_3113;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_3457;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3555;
wire n_3579;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_2459;
wire n_3031;
wire n_3396;
wire n_3701;
wire n_1445;
wire n_3516;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_1079;
wire n_2093;
wire n_2320;
wire n_1045;
wire n_1208;
wire n_2473;
wire n_2038;
wire n_2339;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_1159;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3149;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_2418;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3411;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_3645;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_3474;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_1015;
wire n_1140;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_3679;
wire n_2464;
wire n_3422;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_3229;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1534;
wire n_1354;
wire n_2288;
wire n_3421;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3592;
wire n_3618;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_3394;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_3546;
wire n_1206;
wire n_2647;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3548;
wire n_2440;
wire n_1699;
wire n_1386;
wire n_3334;
wire n_1442;
wire n_2923;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_1050;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_1305;
wire n_3178;
wire n_1826;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3282;
wire n_2472;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3299;
wire n_3041;
wire n_3274;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1668;
wire n_1363;
wire n_1185;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1439;
wire n_1312;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_2997;
wire n_3327;
wire n_1504;
wire n_3326;
wire n_3572;
wire n_3067;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_3167;
wire n_3400;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_3529;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_3078;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_2280;
wire n_2192;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1865;
wire n_1511;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2318;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_2707;
wire n_2751;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3708;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_2795;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3380;
wire n_3177;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_3393;
wire n_1603;
wire n_1232;
wire n_2638;
wire n_1401;
wire n_3520;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_1122;
wire n_3192;
wire n_2608;
wire n_2657;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1929;
wire n_1392;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_1190;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_2409;
wire n_3450;
wire n_1714;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_3174;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_2217;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1777;
wire n_1335;
wire n_1514;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_2148;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3308;
wire n_2665;
wire n_1543;
wire n_1399;
wire n_1991;
wire n_1979;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_2484;
wire n_3530;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_3534;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_3438;
wire n_2012;
wire n_1291;
wire n_3381;
wire n_3503;
wire n_1753;
wire n_1297;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_2103;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_3397;
wire n_2363;
wire n_2430;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_3431;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_3700;
wire n_3609;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1715;
wire n_1518;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_3584;
wire n_1425;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_1867;
wire n_1330;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_1618;
wire n_2260;
wire n_2447;
wire n_1813;
wire n_2343;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_1873;
wire n_1411;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_3391;
wire n_1567;
wire n_2567;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_1648;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_3627;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_2957;
wire n_1769;
wire n_3551;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3722;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_3251;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_3384;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1028;
wire n_1601;
wire n_3336;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_3250;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_2594;
wire n_3125;
wire n_3114;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_3556;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3591;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3266;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_3726;
wire n_2210;
wire n_3247;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_1558;
wire n_3225;
wire n_3321;
wire n_2166;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_1026;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1180;
wire n_1827;
wire n_3360;
wire n_2524;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_3159;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_624),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_953),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_785),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_207),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_279),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_202),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_639),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_993),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_490),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_329),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1004),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_655),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_99),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_488),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_226),
.Y(n_1027)
);

BUFx3_ASAP7_75t_L g1028 ( 
.A(n_530),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_458),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_610),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_923),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_613),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_630),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_597),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_952),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_310),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_378),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_354),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_738),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_632),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_429),
.Y(n_1041)
);

BUFx5_ASAP7_75t_L g1042 ( 
.A(n_982),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_48),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_676),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_943),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_414),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_618),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_864),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_780),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_856),
.Y(n_1050)
);

BUFx10_ASAP7_75t_L g1051 ( 
.A(n_951),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_93),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_538),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_852),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_905),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_57),
.Y(n_1056)
);

CKINVDCx16_ASAP7_75t_R g1057 ( 
.A(n_595),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_308),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_166),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_451),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_6),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_669),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_921),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_570),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_151),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_726),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_799),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_934),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_328),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_949),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_119),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_763),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_277),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_515),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_277),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_978),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_479),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_524),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_917),
.Y(n_1079)
);

CKINVDCx14_ASAP7_75t_R g1080 ( 
.A(n_689),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_829),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_1003),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_913),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_15),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_880),
.Y(n_1085)
);

CKINVDCx16_ASAP7_75t_R g1086 ( 
.A(n_724),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_411),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_341),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_765),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_927),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_503),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_881),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_6),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_486),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_994),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_184),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_957),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_0),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_989),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_841),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_343),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_695),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_223),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_420),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_572),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_398),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_843),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_176),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_54),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_495),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_838),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_748),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_892),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_629),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_890),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_335),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_631),
.Y(n_1117)
);

BUFx10_ASAP7_75t_L g1118 ( 
.A(n_101),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_770),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_752),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_908),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_186),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_691),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_375),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_625),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_946),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_461),
.Y(n_1127)
);

CKINVDCx20_ASAP7_75t_R g1128 ( 
.A(n_684),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_911),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_924),
.Y(n_1130)
);

BUFx3_ASAP7_75t_L g1131 ( 
.A(n_603),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_193),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_919),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_156),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_459),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_621),
.Y(n_1136)
);

CKINVDCx20_ASAP7_75t_R g1137 ( 
.A(n_860),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_196),
.Y(n_1138)
);

INVx1_ASAP7_75t_SL g1139 ( 
.A(n_998),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_183),
.Y(n_1140)
);

INVxp67_ASAP7_75t_L g1141 ( 
.A(n_956),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_996),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_935),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_965),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_147),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_786),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_266),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_700),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_160),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1002),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_608),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_623),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_947),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_112),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_462),
.Y(n_1155)
);

INVx1_ASAP7_75t_SL g1156 ( 
.A(n_209),
.Y(n_1156)
);

CKINVDCx20_ASAP7_75t_R g1157 ( 
.A(n_177),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_402),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_50),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_14),
.Y(n_1160)
);

CKINVDCx14_ASAP7_75t_R g1161 ( 
.A(n_635),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_363),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_666),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_631),
.Y(n_1164)
);

CKINVDCx20_ASAP7_75t_R g1165 ( 
.A(n_592),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_60),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_959),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_412),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_634),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_12),
.Y(n_1170)
);

BUFx5_ASAP7_75t_L g1171 ( 
.A(n_332),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_906),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_196),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_603),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_516),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_939),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_955),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_810),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_94),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_781),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_914),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_836),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_515),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_922),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_930),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_976),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1009),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_341),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_164),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_699),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_928),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_463),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_995),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_137),
.Y(n_1194)
);

BUFx5_ASAP7_75t_L g1195 ( 
.A(n_647),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_343),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_620),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_320),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_609),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_283),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_532),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_617),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_519),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_159),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_743),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_739),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_635),
.Y(n_1207)
);

INVx1_ASAP7_75t_SL g1208 ( 
.A(n_926),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_263),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_594),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_977),
.Y(n_1211)
);

BUFx10_ASAP7_75t_L g1212 ( 
.A(n_954),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_678),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_790),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_933),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_909),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_615),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_201),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_702),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_594),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_941),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_478),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_207),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_223),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_962),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_418),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_529),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_62),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_434),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_454),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_170),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_971),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_367),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_640),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_664),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_536),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_628),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_108),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1010),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_641),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_214),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_985),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_875),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_139),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_220),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_293),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_174),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_910),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_404),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_747),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_410),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_794),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_997),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_291),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_611),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_344),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_78),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_40),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_903),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_349),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_335),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_105),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_580),
.Y(n_1263)
);

BUFx2_ASAP7_75t_L g1264 ( 
.A(n_191),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_418),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_972),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_685),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_612),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_564),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_286),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_768),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_944),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_324),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_267),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_356),
.Y(n_1275)
);

CKINVDCx16_ASAP7_75t_R g1276 ( 
.A(n_374),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_162),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_518),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_445),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_46),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_622),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_481),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_606),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_735),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_915),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1001),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_820),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_618),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_252),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_529),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_98),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_942),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_821),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_969),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_391),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_987),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_620),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_250),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_471),
.Y(n_1299)
);

CKINVDCx20_ASAP7_75t_R g1300 ( 
.A(n_656),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_925),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_506),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_171),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_1000),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_505),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_576),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_945),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_528),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_99),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1005),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_65),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_761),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_286),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_197),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_1011),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_698),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_975),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_598),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_628),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_642),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_382),
.Y(n_1321)
);

INVx2_ASAP7_75t_L g1322 ( 
.A(n_301),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_643),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_974),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_940),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_983),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_330),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_322),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_461),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_948),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_142),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_600),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_84),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_92),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_897),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_32),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_990),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_309),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_629),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_931),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_912),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_937),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_963),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_531),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_381),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_828),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_577),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_999),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_488),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_517),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_410),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_156),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_287),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_932),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_750),
.Y(n_1355)
);

CKINVDCx20_ASAP7_75t_R g1356 ( 
.A(n_212),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_166),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_970),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_258),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_151),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_633),
.Y(n_1361)
);

BUFx2_ASAP7_75t_SL g1362 ( 
.A(n_503),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_938),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_627),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_824),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_832),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_379),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_420),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_973),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_98),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_746),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_688),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_708),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_179),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_636),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_67),
.Y(n_1376)
);

BUFx3_ASAP7_75t_L g1377 ( 
.A(n_314),
.Y(n_1377)
);

CKINVDCx16_ASAP7_75t_R g1378 ( 
.A(n_968),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_540),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_187),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_518),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_607),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_855),
.Y(n_1383)
);

CKINVDCx16_ASAP7_75t_R g1384 ( 
.A(n_614),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_79),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_346),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_80),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_979),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_80),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_657),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_176),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_205),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_104),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_63),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_263),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_441),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_188),
.Y(n_1397)
);

BUFx10_ASAP7_75t_L g1398 ( 
.A(n_578),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_425),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_809),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_984),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_961),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_88),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_578),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_339),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_395),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_774),
.Y(n_1407)
);

BUFx10_ASAP7_75t_L g1408 ( 
.A(n_66),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_283),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_65),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_487),
.Y(n_1411)
);

BUFx6f_ASAP7_75t_L g1412 ( 
.A(n_960),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_367),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_187),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_887),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_619),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_7),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_319),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_986),
.Y(n_1419)
);

BUFx5_ASAP7_75t_L g1420 ( 
.A(n_68),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_638),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_429),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_536),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_599),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_585),
.Y(n_1425)
);

INVxp67_ASAP7_75t_SL g1426 ( 
.A(n_648),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_532),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_958),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_67),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_626),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_964),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_81),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_382),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_607),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_988),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_825),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_281),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_252),
.Y(n_1438)
);

INVxp67_ASAP7_75t_L g1439 ( 
.A(n_697),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_967),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_869),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_719),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_125),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_632),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_472),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_373),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_31),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_177),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_991),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_653),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_936),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_21),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_528),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_430),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_992),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_118),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_481),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_533),
.Y(n_1458)
);

CKINVDCx20_ASAP7_75t_R g1459 ( 
.A(n_235),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_54),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_637),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_346),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_553),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_311),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_216),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_601),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_138),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_254),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_907),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_158),
.Y(n_1470)
);

CKINVDCx16_ASAP7_75t_R g1471 ( 
.A(n_359),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_438),
.Y(n_1472)
);

BUFx6f_ASAP7_75t_L g1473 ( 
.A(n_602),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_180),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_121),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_523),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_916),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_709),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_464),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_76),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_981),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_195),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_686),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_966),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_587),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_466),
.Y(n_1486)
);

INVxp33_ASAP7_75t_L g1487 ( 
.A(n_423),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_91),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_929),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_598),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_62),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_616),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_950),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_604),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_172),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_723),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_593),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_920),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_605),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_680),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_918),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_721),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_408),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_8),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_458),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_980),
.Y(n_1506)
);

BUFx10_ASAP7_75t_L g1507 ( 
.A(n_434),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_641),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_264),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_766),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_142),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_82),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_413),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_157),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_356),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_139),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_254),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_740),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_727),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1161),
.B(n_0),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1024),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1264),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1035),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1051),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1057),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1171),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1048),
.Y(n_1527)
);

INVxp67_ASAP7_75t_SL g1528 ( 
.A(n_1296),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1020),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_R g1530 ( 
.A(n_1080),
.B(n_1008),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_L g1531 ( 
.A(n_1119),
.B(n_1),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1171),
.Y(n_1532)
);

NOR2xp67_ASAP7_75t_L g1533 ( 
.A(n_1119),
.B(n_1),
.Y(n_1533)
);

INVxp33_ASAP7_75t_L g1534 ( 
.A(n_1353),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1049),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1171),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_1044),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1496),
.B(n_3),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1171),
.Y(n_1539)
);

INVxp33_ASAP7_75t_SL g1540 ( 
.A(n_1367),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1171),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1063),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1062),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1066),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1243),
.B(n_2),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1111),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1070),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1113),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1141),
.B(n_3),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1420),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1420),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1128),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1420),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1079),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1420),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1081),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1051),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1376),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_L g1559 ( 
.A(n_1439),
.B(n_4),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1056),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1137),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1420),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1028),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1052),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_L g1565 ( 
.A(n_1263),
.B(n_2),
.Y(n_1565)
);

INVxp33_ASAP7_75t_SL g1566 ( 
.A(n_1013),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1082),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1052),
.Y(n_1568)
);

INVxp33_ASAP7_75t_SL g1569 ( 
.A(n_1016),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1276),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1052),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1132),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1083),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1085),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1346),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1250),
.Y(n_1576)
);

NOR2xp67_ASAP7_75t_L g1577 ( 
.A(n_1328),
.B(n_4),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1132),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1442),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1487),
.B(n_7),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1132),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1090),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1092),
.Y(n_1583)
);

CKINVDCx5p33_ASAP7_75t_R g1584 ( 
.A(n_1097),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1300),
.Y(n_1585)
);

INVxp67_ASAP7_75t_L g1586 ( 
.A(n_1056),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1383),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1017),
.Y(n_1588)
);

CKINVDCx20_ASAP7_75t_R g1589 ( 
.A(n_1441),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1317),
.B(n_5),
.Y(n_1590)
);

INVxp67_ASAP7_75t_SL g1591 ( 
.A(n_1203),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1099),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1086),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1378),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1118),
.Y(n_1595)
);

BUFx6f_ASAP7_75t_L g1596 ( 
.A(n_1564),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1591),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1568),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1521),
.B(n_1390),
.Y(n_1599)
);

AND2x4_ASAP7_75t_L g1600 ( 
.A(n_1524),
.B(n_1014),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1523),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1571),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1525),
.Y(n_1603)
);

INVxp67_ASAP7_75t_L g1604 ( 
.A(n_1570),
.Y(n_1604)
);

INVx3_ASAP7_75t_L g1605 ( 
.A(n_1572),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1593),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1527),
.B(n_1067),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1535),
.B(n_1206),
.Y(n_1609)
);

INVxp67_ASAP7_75t_L g1610 ( 
.A(n_1563),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1581),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1557),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1526),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1532),
.Y(n_1614)
);

CKINVDCx11_ASAP7_75t_R g1615 ( 
.A(n_1529),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1542),
.B(n_1575),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1536),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1588),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1543),
.B(n_1324),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1539),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1541),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1588),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1550),
.Y(n_1623)
);

NAND2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1520),
.B(n_1203),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_1530),
.B(n_1545),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1551),
.Y(n_1626)
);

AND2x6_ASAP7_75t_L g1627 ( 
.A(n_1553),
.B(n_1219),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1555),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1547),
.B(n_1449),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1562),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1579),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1531),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1590),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1554),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1566),
.B(n_1050),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1533),
.A2(n_1519),
.B(n_1023),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1549),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1559),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1528),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1565),
.Y(n_1640)
);

OA21x2_ASAP7_75t_L g1641 ( 
.A1(n_1538),
.A2(n_1031),
.B(n_1015),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1577),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1556),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1567),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1573),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1560),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1594),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1574),
.Y(n_1648)
);

AND2x6_ASAP7_75t_L g1649 ( 
.A(n_1580),
.B(n_1219),
.Y(n_1649)
);

HB1xp67_ASAP7_75t_L g1650 ( 
.A(n_1586),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1582),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1583),
.Y(n_1652)
);

NAND2xp33_ASAP7_75t_SL g1653 ( 
.A(n_1534),
.B(n_1203),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1584),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1569),
.B(n_1384),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1592),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1522),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1558),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1600),
.B(n_1540),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1616),
.B(n_1139),
.Y(n_1660)
);

INVx4_ASAP7_75t_SL g1661 ( 
.A(n_1654),
.Y(n_1661)
);

AOI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1637),
.A2(n_1417),
.B1(n_1448),
.B2(n_1237),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1613),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1208),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1614),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1617),
.Y(n_1666)
);

INVx4_ASAP7_75t_L g1667 ( 
.A(n_1601),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1620),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1631),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1595),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1596),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1609),
.B(n_1537),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1621),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1632),
.B(n_1131),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1596),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1598),
.Y(n_1676)
);

AND2x6_ASAP7_75t_L g1677 ( 
.A(n_1638),
.B(n_1219),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1605),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1635),
.B(n_1471),
.Y(n_1679)
);

INVx4_ASAP7_75t_L g1680 ( 
.A(n_1645),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_SL g1681 ( 
.A(n_1603),
.B(n_1544),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1602),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1623),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1626),
.Y(n_1684)
);

INVx4_ASAP7_75t_L g1685 ( 
.A(n_1634),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1657),
.B(n_1019),
.C(n_1018),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1630),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1636),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1649),
.B(n_1266),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1606),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1628),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1639),
.B(n_1212),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1610),
.B(n_1118),
.Y(n_1693)
);

BUFx3_ASAP7_75t_L g1694 ( 
.A(n_1597),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1611),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1640),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1641),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1633),
.Y(n_1698)
);

INVx3_ASAP7_75t_L g1699 ( 
.A(n_1642),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1658),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1619),
.Y(n_1701)
);

BUFx6f_ASAP7_75t_L g1702 ( 
.A(n_1627),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1629),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1644),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1618),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1627),
.Y(n_1706)
);

BUFx8_ASAP7_75t_SL g1707 ( 
.A(n_1607),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1627),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1604),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1643),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1622),
.B(n_1612),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1646),
.B(n_1075),
.Y(n_1712)
);

NAND2xp33_ASAP7_75t_L g1713 ( 
.A(n_1649),
.B(n_1599),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1649),
.B(n_1489),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1648),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1624),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1647),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1650),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1651),
.Y(n_1719)
);

INVx4_ASAP7_75t_SL g1720 ( 
.A(n_1652),
.Y(n_1720)
);

INVx4_ASAP7_75t_L g1721 ( 
.A(n_1615),
.Y(n_1721)
);

BUFx6f_ASAP7_75t_L g1722 ( 
.A(n_1656),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1625),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1655),
.Y(n_1724)
);

BUFx4f_ASAP7_75t_L g1725 ( 
.A(n_1653),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1637),
.A2(n_1417),
.B1(n_1448),
.B2(n_1237),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1608),
.B(n_1546),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1613),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1596),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1613),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1616),
.B(n_1338),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1616),
.B(n_1502),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1608),
.B(n_1548),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1613),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1661),
.B(n_1552),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1701),
.B(n_1426),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1703),
.B(n_1723),
.Y(n_1737)
);

CKINVDCx20_ASAP7_75t_R g1738 ( 
.A(n_1707),
.Y(n_1738)
);

AO22x2_ASAP7_75t_L g1739 ( 
.A1(n_1679),
.A2(n_1362),
.B1(n_1156),
.B2(n_1168),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1709),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1663),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1683),
.Y(n_1742)
);

BUFx8_ASAP7_75t_L g1743 ( 
.A(n_1717),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1665),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1687),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1713),
.A2(n_1576),
.B1(n_1585),
.B2(n_1561),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1676),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1670),
.A2(n_1589),
.B1(n_1587),
.B2(n_1107),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1671),
.B(n_1147),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1666),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1668),
.Y(n_1751)
);

OR2x6_ASAP7_75t_L g1752 ( 
.A(n_1721),
.B(n_1152),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1724),
.A2(n_1115),
.B1(n_1120),
.B2(n_1100),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1673),
.Y(n_1754)
);

INVxp67_ASAP7_75t_L g1755 ( 
.A(n_1712),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1691),
.Y(n_1756)
);

BUFx8_ASAP7_75t_L g1757 ( 
.A(n_1718),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1660),
.A2(n_1045),
.B1(n_1054),
.B2(n_1039),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1675),
.B(n_1158),
.Y(n_1759)
);

AO22x2_ASAP7_75t_L g1760 ( 
.A1(n_1659),
.A2(n_1394),
.B1(n_1189),
.B2(n_1255),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1728),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1711),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1730),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1734),
.Y(n_1764)
);

OR2x6_ASAP7_75t_L g1765 ( 
.A(n_1667),
.B(n_1306),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1698),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1731),
.B(n_1338),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_1672),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1669),
.B(n_1055),
.Y(n_1769)
);

NAND2x1p5_ASAP7_75t_L g1770 ( 
.A(n_1680),
.B(n_1068),
.Y(n_1770)
);

AO22x2_ASAP7_75t_L g1771 ( 
.A1(n_1705),
.A2(n_1409),
.B1(n_1108),
.B2(n_1391),
.Y(n_1771)
);

OAI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1732),
.A2(n_1444),
.B1(n_1467),
.B2(n_1290),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1704),
.B(n_1021),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1699),
.B(n_1072),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1727),
.B(n_1022),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1682),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1694),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1700),
.B(n_1321),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1696),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1695),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1733),
.A2(n_1123),
.B1(n_1129),
.B2(n_1121),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1678),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1690),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1729),
.B(n_1368),
.Y(n_1784)
);

AO22x2_ASAP7_75t_L g1785 ( 
.A1(n_1693),
.A2(n_1096),
.B1(n_1138),
.B2(n_1065),
.Y(n_1785)
);

CKINVDCx20_ASAP7_75t_R g1786 ( 
.A(n_1720),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1674),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1664),
.B(n_1398),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1684),
.Y(n_1789)
);

INVx2_ASAP7_75t_L g1790 ( 
.A(n_1684),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1722),
.B(n_1398),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1716),
.Y(n_1792)
);

CKINVDCx5p33_ASAP7_75t_R g1793 ( 
.A(n_1722),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1710),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1715),
.B(n_1076),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1719),
.Y(n_1796)
);

AO22x2_ASAP7_75t_L g1797 ( 
.A1(n_1692),
.A2(n_1114),
.B1(n_1175),
.B2(n_1088),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1697),
.B(n_1089),
.Y(n_1798)
);

AO22x2_ASAP7_75t_L g1799 ( 
.A1(n_1686),
.A2(n_1122),
.B1(n_1385),
.B2(n_1091),
.Y(n_1799)
);

AND2x4_ASAP7_75t_L g1800 ( 
.A(n_1685),
.B(n_1708),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1706),
.B(n_1377),
.Y(n_1801)
);

CKINVDCx20_ASAP7_75t_R g1802 ( 
.A(n_1725),
.Y(n_1802)
);

AND2x2_ASAP7_75t_SL g1803 ( 
.A(n_1681),
.B(n_1237),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1689),
.B(n_1095),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1688),
.Y(n_1805)
);

AO22x2_ASAP7_75t_L g1806 ( 
.A1(n_1714),
.A2(n_1254),
.B1(n_1274),
.B2(n_1218),
.Y(n_1806)
);

AO22x2_ASAP7_75t_L g1807 ( 
.A1(n_1662),
.A2(n_1246),
.B1(n_1268),
.B2(n_1220),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1702),
.B(n_1405),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1688),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1726),
.B(n_1408),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1677),
.Y(n_1811)
);

INVx2_ASAP7_75t_SL g1812 ( 
.A(n_1677),
.Y(n_1812)
);

AO22x2_ASAP7_75t_L g1813 ( 
.A1(n_1677),
.A2(n_1299),
.B1(n_1329),
.B2(n_1229),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1702),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1663),
.Y(n_1815)
);

NOR2x1p5_ASAP7_75t_L g1816 ( 
.A(n_1667),
.B(n_1446),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1663),
.Y(n_1817)
);

HB1xp67_ASAP7_75t_L g1818 ( 
.A(n_1709),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1670),
.B(n_1025),
.Y(n_1819)
);

AO22x2_ASAP7_75t_L g1820 ( 
.A1(n_1679),
.A2(n_1036),
.B1(n_1424),
.B2(n_1406),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1670),
.B(n_1026),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1663),
.Y(n_1822)
);

INVxp67_ASAP7_75t_L g1823 ( 
.A(n_1670),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1709),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1701),
.B(n_1102),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1663),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1663),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1701),
.B(n_1112),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1663),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1670),
.Y(n_1830)
);

AO22x2_ASAP7_75t_L g1831 ( 
.A1(n_1679),
.A2(n_1226),
.B1(n_1269),
.B2(n_1074),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1670),
.B(n_1029),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1663),
.Y(n_1833)
);

INVxp67_ASAP7_75t_SL g1834 ( 
.A(n_1684),
.Y(n_1834)
);

NAND2x1p5_ASAP7_75t_L g1835 ( 
.A(n_1680),
.B(n_1126),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1663),
.Y(n_1836)
);

AO22x2_ASAP7_75t_L g1837 ( 
.A1(n_1679),
.A2(n_1078),
.B1(n_1323),
.B2(n_1059),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1663),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1701),
.B(n_1133),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1711),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1701),
.B(n_1143),
.Y(n_1841)
);

OR2x6_ASAP7_75t_L g1842 ( 
.A(n_1717),
.B(n_1504),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1731),
.B(n_1408),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1701),
.B(n_1146),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1731),
.B(n_1507),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_SL g1846 ( 
.A(n_1722),
.B(n_1518),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1670),
.B(n_1030),
.Y(n_1847)
);

AO22x2_ASAP7_75t_L g1848 ( 
.A1(n_1679),
.A2(n_1134),
.B1(n_1160),
.B2(n_1061),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1660),
.A2(n_1201),
.B1(n_1202),
.B2(n_1197),
.C(n_1155),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1663),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_SL g1851 ( 
.A(n_1722),
.B(n_1506),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1663),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1683),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1663),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1731),
.B(n_1507),
.Y(n_1855)
);

AO22x2_ASAP7_75t_L g1856 ( 
.A1(n_1679),
.A2(n_1319),
.B1(n_1370),
.B2(n_1247),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1663),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1663),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1663),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1723),
.A2(n_1142),
.B1(n_1144),
.B2(n_1130),
.Y(n_1860)
);

AO22x2_ASAP7_75t_L g1861 ( 
.A1(n_1679),
.A2(n_1423),
.B1(n_1327),
.B2(n_1241),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1663),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1711),
.Y(n_1863)
);

OR2x2_ASAP7_75t_SL g1864 ( 
.A(n_1724),
.B(n_1058),
.Y(n_1864)
);

AO22x2_ASAP7_75t_L g1865 ( 
.A1(n_1679),
.A2(n_1207),
.B1(n_1336),
.B2(n_1288),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1663),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1701),
.B(n_1148),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1717),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1663),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1723),
.A2(n_1153),
.B1(n_1163),
.B2(n_1150),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1683),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1663),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1717),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1663),
.Y(n_1874)
);

INVxp67_ASAP7_75t_L g1875 ( 
.A(n_1670),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1663),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1793),
.B(n_1167),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_SL g1878 ( 
.A(n_1803),
.B(n_1840),
.Y(n_1878)
);

NAND2xp33_ASAP7_75t_SL g1879 ( 
.A(n_1802),
.B(n_1027),
.Y(n_1879)
);

NAND2xp33_ASAP7_75t_SL g1880 ( 
.A(n_1786),
.B(n_1106),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1863),
.B(n_1172),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1823),
.B(n_1176),
.Y(n_1882)
);

NAND2xp33_ASAP7_75t_SL g1883 ( 
.A(n_1816),
.B(n_1135),
.Y(n_1883)
);

NAND2xp33_ASAP7_75t_SL g1884 ( 
.A(n_1768),
.B(n_1136),
.Y(n_1884)
);

NAND2xp33_ASAP7_75t_SL g1885 ( 
.A(n_1767),
.B(n_1157),
.Y(n_1885)
);

NAND2xp33_ASAP7_75t_SL g1886 ( 
.A(n_1843),
.B(n_1165),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1830),
.B(n_1180),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_SL g1888 ( 
.A(n_1875),
.B(n_1182),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1737),
.B(n_1184),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1819),
.B(n_1821),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1832),
.B(n_1185),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1847),
.B(n_1186),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_SL g1893 ( 
.A(n_1736),
.B(n_1187),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_SL g1894 ( 
.A(n_1775),
.B(n_1190),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1762),
.B(n_1216),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1791),
.B(n_1225),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1755),
.B(n_1242),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_SL g1898 ( 
.A(n_1777),
.B(n_1252),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1845),
.B(n_1259),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_SL g1900 ( 
.A(n_1855),
.B(n_1267),
.Y(n_1900)
);

NAND2xp33_ASAP7_75t_SL g1901 ( 
.A(n_1814),
.B(n_1230),
.Y(n_1901)
);

NAND2xp33_ASAP7_75t_SL g1902 ( 
.A(n_1788),
.B(n_1812),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_SL g1903 ( 
.A(n_1800),
.B(n_1271),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1834),
.B(n_1339),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1825),
.B(n_1272),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1828),
.B(n_1284),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_SL g1907 ( 
.A(n_1839),
.B(n_1286),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1740),
.B(n_1032),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1841),
.B(n_1292),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1844),
.B(n_1293),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1867),
.B(n_1301),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1818),
.B(n_1356),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1796),
.B(n_1304),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_SL g1914 ( 
.A(n_1794),
.B(n_1310),
.Y(n_1914)
);

NAND2xp33_ASAP7_75t_SL g1915 ( 
.A(n_1810),
.B(n_1374),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1792),
.B(n_1177),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1824),
.B(n_1033),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1748),
.B(n_1034),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1741),
.B(n_1178),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1744),
.B(n_1312),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_SL g1921 ( 
.A(n_1750),
.B(n_1315),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1751),
.B(n_1316),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1754),
.B(n_1756),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1761),
.B(n_1326),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1763),
.B(n_1330),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1764),
.B(n_1340),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_SL g1927 ( 
.A(n_1815),
.B(n_1342),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_SL g1928 ( 
.A(n_1811),
.B(n_1382),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1817),
.B(n_1343),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1822),
.B(n_1348),
.Y(n_1930)
);

NAND2xp33_ASAP7_75t_SL g1931 ( 
.A(n_1735),
.B(n_1389),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1826),
.B(n_1355),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1827),
.B(n_1829),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1833),
.B(n_1181),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1790),
.B(n_1352),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1836),
.B(n_1365),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1838),
.B(n_1371),
.Y(n_1937)
);

NAND2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1787),
.B(n_1459),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1850),
.B(n_1372),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1852),
.B(n_1373),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1854),
.B(n_1388),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1857),
.B(n_1400),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1858),
.B(n_1402),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1859),
.B(n_1407),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1862),
.B(n_1415),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1866),
.B(n_1869),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1872),
.B(n_1191),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_SL g1948 ( 
.A(n_1874),
.B(n_1419),
.Y(n_1948)
);

NAND2xp33_ASAP7_75t_SL g1949 ( 
.A(n_1846),
.B(n_1480),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1876),
.B(n_1431),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1860),
.B(n_1435),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1870),
.B(n_1436),
.Y(n_1952)
);

NAND2xp33_ASAP7_75t_SL g1953 ( 
.A(n_1851),
.B(n_1779),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1753),
.B(n_1450),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1746),
.B(n_1469),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1789),
.B(n_1361),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1804),
.B(n_1781),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1782),
.B(n_1395),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1783),
.B(n_1397),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1868),
.B(n_1037),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_SL g1961 ( 
.A(n_1778),
.B(n_1477),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1766),
.B(n_1478),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1776),
.B(n_1481),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1780),
.B(n_1483),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1773),
.B(n_1484),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_SL g1966 ( 
.A(n_1772),
.B(n_1493),
.Y(n_1966)
);

NAND2xp33_ASAP7_75t_SL g1967 ( 
.A(n_1795),
.B(n_1500),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1873),
.B(n_1038),
.Y(n_1968)
);

NAND2xp33_ASAP7_75t_SL g1969 ( 
.A(n_1808),
.B(n_1501),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1774),
.B(n_1212),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1742),
.B(n_1337),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1769),
.B(n_1193),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1745),
.B(n_1337),
.Y(n_1973)
);

NAND2xp33_ASAP7_75t_SL g1974 ( 
.A(n_1758),
.B(n_1040),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1747),
.B(n_1253),
.Y(n_1975)
);

NAND2xp33_ASAP7_75t_SL g1976 ( 
.A(n_1805),
.B(n_1041),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1853),
.B(n_1871),
.Y(n_1977)
);

NAND2xp33_ASAP7_75t_SL g1978 ( 
.A(n_1809),
.B(n_1043),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1770),
.B(n_1253),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1835),
.B(n_1253),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_SL g1981 ( 
.A(n_1801),
.B(n_1412),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1749),
.B(n_1759),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1798),
.B(n_1205),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1784),
.B(n_1412),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1743),
.B(n_1412),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1820),
.B(n_1211),
.Y(n_1986)
);

AND2x2_ASAP7_75t_SL g1987 ( 
.A(n_1757),
.B(n_1417),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1831),
.B(n_1213),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_SL g1989 ( 
.A(n_1837),
.B(n_1214),
.Y(n_1989)
);

NAND2xp33_ASAP7_75t_SL g1990 ( 
.A(n_1738),
.B(n_1046),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1848),
.B(n_1215),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1856),
.B(n_1221),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1861),
.B(n_1232),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1865),
.B(n_1235),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1739),
.B(n_1239),
.Y(n_1995)
);

NAND2xp33_ASAP7_75t_SL g1996 ( 
.A(n_1864),
.B(n_1047),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1797),
.B(n_1248),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1799),
.B(n_1285),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1807),
.B(n_1287),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1760),
.B(n_1294),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_SL g2001 ( 
.A(n_1785),
.B(n_1307),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1806),
.B(n_1053),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1765),
.B(n_1325),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1765),
.B(n_1335),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_SL g2005 ( 
.A(n_1813),
.B(n_1060),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_SL g2006 ( 
.A(n_1842),
.B(n_1341),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1842),
.B(n_1354),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1752),
.B(n_1399),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1849),
.B(n_1358),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1771),
.B(n_1363),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1752),
.B(n_1366),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1793),
.B(n_1369),
.Y(n_2012)
);

NAND2xp33_ASAP7_75t_SL g2013 ( 
.A(n_1793),
.B(n_1064),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1793),
.B(n_1401),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1737),
.B(n_1428),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1737),
.B(n_1440),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1793),
.B(n_1451),
.Y(n_2017)
);

NAND2xp33_ASAP7_75t_SL g2018 ( 
.A(n_1793),
.B(n_1069),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1793),
.B(n_1455),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1793),
.B(n_1498),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1793),
.B(n_1510),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1737),
.B(n_1042),
.Y(n_2022)
);

NAND2xp33_ASAP7_75t_SL g2023 ( 
.A(n_1793),
.B(n_1071),
.Y(n_2023)
);

NAND2xp33_ASAP7_75t_SL g2024 ( 
.A(n_1793),
.B(n_1073),
.Y(n_2024)
);

NAND2xp33_ASAP7_75t_SL g2025 ( 
.A(n_1793),
.B(n_1077),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1793),
.B(n_1042),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_SL g2027 ( 
.A(n_1793),
.B(n_1042),
.Y(n_2027)
);

NAND2xp33_ASAP7_75t_SL g2028 ( 
.A(n_1793),
.B(n_1084),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1793),
.B(n_1042),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1793),
.B(n_1042),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1793),
.B(n_1195),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1793),
.B(n_1195),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_SL g2033 ( 
.A(n_1793),
.B(n_1195),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1793),
.B(n_1195),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1793),
.B(n_1195),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_SL g2036 ( 
.A(n_1793),
.B(n_1448),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1823),
.B(n_1087),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_SL g2038 ( 
.A(n_1793),
.B(n_1093),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1793),
.B(n_1462),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_1793),
.B(n_1462),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1793),
.B(n_1462),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1793),
.B(n_1473),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1793),
.B(n_1473),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1793),
.B(n_1473),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_SL g2045 ( 
.A(n_1793),
.B(n_1094),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1834),
.B(n_1427),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1793),
.B(n_1101),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1823),
.B(n_1103),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1793),
.B(n_1104),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_SL g2050 ( 
.A(n_1793),
.B(n_1105),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1793),
.B(n_1109),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1737),
.B(n_1110),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1793),
.B(n_1116),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1793),
.B(n_1117),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1793),
.B(n_1124),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1793),
.B(n_1125),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_SL g2057 ( 
.A(n_1793),
.B(n_1140),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1793),
.B(n_1145),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1834),
.B(n_1434),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1823),
.B(n_1149),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1834),
.B(n_1438),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1737),
.B(n_1151),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1793),
.B(n_1154),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1793),
.B(n_1159),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_SL g2065 ( 
.A(n_1793),
.B(n_1162),
.Y(n_2065)
);

NAND2xp33_ASAP7_75t_SL g2066 ( 
.A(n_1793),
.B(n_1164),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_SL g2067 ( 
.A(n_1793),
.B(n_1166),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1793),
.B(n_1169),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1793),
.B(n_1170),
.Y(n_2069)
);

NAND2xp33_ASAP7_75t_SL g2070 ( 
.A(n_1793),
.B(n_1173),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_1793),
.B(n_1174),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1823),
.B(n_1179),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1793),
.B(n_1183),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_SL g2074 ( 
.A(n_1793),
.B(n_1188),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1793),
.B(n_1192),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_1823),
.B(n_1194),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_1823),
.B(n_1196),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1890),
.B(n_1198),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1935),
.Y(n_2079)
);

HB1xp67_ASAP7_75t_L g2080 ( 
.A(n_1904),
.Y(n_2080)
);

AOI21x1_ASAP7_75t_SL g2081 ( 
.A1(n_1986),
.A2(n_1200),
.B(n_1199),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2052),
.B(n_1204),
.Y(n_2082)
);

BUFx12f_ASAP7_75t_L g2083 ( 
.A(n_2008),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1956),
.Y(n_2084)
);

OR2x2_ASAP7_75t_L g2085 ( 
.A(n_1884),
.B(n_1209),
.Y(n_2085)
);

OR2x2_ASAP7_75t_L g2086 ( 
.A(n_2062),
.B(n_1210),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2037),
.B(n_1217),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_SL g2088 ( 
.A(n_1987),
.B(n_1512),
.Y(n_2088)
);

AOI22xp5_ASAP7_75t_L g2089 ( 
.A1(n_1878),
.A2(n_1223),
.B1(n_1224),
.B2(n_1222),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2048),
.B(n_1228),
.Y(n_2090)
);

INVxp67_ASAP7_75t_SL g2091 ( 
.A(n_1923),
.Y(n_2091)
);

AOI21x1_ASAP7_75t_SL g2092 ( 
.A1(n_1988),
.A2(n_1233),
.B(n_1231),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1935),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1958),
.Y(n_2094)
);

OAI22x1_ASAP7_75t_L g2095 ( 
.A1(n_1918),
.A2(n_1236),
.B1(n_1238),
.B2(n_1234),
.Y(n_2095)
);

CKINVDCx5p33_ASAP7_75t_R g2096 ( 
.A(n_1990),
.Y(n_2096)
);

NAND3xp33_ASAP7_75t_SL g2097 ( 
.A(n_2065),
.B(n_1244),
.C(n_1240),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_2022),
.A2(n_1466),
.B(n_1454),
.Y(n_2098)
);

BUFx2_ASAP7_75t_L g2099 ( 
.A(n_1879),
.Y(n_2099)
);

INVx2_ASAP7_75t_SL g2100 ( 
.A(n_1960),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1958),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1977),
.A2(n_1482),
.B(n_1127),
.Y(n_2102)
);

CKINVDCx5p33_ASAP7_75t_R g2103 ( 
.A(n_1880),
.Y(n_2103)
);

A2O1A1Ixp33_ASAP7_75t_L g2104 ( 
.A1(n_1957),
.A2(n_1227),
.B(n_1318),
.C(n_1098),
.Y(n_2104)
);

OAI22xp5_ASAP7_75t_L g2105 ( 
.A1(n_2015),
.A2(n_1249),
.B1(n_1251),
.B2(n_1245),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_1983),
.A2(n_1331),
.B(n_1322),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1959),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_1933),
.A2(n_1946),
.B(n_1934),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_1919),
.A2(n_1393),
.B(n_1387),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2016),
.B(n_1256),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2060),
.B(n_1257),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_1912),
.B(n_1258),
.Y(n_2112)
);

OAI21x1_ASAP7_75t_L g2113 ( 
.A1(n_1947),
.A2(n_1432),
.B(n_1422),
.Y(n_2113)
);

BUFx6f_ASAP7_75t_L g2114 ( 
.A(n_1956),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_1982),
.B(n_1453),
.Y(n_2115)
);

OAI21xp5_ASAP7_75t_L g2116 ( 
.A1(n_1972),
.A2(n_1503),
.B(n_1490),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1953),
.A2(n_645),
.B(n_644),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_SL g2118 ( 
.A1(n_1999),
.A2(n_649),
.B(n_646),
.Y(n_2118)
);

BUFx3_ASAP7_75t_L g2119 ( 
.A(n_1959),
.Y(n_2119)
);

OAI21x1_ASAP7_75t_L g2120 ( 
.A1(n_1916),
.A2(n_1963),
.B(n_1964),
.Y(n_2120)
);

AOI21xp33_ASAP7_75t_L g2121 ( 
.A1(n_1891),
.A2(n_1261),
.B(n_1260),
.Y(n_2121)
);

OR2x2_ASAP7_75t_L g2122 ( 
.A(n_2072),
.B(n_1262),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2076),
.B(n_1265),
.Y(n_2123)
);

OAI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_1892),
.A2(n_1273),
.B(n_1270),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2077),
.B(n_1275),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_1915),
.A2(n_1278),
.B1(n_1279),
.B2(n_1277),
.Y(n_2126)
);

OAI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1889),
.A2(n_1894),
.B(n_1893),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_1903),
.A2(n_651),
.B(n_650),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1904),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_1968),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2046),
.B(n_1280),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1881),
.A2(n_654),
.B(n_652),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_1962),
.A2(n_659),
.B(n_658),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2046),
.B(n_1281),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2059),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_1914),
.A2(n_661),
.B(n_660),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2059),
.B(n_1282),
.Y(n_2137)
);

OAI21x1_ASAP7_75t_L g2138 ( 
.A1(n_1920),
.A2(n_663),
.B(n_662),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_2061),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2061),
.Y(n_2140)
);

AO31x2_ASAP7_75t_L g2141 ( 
.A1(n_1995),
.A2(n_667),
.A3(n_668),
.B(n_665),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_1908),
.B(n_670),
.Y(n_2142)
);

O2A1O1Ixp5_ASAP7_75t_L g2143 ( 
.A1(n_1965),
.A2(n_1906),
.B(n_1907),
.C(n_1905),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1882),
.B(n_1283),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1998),
.Y(n_2145)
);

A2O1A1Ixp33_ASAP7_75t_L g2146 ( 
.A1(n_1949),
.A2(n_1291),
.B(n_1295),
.C(n_1289),
.Y(n_2146)
);

AOI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_1921),
.A2(n_672),
.B(n_671),
.Y(n_2147)
);

CKINVDCx5p33_ASAP7_75t_R g2148 ( 
.A(n_1931),
.Y(n_2148)
);

NAND2xp33_ASAP7_75t_R g2149 ( 
.A(n_1917),
.B(n_673),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1989),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2045),
.B(n_1297),
.Y(n_2151)
);

INVx1_ASAP7_75t_SL g2152 ( 
.A(n_2013),
.Y(n_2152)
);

OAI21x1_ASAP7_75t_L g2153 ( 
.A1(n_1922),
.A2(n_675),
.B(n_674),
.Y(n_2153)
);

AO21x2_ASAP7_75t_L g2154 ( 
.A1(n_1909),
.A2(n_679),
.B(n_677),
.Y(n_2154)
);

AOI31xp67_ASAP7_75t_L g2155 ( 
.A1(n_2000),
.A2(n_682),
.A3(n_683),
.B(n_681),
.Y(n_2155)
);

AOI21x1_ASAP7_75t_L g2156 ( 
.A1(n_1910),
.A2(n_690),
.B(n_687),
.Y(n_2156)
);

INVx3_ASAP7_75t_L g2157 ( 
.A(n_2008),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_SL g2158 ( 
.A(n_1885),
.B(n_1298),
.Y(n_2158)
);

AOI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_1924),
.A2(n_693),
.B(n_692),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_2006),
.Y(n_2160)
);

A2O1A1Ixp33_ASAP7_75t_L g2161 ( 
.A1(n_1928),
.A2(n_1303),
.B(n_1305),
.C(n_1302),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1887),
.B(n_1308),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_1886),
.A2(n_1901),
.B(n_1902),
.C(n_1974),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_1896),
.B(n_694),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1925),
.A2(n_701),
.B(n_696),
.Y(n_2165)
);

NAND3x1_ASAP7_75t_L g2166 ( 
.A(n_1883),
.B(n_1311),
.C(n_1309),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1975),
.Y(n_2167)
);

O2A1O1Ixp5_ASAP7_75t_SL g2168 ( 
.A1(n_2010),
.A2(n_1509),
.B(n_1511),
.C(n_1508),
.Y(n_2168)
);

OAI21xp33_ASAP7_75t_L g2169 ( 
.A1(n_1888),
.A2(n_1314),
.B(n_1313),
.Y(n_2169)
);

INVx2_ASAP7_75t_SL g2170 ( 
.A(n_2047),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1991),
.Y(n_2171)
);

AOI21xp5_ASAP7_75t_L g2172 ( 
.A1(n_1926),
.A2(n_704),
.B(n_703),
.Y(n_2172)
);

NAND3xp33_ASAP7_75t_L g2173 ( 
.A(n_1966),
.B(n_1332),
.C(n_1320),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1899),
.B(n_1333),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_1900),
.A2(n_1344),
.B1(n_1345),
.B2(n_1334),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2049),
.B(n_1347),
.Y(n_2176)
);

NOR2x1_ASAP7_75t_SL g2177 ( 
.A(n_2026),
.B(n_705),
.Y(n_2177)
);

A2O1A1Ixp33_ASAP7_75t_L g2178 ( 
.A1(n_1976),
.A2(n_1350),
.B(n_1351),
.C(n_1349),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_1938),
.B(n_1357),
.Y(n_2179)
);

NOR2xp67_ASAP7_75t_L g2180 ( 
.A(n_1877),
.B(n_706),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_L g2181 ( 
.A1(n_1927),
.A2(n_710),
.B(n_707),
.Y(n_2181)
);

BUFx6f_ASAP7_75t_L g2182 ( 
.A(n_2007),
.Y(n_2182)
);

AO31x2_ASAP7_75t_L g2183 ( 
.A1(n_1992),
.A2(n_712),
.A3(n_713),
.B(n_711),
.Y(n_2183)
);

NAND3xp33_ASAP7_75t_L g2184 ( 
.A(n_2018),
.B(n_1360),
.C(n_1359),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1993),
.Y(n_2185)
);

AO21x1_ASAP7_75t_L g2186 ( 
.A1(n_1994),
.A2(n_5),
.B(n_8),
.Y(n_2186)
);

NAND2x1p5_ASAP7_75t_L g2187 ( 
.A(n_2003),
.B(n_714),
.Y(n_2187)
);

INVx8_ASAP7_75t_L g2188 ( 
.A(n_1969),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_1897),
.B(n_1364),
.Y(n_2189)
);

INVx4_ASAP7_75t_L g2190 ( 
.A(n_2023),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_1929),
.A2(n_1932),
.B(n_1930),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1911),
.B(n_1936),
.Y(n_2192)
);

OR2x6_ASAP7_75t_L g2193 ( 
.A(n_2011),
.B(n_9),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1997),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1981),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_1937),
.A2(n_1940),
.B(n_1939),
.Y(n_2196)
);

AO31x2_ASAP7_75t_L g2197 ( 
.A1(n_2002),
.A2(n_716),
.A3(n_717),
.B(n_715),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2001),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1984),
.Y(n_2199)
);

BUFx2_ASAP7_75t_L g2200 ( 
.A(n_1978),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2027),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_1941),
.A2(n_720),
.B(n_718),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_L g2203 ( 
.A1(n_1942),
.A2(n_725),
.B(n_722),
.Y(n_2203)
);

NOR4xp25_ASAP7_75t_L g2204 ( 
.A(n_2009),
.B(n_1379),
.C(n_1380),
.D(n_1375),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1943),
.B(n_1944),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_1945),
.A2(n_729),
.B(n_728),
.Y(n_2206)
);

OAI21x1_ASAP7_75t_L g2207 ( 
.A1(n_1948),
.A2(n_731),
.B(n_730),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_2024),
.Y(n_2208)
);

AOI21x1_ASAP7_75t_L g2209 ( 
.A1(n_1950),
.A2(n_1898),
.B(n_2029),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2030),
.B(n_1381),
.Y(n_2210)
);

O2A1O1Ixp33_ASAP7_75t_SL g2211 ( 
.A1(n_1951),
.A2(n_733),
.B(n_734),
.C(n_732),
.Y(n_2211)
);

INVx2_ASAP7_75t_SL g2212 ( 
.A(n_2050),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_L g2213 ( 
.A(n_2031),
.B(n_1386),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_SL g2214 ( 
.A(n_2025),
.B(n_1392),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_2036),
.Y(n_2215)
);

OAI21x1_ASAP7_75t_L g2216 ( 
.A1(n_2032),
.A2(n_737),
.B(n_736),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_1895),
.A2(n_742),
.B(n_741),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_2012),
.B(n_744),
.Y(n_2218)
);

OAI21x1_ASAP7_75t_SL g2219 ( 
.A1(n_2033),
.A2(n_2035),
.B(n_2034),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_1913),
.A2(n_749),
.B(n_745),
.Y(n_2220)
);

AO32x2_ASAP7_75t_L g2221 ( 
.A1(n_2005),
.A2(n_11),
.A3(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1955),
.B(n_1396),
.Y(n_2222)
);

BUFx12f_ASAP7_75t_L g2223 ( 
.A(n_2028),
.Y(n_2223)
);

AOI21xp33_ASAP7_75t_L g2224 ( 
.A1(n_1952),
.A2(n_1404),
.B(n_1403),
.Y(n_2224)
);

CKINVDCx5p33_ASAP7_75t_R g2225 ( 
.A(n_2038),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2039),
.Y(n_2226)
);

INVx1_ASAP7_75t_SL g2227 ( 
.A(n_2066),
.Y(n_2227)
);

AO21x2_ASAP7_75t_L g2228 ( 
.A1(n_1954),
.A2(n_753),
.B(n_751),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2014),
.B(n_1410),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_L g2230 ( 
.A1(n_1979),
.A2(n_755),
.B(n_754),
.Y(n_2230)
);

OAI21x1_ASAP7_75t_L g2231 ( 
.A1(n_1980),
.A2(n_757),
.B(n_756),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2145),
.Y(n_2232)
);

OAI21x1_ASAP7_75t_L g2233 ( 
.A1(n_2102),
.A2(n_1970),
.B(n_2040),
.Y(n_2233)
);

AND2x2_ASAP7_75t_L g2234 ( 
.A(n_2087),
.B(n_2074),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2185),
.Y(n_2235)
);

CKINVDCx20_ASAP7_75t_R g2236 ( 
.A(n_2096),
.Y(n_2236)
);

OAI21x1_ASAP7_75t_L g2237 ( 
.A1(n_2109),
.A2(n_2042),
.B(n_2041),
.Y(n_2237)
);

OAI21x1_ASAP7_75t_L g2238 ( 
.A1(n_2113),
.A2(n_2044),
.B(n_2043),
.Y(n_2238)
);

INVx2_ASAP7_75t_SL g2239 ( 
.A(n_2083),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_2082),
.B(n_2017),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2112),
.B(n_2019),
.Y(n_2241)
);

OA21x2_ASAP7_75t_L g2242 ( 
.A1(n_2106),
.A2(n_2098),
.B(n_2108),
.Y(n_2242)
);

NAND3xp33_ASAP7_75t_L g2243 ( 
.A(n_2124),
.B(n_2071),
.C(n_2070),
.Y(n_2243)
);

OA21x2_ASAP7_75t_L g2244 ( 
.A1(n_2120),
.A2(n_2021),
.B(n_2020),
.Y(n_2244)
);

OA21x2_ASAP7_75t_L g2245 ( 
.A1(n_2191),
.A2(n_1973),
.B(n_1971),
.Y(n_2245)
);

AND2x4_ASAP7_75t_L g2246 ( 
.A(n_2119),
.B(n_2051),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_2138),
.A2(n_2054),
.B(n_2053),
.Y(n_2247)
);

NAND2x1p5_ASAP7_75t_L g2248 ( 
.A(n_2100),
.B(n_1985),
.Y(n_2248)
);

OAI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_2088),
.A2(n_2055),
.B1(n_2057),
.B2(n_2056),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2110),
.B(n_2058),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_2129),
.Y(n_2251)
);

AO31x2_ASAP7_75t_L g2252 ( 
.A1(n_2104),
.A2(n_1967),
.A3(n_1996),
.B(n_1961),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2090),
.B(n_2063),
.Y(n_2253)
);

NOR2x1_ASAP7_75t_SL g2254 ( 
.A(n_2228),
.B(n_2004),
.Y(n_2254)
);

BUFx3_ASAP7_75t_L g2255 ( 
.A(n_2130),
.Y(n_2255)
);

AOI21x1_ASAP7_75t_L g2256 ( 
.A1(n_2209),
.A2(n_2067),
.B(n_2064),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2150),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2080),
.B(n_2068),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2171),
.Y(n_2259)
);

OA21x2_ASAP7_75t_L g2260 ( 
.A1(n_2196),
.A2(n_2073),
.B(n_2069),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2194),
.Y(n_2261)
);

BUFx12f_ASAP7_75t_L g2262 ( 
.A(n_2223),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2198),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2114),
.Y(n_2264)
);

OAI21xp5_ASAP7_75t_L g2265 ( 
.A1(n_2143),
.A2(n_2168),
.B(n_2127),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2153),
.A2(n_2075),
.B(n_759),
.Y(n_2266)
);

BUFx2_ASAP7_75t_L g2267 ( 
.A(n_2114),
.Y(n_2267)
);

CKINVDCx16_ASAP7_75t_R g2268 ( 
.A(n_2149),
.Y(n_2268)
);

NAND3xp33_ASAP7_75t_L g2269 ( 
.A(n_2146),
.B(n_1413),
.C(n_1411),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2091),
.Y(n_2270)
);

NAND2x1_ASAP7_75t_L g2271 ( 
.A(n_2219),
.B(n_758),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2157),
.Y(n_2272)
);

INVx2_ASAP7_75t_SL g2273 ( 
.A(n_2160),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2079),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2093),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2107),
.Y(n_2276)
);

INVxp67_ASAP7_75t_SL g2277 ( 
.A(n_2135),
.Y(n_2277)
);

AO21x2_ASAP7_75t_L g2278 ( 
.A1(n_2118),
.A2(n_762),
.B(n_760),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2140),
.Y(n_2279)
);

AO31x2_ASAP7_75t_L g2280 ( 
.A1(n_2186),
.A2(n_767),
.A3(n_769),
.B(n_764),
.Y(n_2280)
);

INVxp67_ASAP7_75t_SL g2281 ( 
.A(n_2139),
.Y(n_2281)
);

OAI21x1_ASAP7_75t_L g2282 ( 
.A1(n_2181),
.A2(n_772),
.B(n_771),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2094),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2101),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2084),
.Y(n_2285)
);

OR2x2_ASAP7_75t_L g2286 ( 
.A(n_2122),
.B(n_2111),
.Y(n_2286)
);

NOR2xp33_ASAP7_75t_L g2287 ( 
.A(n_2086),
.B(n_2099),
.Y(n_2287)
);

INVx2_ASAP7_75t_SL g2288 ( 
.A(n_2160),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2199),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2167),
.Y(n_2290)
);

INVx4_ASAP7_75t_L g2291 ( 
.A(n_2182),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2195),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2201),
.Y(n_2293)
);

OAI21x1_ASAP7_75t_L g2294 ( 
.A1(n_2202),
.A2(n_775),
.B(n_773),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2123),
.B(n_2125),
.Y(n_2295)
);

OAI21x1_ASAP7_75t_L g2296 ( 
.A1(n_2203),
.A2(n_777),
.B(n_776),
.Y(n_2296)
);

OAI21x1_ASAP7_75t_SL g2297 ( 
.A1(n_2177),
.A2(n_779),
.B(n_778),
.Y(n_2297)
);

INVx6_ASAP7_75t_L g2298 ( 
.A(n_2182),
.Y(n_2298)
);

CKINVDCx16_ASAP7_75t_R g2299 ( 
.A(n_2085),
.Y(n_2299)
);

AO21x2_ASAP7_75t_L g2300 ( 
.A1(n_2117),
.A2(n_783),
.B(n_782),
.Y(n_2300)
);

OAI21x1_ASAP7_75t_SL g2301 ( 
.A1(n_2156),
.A2(n_787),
.B(n_784),
.Y(n_2301)
);

OAI21x1_ASAP7_75t_L g2302 ( 
.A1(n_2206),
.A2(n_789),
.B(n_788),
.Y(n_2302)
);

AND2x4_ASAP7_75t_L g2303 ( 
.A(n_2170),
.B(n_791),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2097),
.A2(n_1416),
.B1(n_1418),
.B2(n_1414),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2131),
.B(n_1421),
.Y(n_2305)
);

OAI21x1_ASAP7_75t_L g2306 ( 
.A1(n_2207),
.A2(n_793),
.B(n_792),
.Y(n_2306)
);

AOI21xp5_ASAP7_75t_SL g2307 ( 
.A1(n_2163),
.A2(n_796),
.B(n_795),
.Y(n_2307)
);

OA21x2_ASAP7_75t_L g2308 ( 
.A1(n_2133),
.A2(n_1429),
.B(n_1425),
.Y(n_2308)
);

BUFx6f_ASAP7_75t_SL g2309 ( 
.A(n_2212),
.Y(n_2309)
);

NOR2xp33_ASAP7_75t_SL g2310 ( 
.A(n_2103),
.B(n_1430),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2225),
.Y(n_2311)
);

AO21x2_ASAP7_75t_L g2312 ( 
.A1(n_2204),
.A2(n_798),
.B(n_797),
.Y(n_2312)
);

O2A1O1Ixp33_ASAP7_75t_L g2313 ( 
.A1(n_2161),
.A2(n_1437),
.B(n_1443),
.C(n_1433),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2151),
.B(n_1445),
.Y(n_2314)
);

NOR2xp67_ASAP7_75t_L g2315 ( 
.A(n_2190),
.B(n_800),
.Y(n_2315)
);

AOI31xp67_ASAP7_75t_L g2316 ( 
.A1(n_2155),
.A2(n_802),
.A3(n_803),
.B(n_801),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2226),
.Y(n_2317)
);

INVx3_ASAP7_75t_L g2318 ( 
.A(n_2215),
.Y(n_2318)
);

OAI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_2205),
.A2(n_1452),
.B(n_1447),
.Y(n_2319)
);

CKINVDCx20_ASAP7_75t_R g2320 ( 
.A(n_2148),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2216),
.Y(n_2321)
);

OR2x2_ASAP7_75t_L g2322 ( 
.A(n_2134),
.B(n_1456),
.Y(n_2322)
);

NAND2x1p5_ASAP7_75t_L g2323 ( 
.A(n_2152),
.B(n_807),
.Y(n_2323)
);

BUFx6f_ASAP7_75t_L g2324 ( 
.A(n_2215),
.Y(n_2324)
);

OAI22xp5_ASAP7_75t_L g2325 ( 
.A1(n_2192),
.A2(n_1458),
.B1(n_1460),
.B2(n_1457),
.Y(n_2325)
);

CKINVDCx20_ASAP7_75t_R g2326 ( 
.A(n_2208),
.Y(n_2326)
);

OAI22xp5_ASAP7_75t_L g2327 ( 
.A1(n_2227),
.A2(n_1463),
.B1(n_1464),
.B2(n_1461),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_2116),
.Y(n_2328)
);

INVx1_ASAP7_75t_SL g2329 ( 
.A(n_2115),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2136),
.Y(n_2330)
);

NOR2x1_ASAP7_75t_SL g2331 ( 
.A(n_2154),
.B(n_804),
.Y(n_2331)
);

BUFx2_ASAP7_75t_L g2332 ( 
.A(n_2142),
.Y(n_2332)
);

INVx2_ASAP7_75t_SL g2333 ( 
.A(n_2188),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2193),
.Y(n_2334)
);

NOR2xp33_ASAP7_75t_L g2335 ( 
.A(n_2078),
.B(n_1465),
.Y(n_2335)
);

AO31x2_ASAP7_75t_L g2336 ( 
.A1(n_2095),
.A2(n_2217),
.A3(n_2128),
.B(n_2132),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2141),
.Y(n_2337)
);

AOI21x1_ASAP7_75t_L g2338 ( 
.A1(n_2173),
.A2(n_806),
.B(n_805),
.Y(n_2338)
);

OAI21x1_ASAP7_75t_L g2339 ( 
.A1(n_2230),
.A2(n_811),
.B(n_808),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2200),
.B(n_1468),
.Y(n_2340)
);

OR2x6_ASAP7_75t_L g2341 ( 
.A(n_2188),
.B(n_812),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2221),
.Y(n_2342)
);

AOI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2211),
.A2(n_814),
.B(n_813),
.Y(n_2343)
);

BUFx12f_ASAP7_75t_L g2344 ( 
.A(n_2193),
.Y(n_2344)
);

OA21x2_ASAP7_75t_L g2345 ( 
.A1(n_2231),
.A2(n_1472),
.B(n_1470),
.Y(n_2345)
);

INVx2_ASAP7_75t_SL g2346 ( 
.A(n_2164),
.Y(n_2346)
);

OA21x2_ASAP7_75t_L g2347 ( 
.A1(n_2220),
.A2(n_1475),
.B(n_1474),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2081),
.A2(n_816),
.B(n_815),
.Y(n_2348)
);

AOI22xp33_ASAP7_75t_L g2349 ( 
.A1(n_2224),
.A2(n_1479),
.B1(n_1485),
.B2(n_1476),
.Y(n_2349)
);

A2O1A1Ixp33_ASAP7_75t_L g2350 ( 
.A1(n_2121),
.A2(n_1488),
.B(n_1491),
.C(n_1486),
.Y(n_2350)
);

BUFx2_ASAP7_75t_R g2351 ( 
.A(n_2158),
.Y(n_2351)
);

OAI21x1_ASAP7_75t_L g2352 ( 
.A1(n_2092),
.A2(n_818),
.B(n_817),
.Y(n_2352)
);

AOI22xp33_ASAP7_75t_SL g2353 ( 
.A1(n_2176),
.A2(n_2218),
.B1(n_2162),
.B2(n_2144),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_R g2354 ( 
.A(n_2222),
.B(n_819),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2221),
.Y(n_2355)
);

INVx2_ASAP7_75t_L g2356 ( 
.A(n_2141),
.Y(n_2356)
);

BUFx3_ASAP7_75t_L g2357 ( 
.A(n_2137),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_2183),
.Y(n_2358)
);

OAI21x1_ASAP7_75t_L g2359 ( 
.A1(n_2147),
.A2(n_823),
.B(n_822),
.Y(n_2359)
);

OAI21x1_ASAP7_75t_L g2360 ( 
.A1(n_2159),
.A2(n_827),
.B(n_826),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2183),
.Y(n_2361)
);

OAI21x1_ASAP7_75t_SL g2362 ( 
.A1(n_2165),
.A2(n_831),
.B(n_830),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2210),
.Y(n_2363)
);

BUFx4f_ASAP7_75t_L g2364 ( 
.A(n_2187),
.Y(n_2364)
);

NOR2xp33_ASAP7_75t_SL g2365 ( 
.A(n_2180),
.B(n_1492),
.Y(n_2365)
);

OA21x2_ASAP7_75t_L g2366 ( 
.A1(n_2172),
.A2(n_2213),
.B(n_2169),
.Y(n_2366)
);

HB1xp67_ASAP7_75t_L g2367 ( 
.A(n_2189),
.Y(n_2367)
);

OAI22x1_ASAP7_75t_L g2368 ( 
.A1(n_2179),
.A2(n_1495),
.B1(n_1497),
.B2(n_1494),
.Y(n_2368)
);

OA21x2_ASAP7_75t_L g2369 ( 
.A1(n_2174),
.A2(n_1505),
.B(n_1499),
.Y(n_2369)
);

CKINVDCx11_ASAP7_75t_R g2370 ( 
.A(n_2175),
.Y(n_2370)
);

OAI21x1_ASAP7_75t_L g2371 ( 
.A1(n_2214),
.A2(n_834),
.B(n_833),
.Y(n_2371)
);

AO21x2_ASAP7_75t_L g2372 ( 
.A1(n_2178),
.A2(n_837),
.B(n_835),
.Y(n_2372)
);

AO21x2_ASAP7_75t_L g2373 ( 
.A1(n_2184),
.A2(n_840),
.B(n_839),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_2229),
.Y(n_2374)
);

NAND2x1p5_ASAP7_75t_L g2375 ( 
.A(n_2089),
.B(n_846),
.Y(n_2375)
);

CKINVDCx20_ASAP7_75t_R g2376 ( 
.A(n_2105),
.Y(n_2376)
);

OAI21x1_ASAP7_75t_SL g2377 ( 
.A1(n_2197),
.A2(n_844),
.B(n_842),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2197),
.B(n_845),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2126),
.A2(n_848),
.B(n_847),
.Y(n_2379)
);

AOI221xp5_ASAP7_75t_L g2380 ( 
.A1(n_2166),
.A2(n_1515),
.B1(n_1516),
.B2(n_1514),
.C(n_1513),
.Y(n_2380)
);

AO21x2_ASAP7_75t_L g2381 ( 
.A1(n_2127),
.A2(n_850),
.B(n_849),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_L g2382 ( 
.A1(n_2102),
.A2(n_853),
.B(n_851),
.Y(n_2382)
);

OAI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2143),
.A2(n_1517),
.B(n_857),
.Y(n_2383)
);

OAI21x1_ASAP7_75t_L g2384 ( 
.A1(n_2102),
.A2(n_858),
.B(n_854),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2145),
.Y(n_2385)
);

BUFx12f_ASAP7_75t_L g2386 ( 
.A(n_2083),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2145),
.Y(n_2387)
);

OAI21x1_ASAP7_75t_L g2388 ( 
.A1(n_2102),
.A2(n_861),
.B(n_859),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2145),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2257),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2232),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2255),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2385),
.Y(n_2393)
);

BUFx3_ASAP7_75t_L g2394 ( 
.A(n_2298),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2259),
.Y(n_2395)
);

INVx5_ASAP7_75t_L g2396 ( 
.A(n_2262),
.Y(n_2396)
);

AO21x2_ASAP7_75t_L g2397 ( 
.A1(n_2383),
.A2(n_863),
.B(n_862),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_2279),
.Y(n_2398)
);

OAI21x1_ASAP7_75t_L g2399 ( 
.A1(n_2382),
.A2(n_866),
.B(n_865),
.Y(n_2399)
);

BUFx2_ASAP7_75t_L g2400 ( 
.A(n_2270),
.Y(n_2400)
);

BUFx2_ASAP7_75t_L g2401 ( 
.A(n_2265),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2261),
.Y(n_2402)
);

AOI21xp5_ASAP7_75t_L g2403 ( 
.A1(n_2366),
.A2(n_1007),
.B(n_1006),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2324),
.Y(n_2404)
);

NAND4xp25_ASAP7_75t_SL g2405 ( 
.A(n_2241),
.B(n_13),
.C(n_10),
.D(n_11),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2387),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2263),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2235),
.Y(n_2408)
);

AO21x2_ASAP7_75t_L g2409 ( 
.A1(n_2361),
.A2(n_868),
.B(n_867),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2293),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2389),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2290),
.Y(n_2412)
);

INVx3_ASAP7_75t_L g2413 ( 
.A(n_2291),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2317),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2289),
.Y(n_2415)
);

NAND2xp33_ASAP7_75t_R g2416 ( 
.A(n_2311),
.B(n_1012),
.Y(n_2416)
);

OA21x2_ASAP7_75t_L g2417 ( 
.A1(n_2337),
.A2(n_871),
.B(n_870),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_2314),
.B(n_13),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2268),
.B(n_14),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2292),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2251),
.Y(n_2421)
);

INVx2_ASAP7_75t_L g2422 ( 
.A(n_2276),
.Y(n_2422)
);

BUFx3_ASAP7_75t_L g2423 ( 
.A(n_2324),
.Y(n_2423)
);

OAI21x1_ASAP7_75t_L g2424 ( 
.A1(n_2384),
.A2(n_873),
.B(n_872),
.Y(n_2424)
);

OAI21xp5_ASAP7_75t_L g2425 ( 
.A1(n_2240),
.A2(n_15),
.B(n_16),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2274),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2275),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2283),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2273),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_2386),
.Y(n_2430)
);

OA21x2_ASAP7_75t_L g2431 ( 
.A1(n_2356),
.A2(n_876),
.B(n_874),
.Y(n_2431)
);

AO21x2_ASAP7_75t_L g2432 ( 
.A1(n_2358),
.A2(n_878),
.B(n_877),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2284),
.Y(n_2433)
);

AOI21x1_ASAP7_75t_L g2434 ( 
.A1(n_2256),
.A2(n_882),
.B(n_879),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2234),
.B(n_16),
.Y(n_2435)
);

BUFx6f_ASAP7_75t_L g2436 ( 
.A(n_2288),
.Y(n_2436)
);

INVx4_ASAP7_75t_L g2437 ( 
.A(n_2318),
.Y(n_2437)
);

INVx2_ASAP7_75t_SL g2438 ( 
.A(n_2333),
.Y(n_2438)
);

HB1xp67_ASAP7_75t_L g2439 ( 
.A(n_2329),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2264),
.Y(n_2440)
);

OAI21x1_ASAP7_75t_L g2441 ( 
.A1(n_2388),
.A2(n_884),
.B(n_883),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2285),
.Y(n_2442)
);

NOR2xp33_ASAP7_75t_L g2443 ( 
.A(n_2295),
.B(n_885),
.Y(n_2443)
);

BUFx2_ASAP7_75t_SL g2444 ( 
.A(n_2309),
.Y(n_2444)
);

INVx2_ASAP7_75t_L g2445 ( 
.A(n_2363),
.Y(n_2445)
);

INVx3_ASAP7_75t_L g2446 ( 
.A(n_2246),
.Y(n_2446)
);

OAI21xp5_ASAP7_75t_L g2447 ( 
.A1(n_2250),
.A2(n_17),
.B(n_18),
.Y(n_2447)
);

INVx6_ASAP7_75t_L g2448 ( 
.A(n_2374),
.Y(n_2448)
);

AND2x4_ASAP7_75t_L g2449 ( 
.A(n_2267),
.B(n_2239),
.Y(n_2449)
);

AO21x2_ASAP7_75t_L g2450 ( 
.A1(n_2377),
.A2(n_888),
.B(n_886),
.Y(n_2450)
);

HB1xp67_ASAP7_75t_L g2451 ( 
.A(n_2258),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2277),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2374),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2281),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2342),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2244),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2355),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2260),
.Y(n_2458)
);

HB1xp67_ASAP7_75t_L g2459 ( 
.A(n_2367),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_2272),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2328),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2280),
.Y(n_2462)
);

OAI21x1_ASAP7_75t_L g2463 ( 
.A1(n_2266),
.A2(n_891),
.B(n_889),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2301),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2242),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2321),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2280),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_2247),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_2312),
.Y(n_2469)
);

INVx3_ASAP7_75t_L g2470 ( 
.A(n_2332),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2330),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2237),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2245),
.Y(n_2473)
);

INVx2_ASAP7_75t_SL g2474 ( 
.A(n_2320),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2359),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2357),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2238),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2360),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2271),
.Y(n_2479)
);

AO21x1_ASAP7_75t_SL g2480 ( 
.A1(n_2253),
.A2(n_894),
.B(n_893),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2371),
.Y(n_2481)
);

HB1xp67_ASAP7_75t_L g2482 ( 
.A(n_2346),
.Y(n_2482)
);

NOR2xp67_ASAP7_75t_R g2483 ( 
.A(n_2344),
.B(n_17),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2348),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2352),
.Y(n_2485)
);

AO21x2_ASAP7_75t_L g2486 ( 
.A1(n_2254),
.A2(n_896),
.B(n_895),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2381),
.Y(n_2487)
);

HB1xp67_ASAP7_75t_L g2488 ( 
.A(n_2286),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2282),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2294),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2303),
.Y(n_2491)
);

OAI21x1_ASAP7_75t_L g2492 ( 
.A1(n_2296),
.A2(n_899),
.B(n_898),
.Y(n_2492)
);

OAI21x1_ASAP7_75t_L g2493 ( 
.A1(n_2302),
.A2(n_901),
.B(n_900),
.Y(n_2493)
);

XNOR2xp5_ASAP7_75t_L g2494 ( 
.A(n_2474),
.B(n_2236),
.Y(n_2494)
);

AND2x4_ASAP7_75t_L g2495 ( 
.A(n_2453),
.B(n_2341),
.Y(n_2495)
);

XNOR2xp5_ASAP7_75t_L g2496 ( 
.A(n_2451),
.B(n_2326),
.Y(n_2496)
);

XNOR2xp5_ASAP7_75t_L g2497 ( 
.A(n_2419),
.B(n_2376),
.Y(n_2497)
);

OR2x6_ASAP7_75t_L g2498 ( 
.A(n_2444),
.B(n_2341),
.Y(n_2498)
);

OR2x6_ASAP7_75t_L g2499 ( 
.A(n_2448),
.B(n_2307),
.Y(n_2499)
);

NAND2xp33_ASAP7_75t_R g2500 ( 
.A(n_2446),
.B(n_2354),
.Y(n_2500)
);

AND2x2_ASAP7_75t_L g2501 ( 
.A(n_2435),
.B(n_2299),
.Y(n_2501)
);

NAND2xp33_ASAP7_75t_R g2502 ( 
.A(n_2401),
.B(n_2334),
.Y(n_2502)
);

NOR2xp33_ASAP7_75t_R g2503 ( 
.A(n_2416),
.B(n_2310),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2488),
.B(n_2353),
.Y(n_2504)
);

NAND2xp33_ASAP7_75t_R g2505 ( 
.A(n_2401),
.B(n_2287),
.Y(n_2505)
);

INVxp67_ASAP7_75t_L g2506 ( 
.A(n_2459),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2470),
.B(n_2315),
.Y(n_2507)
);

NAND2xp33_ASAP7_75t_R g2508 ( 
.A(n_2413),
.B(n_2449),
.Y(n_2508)
);

CKINVDCx8_ASAP7_75t_R g2509 ( 
.A(n_2396),
.Y(n_2509)
);

XOR2xp5_ASAP7_75t_L g2510 ( 
.A(n_2430),
.B(n_2351),
.Y(n_2510)
);

INVxp67_ASAP7_75t_L g2511 ( 
.A(n_2439),
.Y(n_2511)
);

AND2x2_ASAP7_75t_L g2512 ( 
.A(n_2445),
.B(n_2369),
.Y(n_2512)
);

AND2x4_ASAP7_75t_L g2513 ( 
.A(n_2423),
.B(n_2243),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2391),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2392),
.B(n_2269),
.Y(n_2515)
);

INVxp67_ASAP7_75t_L g2516 ( 
.A(n_2476),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_R g2517 ( 
.A(n_2394),
.B(n_2370),
.Y(n_2517)
);

CKINVDCx20_ASAP7_75t_R g2518 ( 
.A(n_2448),
.Y(n_2518)
);

NAND2xp33_ASAP7_75t_R g2519 ( 
.A(n_2443),
.B(n_2340),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2460),
.B(n_2252),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2390),
.B(n_2249),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2395),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2418),
.B(n_2421),
.Y(n_2523)
);

BUFx3_ASAP7_75t_L g2524 ( 
.A(n_2404),
.Y(n_2524)
);

NAND2xp5_ASAP7_75t_L g2525 ( 
.A(n_2402),
.B(n_2407),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2410),
.B(n_2335),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_R g2527 ( 
.A(n_2404),
.B(n_2365),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2398),
.B(n_2319),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_2429),
.Y(n_2529)
);

XOR2x2_ASAP7_75t_SL g2530 ( 
.A(n_2405),
.B(n_2325),
.Y(n_2530)
);

INVx5_ASAP7_75t_L g2531 ( 
.A(n_2436),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_R g2532 ( 
.A(n_2396),
.B(n_2364),
.Y(n_2532)
);

XNOR2xp5_ASAP7_75t_L g2533 ( 
.A(n_2482),
.B(n_2368),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2420),
.B(n_2323),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2491),
.B(n_2252),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2393),
.Y(n_2536)
);

NAND2xp33_ASAP7_75t_R g2537 ( 
.A(n_2400),
.B(n_2305),
.Y(n_2537)
);

AND2x4_ASAP7_75t_L g2538 ( 
.A(n_2437),
.B(n_2372),
.Y(n_2538)
);

NOR2xp33_ASAP7_75t_R g2539 ( 
.A(n_2436),
.B(n_2338),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2440),
.Y(n_2540)
);

NOR2xp33_ASAP7_75t_R g2541 ( 
.A(n_2430),
.B(n_2322),
.Y(n_2541)
);

AND2x4_ASAP7_75t_L g2542 ( 
.A(n_2438),
.B(n_2233),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2408),
.B(n_2412),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_2422),
.B(n_2378),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_2442),
.B(n_2248),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2406),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_R g2547 ( 
.A(n_2452),
.B(n_2454),
.Y(n_2547)
);

XNOR2xp5_ASAP7_75t_L g2548 ( 
.A(n_2426),
.B(n_2327),
.Y(n_2548)
);

XOR2xp5_ASAP7_75t_L g2549 ( 
.A(n_2425),
.B(n_2375),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2411),
.B(n_2380),
.Y(n_2550)
);

AND2x2_ASAP7_75t_SL g2551 ( 
.A(n_2400),
.B(n_2347),
.Y(n_2551)
);

OR2x6_ASAP7_75t_L g2552 ( 
.A(n_2447),
.B(n_2297),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2414),
.B(n_2349),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2514),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2520),
.B(n_2455),
.Y(n_2555)
);

OR2x2_ASAP7_75t_L g2556 ( 
.A(n_2504),
.B(n_2546),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2535),
.B(n_2457),
.Y(n_2557)
);

OR2x2_ASAP7_75t_L g2558 ( 
.A(n_2536),
.B(n_2461),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2523),
.B(n_2415),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2501),
.B(n_2427),
.Y(n_2560)
);

BUFx2_ASAP7_75t_L g2561 ( 
.A(n_2547),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2545),
.B(n_2428),
.Y(n_2562)
);

INVxp67_ASAP7_75t_SL g2563 ( 
.A(n_2506),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_SL g2564 ( 
.A(n_2530),
.B(n_2479),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2512),
.B(n_2433),
.Y(n_2565)
);

AND2x2_ASAP7_75t_L g2566 ( 
.A(n_2516),
.B(n_2469),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2511),
.B(n_2466),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2513),
.B(n_2469),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2522),
.Y(n_2569)
);

HB1xp67_ASAP7_75t_L g2570 ( 
.A(n_2537),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2525),
.Y(n_2571)
);

AND2x2_ASAP7_75t_L g2572 ( 
.A(n_2544),
.B(n_2487),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2543),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2542),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2515),
.B(n_2462),
.Y(n_2575)
);

INVxp67_ASAP7_75t_SL g2576 ( 
.A(n_2521),
.Y(n_2576)
);

INVx1_ASAP7_75t_SL g2577 ( 
.A(n_2496),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2528),
.B(n_2471),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2495),
.B(n_2467),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2526),
.B(n_2464),
.Y(n_2580)
);

AND2x2_ASAP7_75t_L g2581 ( 
.A(n_2529),
.B(n_2480),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2534),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2551),
.B(n_2480),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2550),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2553),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2538),
.Y(n_2586)
);

BUFx3_ASAP7_75t_L g2587 ( 
.A(n_2518),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2507),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2548),
.Y(n_2589)
);

AND2x2_ASAP7_75t_L g2590 ( 
.A(n_2533),
.B(n_2450),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2549),
.B(n_2552),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2552),
.B(n_2483),
.Y(n_2592)
);

OAI221xp5_ASAP7_75t_SL g2593 ( 
.A1(n_2498),
.A2(n_2304),
.B1(n_2350),
.B2(n_2313),
.C(n_2379),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_SL g2594 ( 
.A(n_2503),
.B(n_2541),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2524),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2540),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2498),
.B(n_2458),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2497),
.B(n_2397),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2499),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2499),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2531),
.B(n_2456),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2494),
.B(n_2484),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2531),
.B(n_2473),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2539),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2509),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2505),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2519),
.A2(n_2500),
.B1(n_2502),
.B2(n_2508),
.Y(n_2607)
);

INVx4_ASAP7_75t_L g2608 ( 
.A(n_2532),
.Y(n_2608)
);

INVx5_ASAP7_75t_L g2609 ( 
.A(n_2527),
.Y(n_2609)
);

OR2x2_ASAP7_75t_L g2610 ( 
.A(n_2510),
.B(n_2472),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2517),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2506),
.B(n_2485),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_2546),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2523),
.B(n_2409),
.Y(n_2614)
);

INVx4_ASAP7_75t_L g2615 ( 
.A(n_2609),
.Y(n_2615)
);

INVx5_ASAP7_75t_L g2616 ( 
.A(n_2609),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2554),
.Y(n_2617)
);

INVx2_ASAP7_75t_SL g2618 ( 
.A(n_2595),
.Y(n_2618)
);

INVx2_ASAP7_75t_SL g2619 ( 
.A(n_2596),
.Y(n_2619)
);

INVx1_ASAP7_75t_SL g2620 ( 
.A(n_2561),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2566),
.Y(n_2621)
);

AND2x2_ASAP7_75t_L g2622 ( 
.A(n_2570),
.B(n_2477),
.Y(n_2622)
);

AO21x2_ASAP7_75t_L g2623 ( 
.A1(n_2592),
.A2(n_2468),
.B(n_2403),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2613),
.Y(n_2624)
);

OAI221xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2607),
.A2(n_2343),
.B1(n_2481),
.B2(n_2478),
.C(n_2475),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2602),
.B(n_2465),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2606),
.B(n_2561),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2568),
.B(n_2486),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2558),
.Y(n_2629)
);

AND2x2_ASAP7_75t_L g2630 ( 
.A(n_2588),
.B(n_2432),
.Y(n_2630)
);

AND2x2_ASAP7_75t_L g2631 ( 
.A(n_2563),
.B(n_2373),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2612),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2560),
.B(n_2278),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_2576),
.B(n_2489),
.Y(n_2634)
);

AOI22xp33_ASAP7_75t_L g2635 ( 
.A1(n_2590),
.A2(n_2362),
.B1(n_2300),
.B2(n_2308),
.Y(n_2635)
);

NOR2xp33_ASAP7_75t_R g2636 ( 
.A(n_2609),
.B(n_18),
.Y(n_2636)
);

INVx2_ASAP7_75t_SL g2637 ( 
.A(n_2587),
.Y(n_2637)
);

CKINVDCx20_ASAP7_75t_R g2638 ( 
.A(n_2577),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2569),
.Y(n_2639)
);

INVx2_ASAP7_75t_SL g2640 ( 
.A(n_2559),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2582),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2575),
.B(n_2490),
.Y(n_2642)
);

OR2x2_ASAP7_75t_L g2643 ( 
.A(n_2556),
.B(n_2336),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2565),
.Y(n_2644)
);

AO21x2_ASAP7_75t_L g2645 ( 
.A1(n_2601),
.A2(n_2434),
.B(n_2424),
.Y(n_2645)
);

AND2x2_ASAP7_75t_L g2646 ( 
.A(n_2610),
.B(n_2417),
.Y(n_2646)
);

INVxp67_ASAP7_75t_SL g2647 ( 
.A(n_2578),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2555),
.Y(n_2648)
);

INVxp67_ASAP7_75t_SL g2649 ( 
.A(n_2603),
.Y(n_2649)
);

OR2x2_ASAP7_75t_L g2650 ( 
.A(n_2585),
.B(n_2336),
.Y(n_2650)
);

AND2x2_ASAP7_75t_L g2651 ( 
.A(n_2579),
.B(n_2431),
.Y(n_2651)
);

NOR2xp67_ASAP7_75t_SL g2652 ( 
.A(n_2608),
.B(n_2345),
.Y(n_2652)
);

NAND2xp5_ASAP7_75t_L g2653 ( 
.A(n_2584),
.B(n_19),
.Y(n_2653)
);

AO21x2_ASAP7_75t_L g2654 ( 
.A1(n_2591),
.A2(n_2441),
.B(n_2399),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2555),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2557),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2571),
.Y(n_2657)
);

OAI221xp5_ASAP7_75t_L g2658 ( 
.A1(n_2593),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.C(n_22),
.Y(n_2658)
);

BUFx3_ASAP7_75t_L g2659 ( 
.A(n_2611),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2562),
.B(n_2463),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2557),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2573),
.Y(n_2662)
);

HB1xp67_ASAP7_75t_L g2663 ( 
.A(n_2580),
.Y(n_2663)
);

OAI22xp5_ASAP7_75t_L g2664 ( 
.A1(n_2594),
.A2(n_2331),
.B1(n_2316),
.B2(n_2492),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2586),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2574),
.Y(n_2666)
);

INVx1_ASAP7_75t_SL g2667 ( 
.A(n_2605),
.Y(n_2667)
);

BUFx6f_ASAP7_75t_L g2668 ( 
.A(n_2567),
.Y(n_2668)
);

AO21x2_ASAP7_75t_L g2669 ( 
.A1(n_2604),
.A2(n_2493),
.B(n_2306),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2597),
.B(n_2572),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2614),
.B(n_2339),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2599),
.Y(n_2672)
);

NOR2xp67_ASAP7_75t_SL g2673 ( 
.A(n_2564),
.B(n_902),
.Y(n_2673)
);

BUFx3_ASAP7_75t_L g2674 ( 
.A(n_2581),
.Y(n_2674)
);

INVxp67_ASAP7_75t_SL g2675 ( 
.A(n_2600),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2583),
.Y(n_2676)
);

INVx3_ASAP7_75t_L g2677 ( 
.A(n_2589),
.Y(n_2677)
);

INVxp67_ASAP7_75t_L g2678 ( 
.A(n_2598),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2570),
.B(n_20),
.Y(n_2679)
);

AOI33xp33_ASAP7_75t_L g2680 ( 
.A1(n_2584),
.A2(n_24),
.A3(n_26),
.B1(n_22),
.B2(n_23),
.B3(n_25),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2554),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2613),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2613),
.Y(n_2683)
);

HB1xp67_ASAP7_75t_L g2684 ( 
.A(n_2566),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2613),
.Y(n_2685)
);

BUFx2_ASAP7_75t_L g2686 ( 
.A(n_2561),
.Y(n_2686)
);

AOI221xp5_ASAP7_75t_L g2687 ( 
.A1(n_2584),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.C(n_26),
.Y(n_2687)
);

HB1xp67_ASAP7_75t_L g2688 ( 
.A(n_2566),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2613),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2570),
.B(n_27),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2576),
.B(n_27),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2570),
.B(n_28),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2554),
.Y(n_2693)
);

NAND3xp33_ASAP7_75t_SL g2694 ( 
.A(n_2607),
.B(n_28),
.C(n_29),
.Y(n_2694)
);

INVxp67_ASAP7_75t_SL g2695 ( 
.A(n_2576),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2554),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2663),
.B(n_29),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2641),
.Y(n_2698)
);

NAND2x1_ASAP7_75t_L g2699 ( 
.A(n_2686),
.B(n_30),
.Y(n_2699)
);

NOR2x1_ASAP7_75t_SL g2700 ( 
.A(n_2616),
.B(n_2615),
.Y(n_2700)
);

OR2x2_ASAP7_75t_L g2701 ( 
.A(n_2621),
.B(n_30),
.Y(n_2701)
);

NAND2x1p5_ASAP7_75t_L g2702 ( 
.A(n_2616),
.B(n_904),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2617),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2684),
.B(n_31),
.Y(n_2704)
);

AND2x4_ASAP7_75t_L g2705 ( 
.A(n_2656),
.B(n_32),
.Y(n_2705)
);

AND2x2_ASAP7_75t_L g2706 ( 
.A(n_2688),
.B(n_33),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2658),
.A2(n_2694),
.B1(n_2678),
.B2(n_2687),
.Y(n_2707)
);

NOR2xp33_ASAP7_75t_SL g2708 ( 
.A(n_2616),
.B(n_33),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2665),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2647),
.B(n_34),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2676),
.B(n_34),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2674),
.B(n_35),
.Y(n_2712)
);

AND2x4_ASAP7_75t_L g2713 ( 
.A(n_2661),
.B(n_35),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2649),
.B(n_36),
.Y(n_2714)
);

AND2x2_ASAP7_75t_L g2715 ( 
.A(n_2670),
.B(n_2648),
.Y(n_2715)
);

OAI21xp5_ASAP7_75t_L g2716 ( 
.A1(n_2691),
.A2(n_36),
.B(n_37),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2655),
.B(n_37),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2629),
.B(n_2632),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2695),
.B(n_38),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2665),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2627),
.B(n_38),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2620),
.B(n_39),
.Y(n_2722)
);

AND2x2_ASAP7_75t_L g2723 ( 
.A(n_2666),
.B(n_39),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2681),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2666),
.B(n_40),
.Y(n_2725)
);

OR2x2_ASAP7_75t_L g2726 ( 
.A(n_2643),
.B(n_41),
.Y(n_2726)
);

AND2x2_ASAP7_75t_L g2727 ( 
.A(n_2640),
.B(n_41),
.Y(n_2727)
);

OR2x2_ASAP7_75t_L g2728 ( 
.A(n_2644),
.B(n_2672),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2675),
.B(n_42),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2668),
.B(n_42),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2693),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2696),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2639),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2668),
.B(n_43),
.Y(n_2734)
);

HB1xp67_ASAP7_75t_L g2735 ( 
.A(n_2622),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2624),
.Y(n_2736)
);

AND2x2_ASAP7_75t_L g2737 ( 
.A(n_2626),
.B(n_43),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2619),
.B(n_44),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2628),
.B(n_44),
.Y(n_2739)
);

INVxp67_ASAP7_75t_L g2740 ( 
.A(n_2618),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2657),
.B(n_45),
.Y(n_2741)
);

OR2x2_ASAP7_75t_L g2742 ( 
.A(n_2662),
.B(n_45),
.Y(n_2742)
);

OR2x2_ASAP7_75t_L g2743 ( 
.A(n_2634),
.B(n_46),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2682),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2683),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_2685),
.B(n_47),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2689),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_SL g2748 ( 
.A(n_2636),
.B(n_47),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2650),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2642),
.Y(n_2750)
);

O2A1O1Ixp33_ASAP7_75t_L g2751 ( 
.A1(n_2625),
.A2(n_50),
.B(n_48),
.C(n_49),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2631),
.Y(n_2752)
);

BUFx2_ASAP7_75t_L g2753 ( 
.A(n_2623),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2633),
.B(n_49),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2630),
.Y(n_2755)
);

AND2x4_ASAP7_75t_L g2756 ( 
.A(n_2660),
.B(n_51),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2651),
.Y(n_2757)
);

INVxp67_ASAP7_75t_SL g2758 ( 
.A(n_2646),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2671),
.B(n_51),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2653),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2667),
.B(n_2677),
.Y(n_2761)
);

OR2x2_ASAP7_75t_L g2762 ( 
.A(n_2679),
.B(n_52),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2659),
.B(n_2637),
.Y(n_2763)
);

OR2x2_ASAP7_75t_L g2764 ( 
.A(n_2690),
.B(n_52),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2645),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2692),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2654),
.Y(n_2767)
);

INVx4_ASAP7_75t_L g2768 ( 
.A(n_2669),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2680),
.B(n_53),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2638),
.B(n_53),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2664),
.Y(n_2771)
);

INVxp67_ASAP7_75t_L g2772 ( 
.A(n_2673),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2635),
.B(n_55),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2652),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2647),
.B(n_55),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2617),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_2641),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2621),
.B(n_56),
.Y(n_2778)
);

AND2x2_ASAP7_75t_L g2779 ( 
.A(n_2663),
.B(n_56),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2617),
.Y(n_2780)
);

HB1xp67_ASAP7_75t_L g2781 ( 
.A(n_2663),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2641),
.Y(n_2782)
);

AND2x2_ASAP7_75t_L g2783 ( 
.A(n_2663),
.B(n_57),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2617),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2617),
.Y(n_2785)
);

INVxp67_ASAP7_75t_L g2786 ( 
.A(n_2649),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2641),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2621),
.B(n_58),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2617),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_2621),
.B(n_58),
.Y(n_2790)
);

NAND2xp5_ASAP7_75t_L g2791 ( 
.A(n_2647),
.B(n_59),
.Y(n_2791)
);

NOR2x1p5_ASAP7_75t_L g2792 ( 
.A(n_2615),
.B(n_59),
.Y(n_2792)
);

NAND4xp25_ASAP7_75t_L g2793 ( 
.A(n_2658),
.B(n_63),
.C(n_60),
.D(n_61),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2617),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2641),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2617),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2641),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2663),
.B(n_61),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2663),
.B(n_64),
.Y(n_2799)
);

NAND2x1_ASAP7_75t_L g2800 ( 
.A(n_2686),
.B(n_64),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2647),
.B(n_66),
.Y(n_2801)
);

OR2x2_ASAP7_75t_L g2802 ( 
.A(n_2621),
.B(n_68),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2617),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2617),
.Y(n_2804)
);

AND2x2_ASAP7_75t_SL g2805 ( 
.A(n_2615),
.B(n_69),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2621),
.B(n_69),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2617),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2663),
.B(n_70),
.Y(n_2808)
);

INVxp67_ASAP7_75t_L g2809 ( 
.A(n_2649),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2647),
.B(n_70),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2617),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2641),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2641),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2663),
.B(n_71),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2786),
.B(n_71),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2809),
.B(n_72),
.Y(n_2816)
);

AO221x2_ASAP7_75t_L g2817 ( 
.A1(n_2716),
.A2(n_74),
.B1(n_76),
.B2(n_73),
.C(n_75),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2760),
.B(n_72),
.Y(n_2818)
);

OR2x2_ASAP7_75t_L g2819 ( 
.A(n_2781),
.B(n_73),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2758),
.B(n_74),
.Y(n_2820)
);

NOR2xp33_ASAP7_75t_R g2821 ( 
.A(n_2708),
.B(n_75),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2709),
.Y(n_2822)
);

NAND2xp33_ASAP7_75t_R g2823 ( 
.A(n_2756),
.B(n_77),
.Y(n_2823)
);

AO221x2_ASAP7_75t_L g2824 ( 
.A1(n_2769),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.C(n_81),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2752),
.B(n_2726),
.Y(n_2825)
);

OAI22xp33_ASAP7_75t_L g2826 ( 
.A1(n_2793),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_2826)
);

CKINVDCx5p33_ASAP7_75t_R g2827 ( 
.A(n_2805),
.Y(n_2827)
);

NAND2xp33_ASAP7_75t_L g2828 ( 
.A(n_2792),
.B(n_83),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2771),
.B(n_85),
.Y(n_2829)
);

AO221x2_ASAP7_75t_L g2830 ( 
.A1(n_2766),
.A2(n_2714),
.B1(n_2719),
.B2(n_2775),
.C(n_2710),
.Y(n_2830)
);

AO221x2_ASAP7_75t_L g2831 ( 
.A1(n_2791),
.A2(n_87),
.B1(n_89),
.B2(n_86),
.C(n_88),
.Y(n_2831)
);

CKINVDCx5p33_ASAP7_75t_R g2832 ( 
.A(n_2770),
.Y(n_2832)
);

AO221x2_ASAP7_75t_L g2833 ( 
.A1(n_2801),
.A2(n_87),
.B1(n_90),
.B2(n_86),
.C(n_89),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2749),
.B(n_85),
.Y(n_2834)
);

AO221x2_ASAP7_75t_L g2835 ( 
.A1(n_2810),
.A2(n_92),
.B1(n_90),
.B2(n_91),
.C(n_93),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2761),
.B(n_2735),
.Y(n_2836)
);

NAND2xp33_ASAP7_75t_SL g2837 ( 
.A(n_2699),
.B(n_94),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_L g2838 ( 
.A(n_2718),
.B(n_95),
.Y(n_2838)
);

AO221x2_ASAP7_75t_L g2839 ( 
.A1(n_2754),
.A2(n_97),
.B1(n_101),
.B2(n_96),
.C(n_100),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_2750),
.B(n_95),
.Y(n_2840)
);

AND2x4_ASAP7_75t_SL g2841 ( 
.A(n_2763),
.B(n_96),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2743),
.B(n_97),
.Y(n_2842)
);

AO221x2_ASAP7_75t_L g2843 ( 
.A1(n_2734),
.A2(n_103),
.B1(n_105),
.B2(n_102),
.C(n_104),
.Y(n_2843)
);

AOI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2707),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_2844)
);

OAI221xp5_ASAP7_75t_L g2845 ( 
.A1(n_2773),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.C(n_109),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2733),
.B(n_106),
.Y(n_2846)
);

NOR2xp33_ASAP7_75t_SL g2847 ( 
.A(n_2772),
.B(n_107),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2703),
.B(n_109),
.Y(n_2848)
);

NOR2x1_ASAP7_75t_L g2849 ( 
.A(n_2753),
.B(n_110),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2774),
.B(n_110),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2724),
.B(n_111),
.Y(n_2851)
);

OAI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2800),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2731),
.B(n_113),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2732),
.B(n_114),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2720),
.Y(n_2855)
);

NAND2xp33_ASAP7_75t_SL g2856 ( 
.A(n_2748),
.B(n_114),
.Y(n_2856)
);

AO221x2_ASAP7_75t_L g2857 ( 
.A1(n_2759),
.A2(n_117),
.B1(n_119),
.B2(n_116),
.C(n_118),
.Y(n_2857)
);

AOI22xp5_ASAP7_75t_L g2858 ( 
.A1(n_2756),
.A2(n_2739),
.B1(n_2740),
.B2(n_2730),
.Y(n_2858)
);

OAI221xp5_ASAP7_75t_L g2859 ( 
.A1(n_2751),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.C(n_120),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2757),
.A2(n_121),
.B1(n_115),
.B2(n_120),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2776),
.B(n_122),
.Y(n_2861)
);

OAI22xp33_ASAP7_75t_L g2862 ( 
.A1(n_2701),
.A2(n_124),
.B1(n_122),
.B2(n_123),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2780),
.B(n_123),
.Y(n_2863)
);

OAI221xp5_ASAP7_75t_L g2864 ( 
.A1(n_2741),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.C(n_127),
.Y(n_2864)
);

CKINVDCx5p33_ASAP7_75t_R g2865 ( 
.A(n_2722),
.Y(n_2865)
);

NAND2xp33_ASAP7_75t_SL g2866 ( 
.A(n_2729),
.B(n_126),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2762),
.B(n_127),
.Y(n_2867)
);

HB1xp67_ASAP7_75t_L g2868 ( 
.A(n_2736),
.Y(n_2868)
);

NOR2xp33_ASAP7_75t_L g2869 ( 
.A(n_2764),
.B(n_2742),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2784),
.B(n_128),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2785),
.B(n_128),
.Y(n_2871)
);

AOI22xp5_ASAP7_75t_L g2872 ( 
.A1(n_2721),
.A2(n_2705),
.B1(n_2713),
.B2(n_2737),
.Y(n_2872)
);

AO221x2_ASAP7_75t_L g2873 ( 
.A1(n_2755),
.A2(n_131),
.B1(n_133),
.B2(n_130),
.C(n_132),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2715),
.B(n_2700),
.Y(n_2874)
);

AOI22xp5_ASAP7_75t_L g2875 ( 
.A1(n_2697),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2789),
.B(n_129),
.Y(n_2876)
);

AO221x2_ASAP7_75t_L g2877 ( 
.A1(n_2746),
.A2(n_134),
.B1(n_136),
.B2(n_133),
.C(n_135),
.Y(n_2877)
);

INVxp67_ASAP7_75t_L g2878 ( 
.A(n_2728),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2794),
.B(n_132),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2796),
.Y(n_2880)
);

AND2x2_ASAP7_75t_L g2881 ( 
.A(n_2745),
.B(n_134),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2803),
.B(n_135),
.Y(n_2882)
);

AOI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2779),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2804),
.B(n_2807),
.Y(n_2884)
);

OAI221xp5_ASAP7_75t_L g2885 ( 
.A1(n_2767),
.A2(n_143),
.B1(n_140),
.B2(n_141),
.C(n_144),
.Y(n_2885)
);

NAND2xp33_ASAP7_75t_SL g2886 ( 
.A(n_2723),
.B(n_140),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2811),
.B(n_141),
.Y(n_2887)
);

INVxp67_ASAP7_75t_L g2888 ( 
.A(n_2725),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2698),
.B(n_2777),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2782),
.B(n_143),
.Y(n_2890)
);

OAI22xp33_ASAP7_75t_L g2891 ( 
.A1(n_2778),
.A2(n_146),
.B1(n_144),
.B2(n_145),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2787),
.B(n_145),
.Y(n_2892)
);

NAND2xp5_ASAP7_75t_L g2893 ( 
.A(n_2795),
.B(n_146),
.Y(n_2893)
);

NAND2xp33_ASAP7_75t_SL g2894 ( 
.A(n_2712),
.B(n_147),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2797),
.B(n_2812),
.Y(n_2895)
);

OR2x2_ASAP7_75t_L g2896 ( 
.A(n_2747),
.B(n_148),
.Y(n_2896)
);

OAI221xp5_ASAP7_75t_L g2897 ( 
.A1(n_2702),
.A2(n_2788),
.B1(n_2806),
.B2(n_2802),
.C(n_2790),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2813),
.B(n_148),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2744),
.B(n_149),
.Y(n_2899)
);

NAND2xp33_ASAP7_75t_R g2900 ( 
.A(n_2783),
.B(n_149),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2753),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_2798),
.A2(n_153),
.B1(n_150),
.B2(n_152),
.Y(n_2902)
);

NAND2xp33_ASAP7_75t_R g2903 ( 
.A(n_2799),
.B(n_150),
.Y(n_2903)
);

BUFx2_ASAP7_75t_L g2904 ( 
.A(n_2808),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2765),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2814),
.B(n_152),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2704),
.B(n_153),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2706),
.B(n_154),
.Y(n_2908)
);

INVx2_ASAP7_75t_SL g2909 ( 
.A(n_2738),
.Y(n_2909)
);

INVxp67_ASAP7_75t_L g2910 ( 
.A(n_2717),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_SL g2911 ( 
.A(n_2768),
.B(n_2727),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2711),
.B(n_154),
.Y(n_2912)
);

NOR2x1_ASAP7_75t_L g2913 ( 
.A(n_2753),
.B(n_155),
.Y(n_2913)
);

NAND2xp5_ASAP7_75t_L g2914 ( 
.A(n_2786),
.B(n_155),
.Y(n_2914)
);

AO221x2_ASAP7_75t_L g2915 ( 
.A1(n_2716),
.A2(n_159),
.B1(n_161),
.B2(n_158),
.C(n_160),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2760),
.B(n_157),
.Y(n_2916)
);

AO221x2_ASAP7_75t_L g2917 ( 
.A1(n_2716),
.A2(n_163),
.B1(n_165),
.B2(n_162),
.C(n_164),
.Y(n_2917)
);

AO221x2_ASAP7_75t_L g2918 ( 
.A1(n_2716),
.A2(n_165),
.B1(n_168),
.B2(n_163),
.C(n_167),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2786),
.B(n_161),
.Y(n_2919)
);

NOR4xp25_ASAP7_75t_SL g2920 ( 
.A(n_2753),
.B(n_169),
.C(n_167),
.D(n_168),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2786),
.B(n_169),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2786),
.B(n_170),
.Y(n_2922)
);

AO221x2_ASAP7_75t_L g2923 ( 
.A1(n_2716),
.A2(n_173),
.B1(n_175),
.B2(n_172),
.C(n_174),
.Y(n_2923)
);

AO221x2_ASAP7_75t_L g2924 ( 
.A1(n_2716),
.A2(n_175),
.B1(n_179),
.B2(n_173),
.C(n_178),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2786),
.B(n_171),
.Y(n_2925)
);

NOR4xp25_ASAP7_75t_SL g2926 ( 
.A(n_2753),
.B(n_181),
.C(n_178),
.D(n_180),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2786),
.B(n_181),
.Y(n_2927)
);

AOI22xp5_ASAP7_75t_L g2928 ( 
.A1(n_2793),
.A2(n_184),
.B1(n_182),
.B2(n_183),
.Y(n_2928)
);

OAI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2707),
.A2(n_186),
.B1(n_182),
.B2(n_185),
.Y(n_2929)
);

AOI22xp5_ASAP7_75t_L g2930 ( 
.A1(n_2793),
.A2(n_189),
.B1(n_185),
.B2(n_188),
.Y(n_2930)
);

AO221x2_ASAP7_75t_L g2931 ( 
.A1(n_2716),
.A2(n_191),
.B1(n_193),
.B2(n_190),
.C(n_192),
.Y(n_2931)
);

AO221x2_ASAP7_75t_L g2932 ( 
.A1(n_2716),
.A2(n_192),
.B1(n_195),
.B2(n_190),
.C(n_194),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2786),
.B(n_189),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2786),
.B(n_194),
.Y(n_2934)
);

NOR2xp33_ASAP7_75t_SL g2935 ( 
.A(n_2805),
.B(n_197),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2781),
.Y(n_2936)
);

NOR2x1_ASAP7_75t_L g2937 ( 
.A(n_2753),
.B(n_198),
.Y(n_2937)
);

OR2x2_ASAP7_75t_L g2938 ( 
.A(n_2781),
.B(n_198),
.Y(n_2938)
);

AO221x2_ASAP7_75t_L g2939 ( 
.A1(n_2716),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.C(n_202),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2786),
.B(n_199),
.Y(n_2940)
);

AO221x2_ASAP7_75t_L g2941 ( 
.A1(n_2716),
.A2(n_204),
.B1(n_206),
.B2(n_203),
.C(n_205),
.Y(n_2941)
);

AOI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2793),
.A2(n_204),
.B1(n_200),
.B2(n_203),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2786),
.B(n_206),
.Y(n_2943)
);

AOI22xp5_ASAP7_75t_L g2944 ( 
.A1(n_2793),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2944)
);

OAI221xp5_ASAP7_75t_L g2945 ( 
.A1(n_2707),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.C(n_212),
.Y(n_2945)
);

OAI22xp33_ASAP7_75t_L g2946 ( 
.A1(n_2793),
.A2(n_214),
.B1(n_211),
.B2(n_213),
.Y(n_2946)
);

NOR2x1_ASAP7_75t_L g2947 ( 
.A(n_2753),
.B(n_213),
.Y(n_2947)
);

NOR2x1_ASAP7_75t_L g2948 ( 
.A(n_2753),
.B(n_215),
.Y(n_2948)
);

NAND2xp33_ASAP7_75t_SL g2949 ( 
.A(n_2699),
.B(n_215),
.Y(n_2949)
);

NAND2xp33_ASAP7_75t_SL g2950 ( 
.A(n_2699),
.B(n_216),
.Y(n_2950)
);

AOI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2793),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_2951)
);

AND2x4_ASAP7_75t_L g2952 ( 
.A(n_2761),
.B(n_217),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2786),
.B(n_218),
.Y(n_2953)
);

NOR2x1_ASAP7_75t_L g2954 ( 
.A(n_2753),
.B(n_219),
.Y(n_2954)
);

AND2x2_ASAP7_75t_L g2955 ( 
.A(n_2758),
.B(n_220),
.Y(n_2955)
);

INVx2_ASAP7_75t_L g2956 ( 
.A(n_2709),
.Y(n_2956)
);

AO221x2_ASAP7_75t_L g2957 ( 
.A1(n_2716),
.A2(n_224),
.B1(n_226),
.B2(n_222),
.C(n_225),
.Y(n_2957)
);

OAI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_2793),
.A2(n_224),
.B1(n_221),
.B2(n_222),
.Y(n_2958)
);

AO221x2_ASAP7_75t_L g2959 ( 
.A1(n_2716),
.A2(n_227),
.B1(n_229),
.B2(n_225),
.C(n_228),
.Y(n_2959)
);

AOI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2793),
.A2(n_228),
.B1(n_221),
.B2(n_227),
.Y(n_2960)
);

AO221x2_ASAP7_75t_L g2961 ( 
.A1(n_2716),
.A2(n_231),
.B1(n_233),
.B2(n_230),
.C(n_232),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2763),
.Y(n_2962)
);

INVx1_ASAP7_75t_SL g2963 ( 
.A(n_2841),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2880),
.Y(n_2964)
);

INVx1_ASAP7_75t_SL g2965 ( 
.A(n_2827),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2830),
.B(n_229),
.Y(n_2966)
);

INVx1_ASAP7_75t_L g2967 ( 
.A(n_2884),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2868),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2878),
.B(n_230),
.Y(n_2969)
);

OR2x2_ASAP7_75t_L g2970 ( 
.A(n_2825),
.B(n_231),
.Y(n_2970)
);

INVx2_ASAP7_75t_L g2971 ( 
.A(n_2936),
.Y(n_2971)
);

CKINVDCx16_ASAP7_75t_R g2972 ( 
.A(n_2900),
.Y(n_2972)
);

NAND3xp33_ASAP7_75t_L g2973 ( 
.A(n_2928),
.B(n_232),
.C(n_233),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2836),
.Y(n_2974)
);

NOR2x1p5_ASAP7_75t_L g2975 ( 
.A(n_2832),
.B(n_234),
.Y(n_2975)
);

INVxp67_ASAP7_75t_SL g2976 ( 
.A(n_2849),
.Y(n_2976)
);

HB1xp67_ASAP7_75t_L g2977 ( 
.A(n_2913),
.Y(n_2977)
);

OAI21x1_ASAP7_75t_L g2978 ( 
.A1(n_2901),
.A2(n_234),
.B(n_235),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2874),
.B(n_236),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2962),
.B(n_236),
.Y(n_2980)
);

OR2x2_ASAP7_75t_L g2981 ( 
.A(n_2904),
.B(n_2888),
.Y(n_2981)
);

AOI22x1_ASAP7_75t_L g2982 ( 
.A1(n_2955),
.A2(n_239),
.B1(n_237),
.B2(n_238),
.Y(n_2982)
);

AND2x4_ASAP7_75t_L g2983 ( 
.A(n_2909),
.B(n_238),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2905),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2822),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2889),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2895),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2890),
.Y(n_2988)
);

INVx1_ASAP7_75t_SL g2989 ( 
.A(n_2821),
.Y(n_2989)
);

OR2x2_ASAP7_75t_L g2990 ( 
.A(n_2834),
.B(n_237),
.Y(n_2990)
);

NAND2xp33_ASAP7_75t_SL g2991 ( 
.A(n_2823),
.B(n_2903),
.Y(n_2991)
);

AND2x2_ASAP7_75t_L g2992 ( 
.A(n_2911),
.B(n_239),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_2865),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2869),
.B(n_240),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2892),
.Y(n_2995)
);

INVx2_ASAP7_75t_L g2996 ( 
.A(n_2855),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_2866),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2820),
.B(n_240),
.Y(n_2998)
);

AND2x4_ASAP7_75t_L g2999 ( 
.A(n_2910),
.B(n_241),
.Y(n_2999)
);

AND2x2_ASAP7_75t_L g3000 ( 
.A(n_2956),
.B(n_241),
.Y(n_3000)
);

INVx2_ASAP7_75t_L g3001 ( 
.A(n_2896),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2858),
.B(n_242),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2952),
.Y(n_3003)
);

BUFx2_ASAP7_75t_L g3004 ( 
.A(n_2937),
.Y(n_3004)
);

AND2x2_ASAP7_75t_L g3005 ( 
.A(n_2881),
.B(n_242),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2947),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2899),
.B(n_243),
.Y(n_3007)
);

INVx1_ASAP7_75t_SL g3008 ( 
.A(n_2894),
.Y(n_3008)
);

OR2x2_ASAP7_75t_L g3009 ( 
.A(n_2819),
.B(n_243),
.Y(n_3009)
);

AND2x2_ASAP7_75t_L g3010 ( 
.A(n_2872),
.B(n_244),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2948),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_2938),
.B(n_244),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2838),
.B(n_245),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2954),
.Y(n_3014)
);

OAI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2935),
.A2(n_245),
.B(n_246),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2846),
.B(n_246),
.Y(n_3016)
);

INVx1_ASAP7_75t_SL g3017 ( 
.A(n_2886),
.Y(n_3017)
);

OR2x2_ASAP7_75t_L g3018 ( 
.A(n_2840),
.B(n_247),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2893),
.Y(n_3019)
);

CKINVDCx16_ASAP7_75t_R g3020 ( 
.A(n_2847),
.Y(n_3020)
);

AOI21xp5_ASAP7_75t_SL g3021 ( 
.A1(n_2939),
.A2(n_247),
.B(n_248),
.Y(n_3021)
);

INVx3_ASAP7_75t_SL g3022 ( 
.A(n_2850),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2898),
.Y(n_3023)
);

OR2x2_ASAP7_75t_L g3024 ( 
.A(n_2848),
.B(n_248),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2851),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2853),
.Y(n_3026)
);

OR2x2_ASAP7_75t_L g3027 ( 
.A(n_2854),
.B(n_249),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2861),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2863),
.B(n_249),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2829),
.Y(n_3030)
);

AND2x4_ASAP7_75t_SL g3031 ( 
.A(n_2875),
.B(n_250),
.Y(n_3031)
);

HB1xp67_ASAP7_75t_L g3032 ( 
.A(n_2870),
.Y(n_3032)
);

INVx1_ASAP7_75t_L g3033 ( 
.A(n_2871),
.Y(n_3033)
);

INVx1_ASAP7_75t_SL g3034 ( 
.A(n_2837),
.Y(n_3034)
);

INVx2_ASAP7_75t_L g3035 ( 
.A(n_2876),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2879),
.Y(n_3036)
);

INVx4_ASAP7_75t_L g3037 ( 
.A(n_2856),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2882),
.B(n_251),
.Y(n_3038)
);

AND2x2_ASAP7_75t_L g3039 ( 
.A(n_2887),
.B(n_251),
.Y(n_3039)
);

INVx1_ASAP7_75t_SL g3040 ( 
.A(n_2949),
.Y(n_3040)
);

INVx3_ASAP7_75t_L g3041 ( 
.A(n_2835),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2815),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_L g3043 ( 
.A1(n_2939),
.A2(n_256),
.B1(n_253),
.B2(n_255),
.Y(n_3043)
);

INVx1_ASAP7_75t_SL g3044 ( 
.A(n_2950),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2816),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2914),
.B(n_253),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2919),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2921),
.B(n_255),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2922),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2925),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2927),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2818),
.B(n_256),
.Y(n_3052)
);

OR2x2_ASAP7_75t_L g3053 ( 
.A(n_2934),
.B(n_257),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2940),
.B(n_257),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2943),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2953),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2842),
.Y(n_3057)
);

OR2x6_ASAP7_75t_L g3058 ( 
.A(n_2933),
.B(n_258),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2867),
.B(n_259),
.Y(n_3059)
);

OR2x2_ASAP7_75t_L g3060 ( 
.A(n_2897),
.B(n_259),
.Y(n_3060)
);

BUFx2_ASAP7_75t_L g3061 ( 
.A(n_2906),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2916),
.B(n_2907),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_2908),
.B(n_260),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2912),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2835),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2873),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2824),
.B(n_260),
.Y(n_3067)
);

INVx3_ASAP7_75t_L g3068 ( 
.A(n_2831),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_L g3069 ( 
.A(n_2824),
.B(n_261),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2833),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_2860),
.B(n_261),
.Y(n_3071)
);

INVxp67_ASAP7_75t_SL g3072 ( 
.A(n_2828),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2877),
.Y(n_3073)
);

INVx2_ASAP7_75t_L g3074 ( 
.A(n_2843),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_2857),
.Y(n_3075)
);

INVx1_ASAP7_75t_SL g3076 ( 
.A(n_2883),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_2839),
.B(n_262),
.Y(n_3077)
);

OR2x2_ASAP7_75t_L g3078 ( 
.A(n_2902),
.B(n_262),
.Y(n_3078)
);

INVxp33_ASAP7_75t_L g3079 ( 
.A(n_2864),
.Y(n_3079)
);

INVx4_ASAP7_75t_L g3080 ( 
.A(n_2961),
.Y(n_3080)
);

AND2x2_ASAP7_75t_L g3081 ( 
.A(n_2817),
.B(n_264),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2862),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2891),
.B(n_265),
.Y(n_3083)
);

HB1xp67_ASAP7_75t_L g3084 ( 
.A(n_2915),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2917),
.B(n_265),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_L g3086 ( 
.A(n_2918),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2885),
.Y(n_3087)
);

NAND2xp5_ASAP7_75t_L g3088 ( 
.A(n_2923),
.B(n_266),
.Y(n_3088)
);

OAI21xp5_ASAP7_75t_SL g3089 ( 
.A1(n_2930),
.A2(n_267),
.B(n_268),
.Y(n_3089)
);

AOI22xp5_ASAP7_75t_L g3090 ( 
.A1(n_2924),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_3090)
);

INVx1_ASAP7_75t_SL g3091 ( 
.A(n_2844),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2845),
.Y(n_3092)
);

NOR2xp33_ASAP7_75t_L g3093 ( 
.A(n_2942),
.B(n_269),
.Y(n_3093)
);

OAI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_2944),
.A2(n_272),
.B1(n_270),
.B2(n_271),
.Y(n_3094)
);

INVx2_ASAP7_75t_SL g3095 ( 
.A(n_2931),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2932),
.Y(n_3096)
);

INVx1_ASAP7_75t_SL g3097 ( 
.A(n_2951),
.Y(n_3097)
);

AND2x2_ASAP7_75t_L g3098 ( 
.A(n_2941),
.B(n_271),
.Y(n_3098)
);

OAI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2960),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2957),
.B(n_273),
.Y(n_3100)
);

INVx4_ASAP7_75t_L g3101 ( 
.A(n_2959),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2852),
.B(n_274),
.Y(n_3102)
);

INVx1_ASAP7_75t_SL g3103 ( 
.A(n_2929),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2859),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2945),
.Y(n_3105)
);

INVx1_ASAP7_75t_SL g3106 ( 
.A(n_2920),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_2926),
.Y(n_3107)
);

INVx1_ASAP7_75t_L g3108 ( 
.A(n_2958),
.Y(n_3108)
);

NAND2xp33_ASAP7_75t_SL g3109 ( 
.A(n_2826),
.B(n_275),
.Y(n_3109)
);

INVx2_ASAP7_75t_L g3110 ( 
.A(n_2946),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2880),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_2841),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2874),
.B(n_275),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_2841),
.Y(n_3114)
);

AOI22xp5_ASAP7_75t_L g3115 ( 
.A1(n_2939),
.A2(n_279),
.B1(n_276),
.B2(n_278),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2936),
.Y(n_3116)
);

OAI21x1_ASAP7_75t_L g3117 ( 
.A1(n_2901),
.A2(n_276),
.B(n_278),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_2880),
.Y(n_3118)
);

AOI22xp33_ASAP7_75t_L g3119 ( 
.A1(n_2939),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_3119)
);

NOR2x1_ASAP7_75t_L g3120 ( 
.A(n_2849),
.B(n_280),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2880),
.Y(n_3121)
);

CKINVDCx16_ASAP7_75t_R g3122 ( 
.A(n_2900),
.Y(n_3122)
);

AND2x2_ASAP7_75t_L g3123 ( 
.A(n_2874),
.B(n_282),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2827),
.B(n_284),
.Y(n_3124)
);

NOR2x1_ASAP7_75t_L g3125 ( 
.A(n_2849),
.B(n_284),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2880),
.Y(n_3126)
);

NOR2x1_ASAP7_75t_L g3127 ( 
.A(n_2849),
.B(n_285),
.Y(n_3127)
);

OR2x2_ASAP7_75t_L g3128 ( 
.A(n_2825),
.B(n_285),
.Y(n_3128)
);

NOR2x1_ASAP7_75t_L g3129 ( 
.A(n_2849),
.B(n_287),
.Y(n_3129)
);

BUFx2_ASAP7_75t_L g3130 ( 
.A(n_2936),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2874),
.B(n_288),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2880),
.Y(n_3132)
);

OAI221xp5_ASAP7_75t_SL g3133 ( 
.A1(n_2844),
.A2(n_290),
.B1(n_288),
.B2(n_289),
.C(n_291),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2880),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2874),
.B(n_289),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2939),
.A2(n_293),
.B1(n_290),
.B2(n_292),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2936),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2880),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2880),
.Y(n_3139)
);

AOI222xp33_ASAP7_75t_L g3140 ( 
.A1(n_2826),
.A2(n_295),
.B1(n_297),
.B2(n_292),
.C1(n_294),
.C2(n_296),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2880),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2830),
.B(n_294),
.Y(n_3142)
);

AOI22xp33_ASAP7_75t_L g3143 ( 
.A1(n_2939),
.A2(n_297),
.B1(n_295),
.B2(n_296),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2830),
.B(n_298),
.Y(n_3144)
);

INVx1_ASAP7_75t_SL g3145 ( 
.A(n_2841),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2874),
.B(n_298),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2880),
.Y(n_3147)
);

INVx4_ASAP7_75t_L g3148 ( 
.A(n_2841),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2830),
.B(n_299),
.Y(n_3149)
);

INVxp67_ASAP7_75t_L g3150 ( 
.A(n_2849),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2874),
.B(n_299),
.Y(n_3151)
);

AND2x2_ASAP7_75t_L g3152 ( 
.A(n_2874),
.B(n_300),
.Y(n_3152)
);

INVx2_ASAP7_75t_L g3153 ( 
.A(n_2936),
.Y(n_3153)
);

NOR2x1p5_ASAP7_75t_L g3154 ( 
.A(n_2827),
.B(n_300),
.Y(n_3154)
);

HB1xp67_ASAP7_75t_L g3155 ( 
.A(n_2936),
.Y(n_3155)
);

INVx1_ASAP7_75t_SL g3156 ( 
.A(n_2841),
.Y(n_3156)
);

INVx2_ASAP7_75t_L g3157 ( 
.A(n_2936),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2880),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2936),
.Y(n_3159)
);

NOR2xp33_ASAP7_75t_L g3160 ( 
.A(n_2827),
.B(n_301),
.Y(n_3160)
);

INVx3_ASAP7_75t_SL g3161 ( 
.A(n_2841),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_2874),
.B(n_302),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2880),
.Y(n_3163)
);

OR2x2_ASAP7_75t_L g3164 ( 
.A(n_2825),
.B(n_302),
.Y(n_3164)
);

HB1xp67_ASAP7_75t_L g3165 ( 
.A(n_2936),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2880),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2936),
.Y(n_3167)
);

HB1xp67_ASAP7_75t_L g3168 ( 
.A(n_2936),
.Y(n_3168)
);

INVx1_ASAP7_75t_SL g3169 ( 
.A(n_2841),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2964),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3111),
.Y(n_3171)
);

INVx1_ASAP7_75t_L g3172 ( 
.A(n_3118),
.Y(n_3172)
);

OAI21xp5_ASAP7_75t_SL g3173 ( 
.A1(n_3079),
.A2(n_305),
.B(n_304),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2976),
.B(n_303),
.Y(n_3174)
);

AND2x2_ASAP7_75t_L g3175 ( 
.A(n_3130),
.B(n_303),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3121),
.Y(n_3176)
);

NAND2x1p5_ASAP7_75t_L g3177 ( 
.A(n_3004),
.B(n_304),
.Y(n_3177)
);

OAI21xp33_ASAP7_75t_L g3178 ( 
.A1(n_3021),
.A2(n_305),
.B(n_306),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2977),
.B(n_306),
.Y(n_3179)
);

OAI21xp33_ASAP7_75t_L g3180 ( 
.A1(n_3115),
.A2(n_307),
.B(n_308),
.Y(n_3180)
);

AOI22xp5_ASAP7_75t_L g3181 ( 
.A1(n_2991),
.A2(n_310),
.B1(n_307),
.B2(n_309),
.Y(n_3181)
);

AOI321xp33_ASAP7_75t_L g3182 ( 
.A1(n_3094),
.A2(n_313),
.A3(n_315),
.B1(n_311),
.B2(n_312),
.C(n_314),
.Y(n_3182)
);

OR2x2_ASAP7_75t_L g3183 ( 
.A(n_2981),
.B(n_312),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_3126),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_3132),
.Y(n_3185)
);

HB1xp67_ASAP7_75t_L g3186 ( 
.A(n_3155),
.Y(n_3186)
);

OR2x2_ASAP7_75t_L g3187 ( 
.A(n_2971),
.B(n_313),
.Y(n_3187)
);

A2O1A1Ixp33_ASAP7_75t_L g3188 ( 
.A1(n_3041),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_3150),
.B(n_3006),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_3134),
.Y(n_3190)
);

NAND3xp33_ASAP7_75t_SL g3191 ( 
.A(n_3034),
.B(n_316),
.C(n_317),
.Y(n_3191)
);

AOI22xp5_ASAP7_75t_L g3192 ( 
.A1(n_2972),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_3192)
);

OAI22xp33_ASAP7_75t_L g3193 ( 
.A1(n_3122),
.A2(n_322),
.B1(n_318),
.B2(n_321),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_3138),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_3011),
.B(n_321),
.Y(n_3195)
);

OAI222xp33_ASAP7_75t_L g3196 ( 
.A1(n_3080),
.A2(n_325),
.B1(n_327),
.B2(n_328),
.C1(n_324),
.C2(n_326),
.Y(n_3196)
);

INVxp67_ASAP7_75t_L g3197 ( 
.A(n_3072),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3139),
.Y(n_3198)
);

INVx2_ASAP7_75t_L g3199 ( 
.A(n_3116),
.Y(n_3199)
);

OAI322xp33_ASAP7_75t_L g3200 ( 
.A1(n_3101),
.A2(n_330),
.A3(n_329),
.B1(n_326),
.B2(n_323),
.C1(n_325),
.C2(n_327),
.Y(n_3200)
);

INVx1_ASAP7_75t_SL g3201 ( 
.A(n_3161),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3141),
.Y(n_3202)
);

OAI21xp33_ASAP7_75t_SL g3203 ( 
.A1(n_2966),
.A2(n_323),
.B(n_331),
.Y(n_3203)
);

INVx3_ASAP7_75t_L g3204 ( 
.A(n_3148),
.Y(n_3204)
);

AOI21xp5_ASAP7_75t_L g3205 ( 
.A1(n_3109),
.A2(n_331),
.B(n_332),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_3014),
.B(n_3030),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_3147),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_L g3208 ( 
.A(n_3037),
.B(n_333),
.Y(n_3208)
);

AO21x1_ASAP7_75t_L g3209 ( 
.A1(n_3142),
.A2(n_333),
.B(n_334),
.Y(n_3209)
);

AOI22xp5_ASAP7_75t_L g3210 ( 
.A1(n_3084),
.A2(n_337),
.B1(n_334),
.B2(n_336),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_L g3211 ( 
.A(n_3061),
.B(n_336),
.Y(n_3211)
);

OAI222xp33_ASAP7_75t_L g3212 ( 
.A1(n_3086),
.A2(n_339),
.B1(n_342),
.B2(n_344),
.C1(n_338),
.C2(n_340),
.Y(n_3212)
);

OR2x2_ASAP7_75t_L g3213 ( 
.A(n_3137),
.B(n_337),
.Y(n_3213)
);

AOI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_3104),
.A2(n_342),
.B1(n_338),
.B2(n_340),
.Y(n_3214)
);

NAND2xp5_ASAP7_75t_L g3215 ( 
.A(n_3001),
.B(n_345),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_3144),
.A2(n_345),
.B(n_347),
.Y(n_3216)
);

INVx1_ASAP7_75t_L g3217 ( 
.A(n_3158),
.Y(n_3217)
);

AOI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_3105),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.Y(n_3218)
);

AO22x1_ASAP7_75t_L g3219 ( 
.A1(n_3022),
.A2(n_351),
.B1(n_348),
.B2(n_350),
.Y(n_3219)
);

OAI221xp5_ASAP7_75t_L g3220 ( 
.A1(n_3089),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.C(n_353),
.Y(n_3220)
);

OA211x2_ASAP7_75t_L g3221 ( 
.A1(n_3149),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_3065),
.B(n_355),
.Y(n_3222)
);

NAND4xp75_ASAP7_75t_L g3223 ( 
.A(n_3120),
.B(n_358),
.C(n_355),
.D(n_357),
.Y(n_3223)
);

AOI21xp33_ASAP7_75t_L g3224 ( 
.A1(n_3087),
.A2(n_357),
.B(n_358),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3163),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3166),
.Y(n_3226)
);

NAND2xp5_ASAP7_75t_L g3227 ( 
.A(n_3032),
.B(n_359),
.Y(n_3227)
);

INVx1_ASAP7_75t_SL g3228 ( 
.A(n_2989),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3106),
.B(n_360),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2984),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3153),
.Y(n_3231)
);

NAND2xp33_ASAP7_75t_R g3232 ( 
.A(n_3107),
.B(n_360),
.Y(n_3232)
);

OA21x2_ASAP7_75t_L g3233 ( 
.A1(n_3157),
.A2(n_361),
.B(n_362),
.Y(n_3233)
);

OAI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3075),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_3234)
);

NAND2xp33_ASAP7_75t_L g3235 ( 
.A(n_3125),
.B(n_364),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3057),
.B(n_364),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_3045),
.B(n_365),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3047),
.B(n_365),
.Y(n_3238)
);

OR2x2_ASAP7_75t_L g3239 ( 
.A(n_3159),
.B(n_366),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_2974),
.B(n_366),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3049),
.B(n_368),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3167),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_3064),
.B(n_368),
.Y(n_3243)
);

OAI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3127),
.A2(n_369),
.B(n_370),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_3068),
.A2(n_371),
.B1(n_369),
.B2(n_370),
.Y(n_3245)
);

OAI21xp33_ASAP7_75t_SL g3246 ( 
.A1(n_3017),
.A2(n_371),
.B(n_372),
.Y(n_3246)
);

AOI211x1_ASAP7_75t_SL g3247 ( 
.A1(n_3099),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_3247)
);

AOI22xp5_ASAP7_75t_L g3248 ( 
.A1(n_3097),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2986),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_2987),
.Y(n_3250)
);

OAI22xp5_ASAP7_75t_L g3251 ( 
.A1(n_3095),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_3020),
.B(n_3040),
.Y(n_3252)
);

NOR2xp33_ASAP7_75t_L g3253 ( 
.A(n_2997),
.B(n_3008),
.Y(n_3253)
);

NOR4xp25_ASAP7_75t_L g3254 ( 
.A(n_3067),
.B(n_381),
.C(n_379),
.D(n_380),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_2979),
.B(n_380),
.Y(n_3255)
);

INVx1_ASAP7_75t_SL g3256 ( 
.A(n_3044),
.Y(n_3256)
);

NOR2xp33_ASAP7_75t_L g3257 ( 
.A(n_2965),
.B(n_383),
.Y(n_3257)
);

CKINVDCx20_ASAP7_75t_R g3258 ( 
.A(n_2993),
.Y(n_3258)
);

OAI221xp5_ASAP7_75t_L g3259 ( 
.A1(n_3015),
.A2(n_385),
.B1(n_383),
.B2(n_384),
.C(n_386),
.Y(n_3259)
);

OAI22xp33_ASAP7_75t_L g3260 ( 
.A1(n_3090),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_3260)
);

NOR2x1_ASAP7_75t_L g3261 ( 
.A(n_3129),
.B(n_387),
.Y(n_3261)
);

OAI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_2973),
.A2(n_387),
.B(n_388),
.Y(n_3262)
);

AOI21xp33_ASAP7_75t_SL g3263 ( 
.A1(n_3096),
.A2(n_388),
.B(n_389),
.Y(n_3263)
);

OAI21xp33_ASAP7_75t_SL g3264 ( 
.A1(n_3165),
.A2(n_389),
.B(n_390),
.Y(n_3264)
);

AOI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3069),
.A2(n_390),
.B(n_391),
.Y(n_3265)
);

OAI211xp5_ASAP7_75t_L g3266 ( 
.A1(n_3043),
.A2(n_394),
.B(n_392),
.C(n_393),
.Y(n_3266)
);

AOI22xp5_ASAP7_75t_L g3267 ( 
.A1(n_3091),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.Y(n_3267)
);

INVx1_ASAP7_75t_L g3268 ( 
.A(n_3168),
.Y(n_3268)
);

AOI221x1_ASAP7_75t_L g3269 ( 
.A1(n_3088),
.A2(n_3100),
.B1(n_3085),
.B2(n_3098),
.C(n_3081),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2968),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2967),
.Y(n_3271)
);

AND2x4_ASAP7_75t_L g3272 ( 
.A(n_3003),
.B(n_395),
.Y(n_3272)
);

OAI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3093),
.A2(n_396),
.B(n_397),
.Y(n_3273)
);

OR2x2_ASAP7_75t_L g3274 ( 
.A(n_3025),
.B(n_396),
.Y(n_3274)
);

NOR3xp33_ASAP7_75t_L g3275 ( 
.A(n_3133),
.B(n_397),
.C(n_398),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3092),
.B(n_399),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2988),
.Y(n_3277)
);

OR2x2_ASAP7_75t_L g3278 ( 
.A(n_3026),
.B(n_399),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2995),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3019),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3023),
.Y(n_3281)
);

NAND3xp33_ASAP7_75t_SL g3282 ( 
.A(n_3119),
.B(n_400),
.C(n_401),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3028),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_3076),
.B(n_3035),
.Y(n_3284)
);

HB1xp67_ASAP7_75t_L g3285 ( 
.A(n_2985),
.Y(n_3285)
);

AND2x2_ASAP7_75t_L g3286 ( 
.A(n_3113),
.B(n_400),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_2996),
.Y(n_3287)
);

AOI221xp5_ASAP7_75t_L g3288 ( 
.A1(n_3103),
.A2(n_3073),
.B1(n_3108),
.B2(n_3082),
.C(n_3136),
.Y(n_3288)
);

INVx2_ASAP7_75t_SL g3289 ( 
.A(n_3154),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_3123),
.B(n_401),
.Y(n_3290)
);

NOR2x1_ASAP7_75t_L g3291 ( 
.A(n_2975),
.B(n_402),
.Y(n_3291)
);

AND2x2_ASAP7_75t_L g3292 ( 
.A(n_3131),
.B(n_403),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3033),
.Y(n_3293)
);

AOI22xp5_ASAP7_75t_L g3294 ( 
.A1(n_3110),
.A2(n_405),
.B1(n_403),
.B2(n_404),
.Y(n_3294)
);

INVxp67_ASAP7_75t_SL g3295 ( 
.A(n_3066),
.Y(n_3295)
);

INVxp67_ASAP7_75t_SL g3296 ( 
.A(n_3070),
.Y(n_3296)
);

OR2x2_ASAP7_75t_L g3297 ( 
.A(n_2970),
.B(n_405),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3036),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3042),
.B(n_406),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3050),
.Y(n_3300)
);

INVxp67_ASAP7_75t_SL g3301 ( 
.A(n_3074),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3051),
.B(n_406),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3055),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3056),
.Y(n_3304)
);

OR2x2_ASAP7_75t_L g3305 ( 
.A(n_3128),
.B(n_3164),
.Y(n_3305)
);

NAND3xp33_ASAP7_75t_SL g3306 ( 
.A(n_3143),
.B(n_407),
.C(n_408),
.Y(n_3306)
);

OAI211xp5_ASAP7_75t_L g3307 ( 
.A1(n_3140),
.A2(n_411),
.B(n_407),
.C(n_409),
.Y(n_3307)
);

OAI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_3083),
.A2(n_409),
.B(n_412),
.Y(n_3308)
);

OAI21xp33_ASAP7_75t_SL g3309 ( 
.A1(n_3135),
.A2(n_413),
.B(n_414),
.Y(n_3309)
);

OAI21xp33_ASAP7_75t_L g3310 ( 
.A1(n_3102),
.A2(n_415),
.B(n_416),
.Y(n_3310)
);

INVx2_ASAP7_75t_SL g3311 ( 
.A(n_2983),
.Y(n_3311)
);

OAI22xp33_ASAP7_75t_L g3312 ( 
.A1(n_3058),
.A2(n_417),
.B1(n_415),
.B2(n_416),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2969),
.Y(n_3313)
);

AOI21xp33_ASAP7_75t_L g3314 ( 
.A1(n_3078),
.A2(n_417),
.B(n_419),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3146),
.B(n_419),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3000),
.Y(n_3316)
);

NOR2xp33_ASAP7_75t_L g3317 ( 
.A(n_3060),
.B(n_421),
.Y(n_3317)
);

AOI22xp5_ASAP7_75t_L g3318 ( 
.A1(n_3077),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3318)
);

NAND2xp33_ASAP7_75t_L g3319 ( 
.A(n_2992),
.B(n_422),
.Y(n_3319)
);

AND2x2_ASAP7_75t_L g3320 ( 
.A(n_3201),
.B(n_3151),
.Y(n_3320)
);

NOR2xp33_ASAP7_75t_SL g3321 ( 
.A(n_3178),
.B(n_2963),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3186),
.Y(n_3322)
);

AND2x2_ASAP7_75t_L g3323 ( 
.A(n_3204),
.B(n_3152),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3269),
.B(n_3162),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3170),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3295),
.B(n_3062),
.Y(n_3326)
);

NAND2x1p5_ASAP7_75t_L g3327 ( 
.A(n_3261),
.B(n_2983),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3204),
.B(n_3112),
.Y(n_3328)
);

AND2x2_ASAP7_75t_L g3329 ( 
.A(n_3296),
.B(n_3114),
.Y(n_3329)
);

BUFx2_ASAP7_75t_L g3330 ( 
.A(n_3289),
.Y(n_3330)
);

INVx2_ASAP7_75t_SL g3331 ( 
.A(n_3272),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3301),
.B(n_3002),
.Y(n_3332)
);

HB1xp67_ASAP7_75t_L g3333 ( 
.A(n_3197),
.Y(n_3333)
);

INVxp67_ASAP7_75t_L g3334 ( 
.A(n_3232),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_SL g3335 ( 
.A(n_3256),
.B(n_3169),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3171),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_3228),
.B(n_3145),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3216),
.B(n_3010),
.Y(n_3338)
);

INVx3_ASAP7_75t_L g3339 ( 
.A(n_3272),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3172),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_3176),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3184),
.Y(n_3342)
);

AOI222xp33_ASAP7_75t_L g3343 ( 
.A1(n_3288),
.A2(n_3071),
.B1(n_3031),
.B2(n_2994),
.C1(n_3160),
.C2(n_3124),
.Y(n_3343)
);

NOR2x1_ASAP7_75t_L g3344 ( 
.A(n_3191),
.B(n_3058),
.Y(n_3344)
);

NAND3xp33_ASAP7_75t_L g3345 ( 
.A(n_3275),
.B(n_2982),
.C(n_3016),
.Y(n_3345)
);

HB1xp67_ASAP7_75t_L g3346 ( 
.A(n_3233),
.Y(n_3346)
);

NAND2x1_ASAP7_75t_SL g3347 ( 
.A(n_3291),
.B(n_2980),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3253),
.B(n_3156),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3209),
.B(n_3039),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3252),
.B(n_3013),
.Y(n_3350)
);

OR2x2_ASAP7_75t_L g3351 ( 
.A(n_3268),
.B(n_3053),
.Y(n_3351)
);

OR2x2_ASAP7_75t_L g3352 ( 
.A(n_3206),
.B(n_3024),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3311),
.B(n_3046),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3185),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3203),
.B(n_3048),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3316),
.B(n_3063),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_3317),
.B(n_3054),
.Y(n_3357)
);

INVx2_ASAP7_75t_SL g3358 ( 
.A(n_3258),
.Y(n_3358)
);

NOR2xp33_ASAP7_75t_L g3359 ( 
.A(n_3246),
.B(n_3027),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3190),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3265),
.B(n_3059),
.Y(n_3361)
);

INVx2_ASAP7_75t_L g3362 ( 
.A(n_3187),
.Y(n_3362)
);

INVx2_ASAP7_75t_L g3363 ( 
.A(n_3213),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3194),
.Y(n_3364)
);

OAI31xp33_ASAP7_75t_SL g3365 ( 
.A1(n_3307),
.A2(n_3180),
.A3(n_3260),
.B(n_3244),
.Y(n_3365)
);

AND2x2_ASAP7_75t_SL g3366 ( 
.A(n_3235),
.B(n_2999),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_3313),
.B(n_3005),
.Y(n_3367)
);

OR2x2_ASAP7_75t_L g3368 ( 
.A(n_3189),
.B(n_2990),
.Y(n_3368)
);

AOI22xp33_ASAP7_75t_L g3369 ( 
.A1(n_3282),
.A2(n_2998),
.B1(n_3038),
.B2(n_3029),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3199),
.B(n_3018),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3239),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_3254),
.B(n_3009),
.Y(n_3372)
);

NOR2xp33_ASAP7_75t_L g3373 ( 
.A(n_3305),
.B(n_3052),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_3198),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_3219),
.B(n_3007),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3202),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3264),
.B(n_3012),
.Y(n_3377)
);

INVx3_ASAP7_75t_L g3378 ( 
.A(n_3177),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3231),
.B(n_2978),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3242),
.B(n_3117),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3309),
.B(n_424),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_3284),
.B(n_3182),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_SL g3383 ( 
.A(n_3205),
.B(n_424),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3207),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3175),
.B(n_425),
.Y(n_3385)
);

INVx1_ASAP7_75t_L g3386 ( 
.A(n_3217),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3225),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3183),
.B(n_3287),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3179),
.B(n_426),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3294),
.B(n_3174),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3226),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3230),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3318),
.B(n_426),
.Y(n_3393)
);

OR2x2_ASAP7_75t_L g3394 ( 
.A(n_3270),
.B(n_427),
.Y(n_3394)
);

OAI21xp5_ASAP7_75t_SL g3395 ( 
.A1(n_3173),
.A2(n_427),
.B(n_428),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3300),
.B(n_428),
.Y(n_3396)
);

AND2x2_ASAP7_75t_L g3397 ( 
.A(n_3285),
.B(n_430),
.Y(n_3397)
);

AOI22xp33_ASAP7_75t_SL g3398 ( 
.A1(n_3273),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3255),
.B(n_431),
.Y(n_3399)
);

NOR2x1_ASAP7_75t_L g3400 ( 
.A(n_3233),
.B(n_432),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3303),
.B(n_433),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_L g3402 ( 
.A(n_3195),
.B(n_435),
.Y(n_3402)
);

NAND2x1p5_ASAP7_75t_L g3403 ( 
.A(n_3240),
.B(n_435),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3304),
.B(n_436),
.Y(n_3404)
);

AND2x4_ASAP7_75t_SL g3405 ( 
.A(n_3286),
.B(n_436),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3283),
.Y(n_3406)
);

OR2x2_ASAP7_75t_L g3407 ( 
.A(n_3293),
.B(n_437),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3298),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3229),
.B(n_437),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3277),
.B(n_438),
.Y(n_3410)
);

OAI22xp5_ASAP7_75t_L g3411 ( 
.A1(n_3220),
.A2(n_441),
.B1(n_439),
.B2(n_440),
.Y(n_3411)
);

AND2x2_ASAP7_75t_L g3412 ( 
.A(n_3290),
.B(n_439),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3279),
.B(n_440),
.Y(n_3413)
);

NAND2x1_ASAP7_75t_SL g3414 ( 
.A(n_3181),
.B(n_442),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_3280),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3215),
.B(n_442),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3281),
.B(n_443),
.Y(n_3417)
);

INVx1_ASAP7_75t_SL g3418 ( 
.A(n_3292),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3208),
.B(n_3222),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3333),
.Y(n_3420)
);

NOR2xp33_ASAP7_75t_L g3421 ( 
.A(n_3334),
.B(n_3243),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3346),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3358),
.Y(n_3423)
);

CKINVDCx20_ASAP7_75t_R g3424 ( 
.A(n_3335),
.Y(n_3424)
);

INVx2_ASAP7_75t_SL g3425 ( 
.A(n_3339),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_3330),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3322),
.Y(n_3427)
);

INVx2_ASAP7_75t_L g3428 ( 
.A(n_3328),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3397),
.Y(n_3429)
);

HB1xp67_ASAP7_75t_L g3430 ( 
.A(n_3327),
.Y(n_3430)
);

INVx5_ASAP7_75t_L g3431 ( 
.A(n_3339),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3394),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3407),
.Y(n_3433)
);

BUFx4f_ASAP7_75t_SL g3434 ( 
.A(n_3399),
.Y(n_3434)
);

INVx2_ASAP7_75t_L g3435 ( 
.A(n_3378),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3362),
.Y(n_3436)
);

CKINVDCx6p67_ASAP7_75t_R g3437 ( 
.A(n_3412),
.Y(n_3437)
);

CKINVDCx20_ASAP7_75t_R g3438 ( 
.A(n_3348),
.Y(n_3438)
);

INVx1_ASAP7_75t_SL g3439 ( 
.A(n_3347),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3363),
.Y(n_3440)
);

BUFx2_ASAP7_75t_L g3441 ( 
.A(n_3378),
.Y(n_3441)
);

INVx2_ASAP7_75t_SL g3442 ( 
.A(n_3331),
.Y(n_3442)
);

INVx2_ASAP7_75t_L g3443 ( 
.A(n_3320),
.Y(n_3443)
);

BUFx2_ASAP7_75t_L g3444 ( 
.A(n_3329),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3371),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3388),
.Y(n_3446)
);

INVx1_ASAP7_75t_SL g3447 ( 
.A(n_3366),
.Y(n_3447)
);

INVxp33_ASAP7_75t_SL g3448 ( 
.A(n_3337),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3356),
.Y(n_3449)
);

XNOR2xp5_ASAP7_75t_L g3450 ( 
.A(n_3344),
.B(n_3192),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3325),
.Y(n_3451)
);

INVx1_ASAP7_75t_SL g3452 ( 
.A(n_3405),
.Y(n_3452)
);

INVx2_ASAP7_75t_SL g3453 ( 
.A(n_3323),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3336),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3340),
.Y(n_3455)
);

INVxp33_ASAP7_75t_SL g3456 ( 
.A(n_3321),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3341),
.Y(n_3457)
);

CKINVDCx20_ASAP7_75t_R g3458 ( 
.A(n_3355),
.Y(n_3458)
);

INVx2_ASAP7_75t_L g3459 ( 
.A(n_3403),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3342),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3354),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_3370),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_3360),
.Y(n_3463)
);

HB1xp67_ASAP7_75t_L g3464 ( 
.A(n_3400),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3367),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3364),
.Y(n_3466)
);

INVxp33_ASAP7_75t_SL g3467 ( 
.A(n_3359),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_3351),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3374),
.Y(n_3469)
);

NOR2xp33_ASAP7_75t_L g3470 ( 
.A(n_3375),
.B(n_3299),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3376),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3384),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3386),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3365),
.B(n_3263),
.Y(n_3474)
);

INVx2_ASAP7_75t_L g3475 ( 
.A(n_3418),
.Y(n_3475)
);

NOR2x1_ASAP7_75t_L g3476 ( 
.A(n_3345),
.B(n_3223),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_3350),
.Y(n_3477)
);

INVx2_ASAP7_75t_SL g3478 ( 
.A(n_3414),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3380),
.Y(n_3479)
);

CKINVDCx20_ASAP7_75t_R g3480 ( 
.A(n_3382),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3387),
.Y(n_3481)
);

INVxp67_ASAP7_75t_L g3482 ( 
.A(n_3349),
.Y(n_3482)
);

BUFx2_ASAP7_75t_L g3483 ( 
.A(n_3326),
.Y(n_3483)
);

INVx1_ASAP7_75t_SL g3484 ( 
.A(n_3377),
.Y(n_3484)
);

INVx2_ASAP7_75t_L g3485 ( 
.A(n_3353),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3391),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3343),
.B(n_3193),
.Y(n_3487)
);

INVxp67_ASAP7_75t_L g3488 ( 
.A(n_3324),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3392),
.Y(n_3489)
);

XNOR2x1_ASAP7_75t_L g3490 ( 
.A(n_3411),
.B(n_3308),
.Y(n_3490)
);

AND2x2_ASAP7_75t_L g3491 ( 
.A(n_3373),
.B(n_3249),
.Y(n_3491)
);

CKINVDCx6p67_ASAP7_75t_R g3492 ( 
.A(n_3409),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3406),
.Y(n_3493)
);

NAND2x1_ASAP7_75t_SL g3494 ( 
.A(n_3408),
.B(n_3210),
.Y(n_3494)
);

INVx2_ASAP7_75t_SL g3495 ( 
.A(n_3368),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3415),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_SL g3497 ( 
.A(n_3361),
.B(n_3312),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3396),
.Y(n_3498)
);

INVxp67_ASAP7_75t_L g3499 ( 
.A(n_3383),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3372),
.B(n_3237),
.Y(n_3500)
);

CKINVDCx5p33_ASAP7_75t_R g3501 ( 
.A(n_3402),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_3401),
.Y(n_3502)
);

INVxp33_ASAP7_75t_L g3503 ( 
.A(n_3332),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3404),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3410),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_3413),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3417),
.Y(n_3507)
);

AND2x4_ASAP7_75t_SL g3508 ( 
.A(n_3369),
.B(n_3257),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3352),
.Y(n_3509)
);

HB1xp67_ASAP7_75t_L g3510 ( 
.A(n_3379),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3381),
.Y(n_3511)
);

INVx1_ASAP7_75t_SL g3512 ( 
.A(n_3385),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3389),
.Y(n_3513)
);

INVxp67_ASAP7_75t_L g3514 ( 
.A(n_3419),
.Y(n_3514)
);

INVxp67_ASAP7_75t_L g3515 ( 
.A(n_3357),
.Y(n_3515)
);

INVx1_ASAP7_75t_L g3516 ( 
.A(n_3416),
.Y(n_3516)
);

INVxp67_ASAP7_75t_L g3517 ( 
.A(n_3338),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3393),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3390),
.Y(n_3519)
);

INVxp33_ASAP7_75t_SL g3520 ( 
.A(n_3395),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3398),
.Y(n_3521)
);

INVx1_ASAP7_75t_SL g3522 ( 
.A(n_3347),
.Y(n_3522)
);

INVxp67_ASAP7_75t_L g3523 ( 
.A(n_3330),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3358),
.Y(n_3524)
);

OAI221xp5_ASAP7_75t_L g3525 ( 
.A1(n_3494),
.A2(n_3245),
.B1(n_3310),
.B2(n_3262),
.C(n_3218),
.Y(n_3525)
);

INVx1_ASAP7_75t_SL g3526 ( 
.A(n_3438),
.Y(n_3526)
);

NOR2x1_ASAP7_75t_L g3527 ( 
.A(n_3476),
.B(n_3196),
.Y(n_3527)
);

AOI211xp5_ASAP7_75t_L g3528 ( 
.A1(n_3474),
.A2(n_3212),
.B(n_3200),
.C(n_3234),
.Y(n_3528)
);

NAND4xp25_ASAP7_75t_L g3529 ( 
.A(n_3447),
.B(n_3221),
.C(n_3247),
.D(n_3188),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3464),
.Y(n_3530)
);

NAND3xp33_ASAP7_75t_L g3531 ( 
.A(n_3488),
.B(n_3266),
.C(n_3319),
.Y(n_3531)
);

NAND2xp33_ASAP7_75t_L g3532 ( 
.A(n_3478),
.B(n_3274),
.Y(n_3532)
);

NAND3xp33_ASAP7_75t_L g3533 ( 
.A(n_3482),
.B(n_3259),
.C(n_3214),
.Y(n_3533)
);

NOR3xp33_ASAP7_75t_L g3534 ( 
.A(n_3487),
.B(n_3500),
.C(n_3421),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3444),
.B(n_3250),
.Y(n_3535)
);

OR2x2_ASAP7_75t_L g3536 ( 
.A(n_3484),
.B(n_3271),
.Y(n_3536)
);

NOR3xp33_ASAP7_75t_L g3537 ( 
.A(n_3497),
.B(n_3314),
.C(n_3224),
.Y(n_3537)
);

NOR3xp33_ASAP7_75t_L g3538 ( 
.A(n_3514),
.B(n_3306),
.C(n_3251),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_3448),
.B(n_3248),
.Y(n_3539)
);

NAND3xp33_ASAP7_75t_L g3540 ( 
.A(n_3450),
.B(n_3267),
.C(n_3276),
.Y(n_3540)
);

NAND3xp33_ASAP7_75t_L g3541 ( 
.A(n_3431),
.B(n_3211),
.C(n_3227),
.Y(n_3541)
);

NOR3xp33_ASAP7_75t_L g3542 ( 
.A(n_3523),
.B(n_3236),
.C(n_3302),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_SL g3543 ( 
.A(n_3456),
.B(n_3278),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3422),
.Y(n_3544)
);

OAI211xp5_ASAP7_75t_L g3545 ( 
.A1(n_3439),
.A2(n_3241),
.B(n_3238),
.C(n_3315),
.Y(n_3545)
);

NAND4xp25_ASAP7_75t_L g3546 ( 
.A(n_3467),
.B(n_3297),
.C(n_445),
.D(n_443),
.Y(n_3546)
);

NAND4xp25_ASAP7_75t_L g3547 ( 
.A(n_3470),
.B(n_447),
.C(n_444),
.D(n_446),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3452),
.B(n_444),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3425),
.B(n_446),
.Y(n_3549)
);

OAI211xp5_ASAP7_75t_SL g3550 ( 
.A1(n_3517),
.A2(n_449),
.B(n_447),
.C(n_448),
.Y(n_3550)
);

NAND4xp25_ASAP7_75t_SL g3551 ( 
.A(n_3522),
.B(n_3480),
.C(n_3424),
.D(n_3521),
.Y(n_3551)
);

OR2x2_ASAP7_75t_L g3552 ( 
.A(n_3443),
.B(n_448),
.Y(n_3552)
);

NAND3xp33_ASAP7_75t_L g3553 ( 
.A(n_3431),
.B(n_449),
.C(n_450),
.Y(n_3553)
);

A2O1A1Ixp33_ASAP7_75t_L g3554 ( 
.A1(n_3499),
.A2(n_452),
.B(n_450),
.C(n_451),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_SL g3555 ( 
.A(n_3431),
.B(n_452),
.Y(n_3555)
);

NOR3x1_ASAP7_75t_SL g3556 ( 
.A(n_3430),
.B(n_453),
.C(n_454),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3426),
.B(n_453),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3420),
.Y(n_3558)
);

OAI221xp5_ASAP7_75t_L g3559 ( 
.A1(n_3490),
.A2(n_457),
.B1(n_455),
.B2(n_456),
.C(n_459),
.Y(n_3559)
);

A2O1A1Ixp33_ASAP7_75t_L g3560 ( 
.A1(n_3508),
.A2(n_457),
.B(n_455),
.C(n_456),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3475),
.Y(n_3561)
);

AOI211xp5_ASAP7_75t_L g3562 ( 
.A1(n_3503),
.A2(n_463),
.B(n_460),
.C(n_462),
.Y(n_3562)
);

NOR2x1_ASAP7_75t_L g3563 ( 
.A(n_3441),
.B(n_460),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3442),
.B(n_464),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_SL g3565 ( 
.A(n_3434),
.B(n_465),
.Y(n_3565)
);

A2O1A1Ixp33_ASAP7_75t_L g3566 ( 
.A1(n_3518),
.A2(n_467),
.B(n_465),
.C(n_466),
.Y(n_3566)
);

O2A1O1Ixp33_ASAP7_75t_L g3567 ( 
.A1(n_3520),
.A2(n_3519),
.B(n_3511),
.C(n_3510),
.Y(n_3567)
);

AOI211xp5_ASAP7_75t_L g3568 ( 
.A1(n_3423),
.A2(n_3524),
.B(n_3435),
.C(n_3428),
.Y(n_3568)
);

OA21x2_ASAP7_75t_L g3569 ( 
.A1(n_3427),
.A2(n_467),
.B(n_468),
.Y(n_3569)
);

AOI21xp5_ASAP7_75t_L g3570 ( 
.A1(n_3458),
.A2(n_468),
.B(n_469),
.Y(n_3570)
);

NOR3x1_ASAP7_75t_L g3571 ( 
.A(n_3453),
.B(n_469),
.C(n_470),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3437),
.B(n_3477),
.Y(n_3572)
);

NOR2xp67_ASAP7_75t_L g3573 ( 
.A(n_3495),
.B(n_470),
.Y(n_3573)
);

NAND4xp25_ASAP7_75t_SL g3574 ( 
.A(n_3449),
.B(n_3512),
.C(n_3429),
.D(n_3465),
.Y(n_3574)
);

AOI211xp5_ASAP7_75t_L g3575 ( 
.A1(n_3446),
.A2(n_473),
.B(n_471),
.C(n_472),
.Y(n_3575)
);

NOR2xp33_ASAP7_75t_L g3576 ( 
.A(n_3459),
.B(n_473),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_3501),
.A2(n_474),
.B(n_475),
.Y(n_3577)
);

OAI211xp5_ASAP7_75t_SL g3578 ( 
.A1(n_3515),
.A2(n_3509),
.B(n_3485),
.C(n_3468),
.Y(n_3578)
);

NOR2xp67_ASAP7_75t_L g3579 ( 
.A(n_3462),
.B(n_474),
.Y(n_3579)
);

NOR4xp25_ASAP7_75t_L g3580 ( 
.A(n_3436),
.B(n_477),
.C(n_475),
.D(n_476),
.Y(n_3580)
);

NAND4xp25_ASAP7_75t_L g3581 ( 
.A(n_3483),
.B(n_3445),
.C(n_3440),
.D(n_3491),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3432),
.B(n_476),
.Y(n_3582)
);

NOR3xp33_ASAP7_75t_L g3583 ( 
.A(n_3498),
.B(n_477),
.C(n_478),
.Y(n_3583)
);

NOR3xp33_ASAP7_75t_SL g3584 ( 
.A(n_3502),
.B(n_479),
.C(n_480),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3433),
.Y(n_3585)
);

XOR2x2_ASAP7_75t_L g3586 ( 
.A(n_3516),
.B(n_480),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3513),
.A2(n_482),
.B(n_483),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3451),
.Y(n_3588)
);

AOI211xp5_ASAP7_75t_L g3589 ( 
.A1(n_3479),
.A2(n_484),
.B(n_482),
.C(n_483),
.Y(n_3589)
);

OAI32xp33_ASAP7_75t_L g3590 ( 
.A1(n_3504),
.A2(n_486),
.A3(n_484),
.B1(n_485),
.B2(n_487),
.Y(n_3590)
);

BUFx3_ASAP7_75t_L g3591 ( 
.A(n_3492),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_L g3592 ( 
.A(n_3505),
.B(n_485),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3506),
.B(n_489),
.Y(n_3593)
);

AOI31xp33_ASAP7_75t_L g3594 ( 
.A1(n_3507),
.A2(n_491),
.A3(n_489),
.B(n_490),
.Y(n_3594)
);

OAI21xp33_ASAP7_75t_L g3595 ( 
.A1(n_3454),
.A2(n_491),
.B(n_492),
.Y(n_3595)
);

OAI221xp5_ASAP7_75t_L g3596 ( 
.A1(n_3527),
.A2(n_3460),
.B1(n_3461),
.B2(n_3457),
.C(n_3455),
.Y(n_3596)
);

OAI21xp33_ASAP7_75t_SL g3597 ( 
.A1(n_3526),
.A2(n_3466),
.B(n_3463),
.Y(n_3597)
);

AOI211xp5_ASAP7_75t_L g3598 ( 
.A1(n_3531),
.A2(n_3471),
.B(n_3472),
.C(n_3469),
.Y(n_3598)
);

NAND3xp33_ASAP7_75t_SL g3599 ( 
.A(n_3528),
.B(n_3481),
.C(n_3473),
.Y(n_3599)
);

AOI32xp33_ASAP7_75t_L g3600 ( 
.A1(n_3537),
.A2(n_3493),
.A3(n_3496),
.B1(n_3489),
.B2(n_3486),
.Y(n_3600)
);

AOI22xp5_ASAP7_75t_L g3601 ( 
.A1(n_3534),
.A2(n_494),
.B1(n_492),
.B2(n_493),
.Y(n_3601)
);

AOI221xp5_ASAP7_75t_L g3602 ( 
.A1(n_3567),
.A2(n_495),
.B1(n_493),
.B2(n_494),
.C(n_496),
.Y(n_3602)
);

AOI221x1_ASAP7_75t_L g3603 ( 
.A1(n_3530),
.A2(n_498),
.B1(n_496),
.B2(n_497),
.C(n_499),
.Y(n_3603)
);

INVx2_ASAP7_75t_L g3604 ( 
.A(n_3591),
.Y(n_3604)
);

NOR2x1_ASAP7_75t_SL g3605 ( 
.A(n_3555),
.B(n_497),
.Y(n_3605)
);

OA211x2_ASAP7_75t_L g3606 ( 
.A1(n_3551),
.A2(n_3539),
.B(n_3574),
.C(n_3543),
.Y(n_3606)
);

AOI22xp5_ASAP7_75t_L g3607 ( 
.A1(n_3525),
.A2(n_500),
.B1(n_498),
.B2(n_499),
.Y(n_3607)
);

AOI22xp5_ASAP7_75t_L g3608 ( 
.A1(n_3538),
.A2(n_502),
.B1(n_500),
.B2(n_501),
.Y(n_3608)
);

INVx1_ASAP7_75t_L g3609 ( 
.A(n_3535),
.Y(n_3609)
);

INVx1_ASAP7_75t_L g3610 ( 
.A(n_3548),
.Y(n_3610)
);

XOR2x2_ASAP7_75t_L g3611 ( 
.A(n_3540),
.B(n_501),
.Y(n_3611)
);

O2A1O1Ixp33_ASAP7_75t_L g3612 ( 
.A1(n_3594),
.A2(n_505),
.B(n_502),
.C(n_504),
.Y(n_3612)
);

O2A1O1Ixp33_ASAP7_75t_L g3613 ( 
.A1(n_3560),
.A2(n_507),
.B(n_504),
.C(n_506),
.Y(n_3613)
);

AOI211xp5_ASAP7_75t_SL g3614 ( 
.A1(n_3568),
.A2(n_509),
.B(n_507),
.C(n_508),
.Y(n_3614)
);

NAND4xp25_ASAP7_75t_L g3615 ( 
.A(n_3572),
.B(n_510),
.C(n_508),
.D(n_509),
.Y(n_3615)
);

OAI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3529),
.A2(n_512),
.B1(n_510),
.B2(n_511),
.Y(n_3616)
);

AOI211xp5_ASAP7_75t_L g3617 ( 
.A1(n_3533),
.A2(n_513),
.B(n_511),
.C(n_512),
.Y(n_3617)
);

NAND3xp33_ASAP7_75t_L g3618 ( 
.A(n_3532),
.B(n_513),
.C(n_514),
.Y(n_3618)
);

AOI221xp5_ASAP7_75t_L g3619 ( 
.A1(n_3580),
.A2(n_517),
.B1(n_514),
.B2(n_516),
.C(n_519),
.Y(n_3619)
);

AOI211xp5_ASAP7_75t_L g3620 ( 
.A1(n_3578),
.A2(n_522),
.B(n_520),
.C(n_521),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3573),
.B(n_520),
.Y(n_3621)
);

BUFx2_ASAP7_75t_L g3622 ( 
.A(n_3563),
.Y(n_3622)
);

O2A1O1Ixp33_ASAP7_75t_L g3623 ( 
.A1(n_3554),
.A2(n_523),
.B(n_521),
.C(n_522),
.Y(n_3623)
);

AOI211xp5_ASAP7_75t_L g3624 ( 
.A1(n_3559),
.A2(n_526),
.B(n_524),
.C(n_525),
.Y(n_3624)
);

AOI211xp5_ASAP7_75t_SL g3625 ( 
.A1(n_3561),
.A2(n_527),
.B(n_525),
.C(n_526),
.Y(n_3625)
);

OAI211xp5_ASAP7_75t_SL g3626 ( 
.A1(n_3545),
.A2(n_531),
.B(n_527),
.C(n_530),
.Y(n_3626)
);

NOR2x1_ASAP7_75t_L g3627 ( 
.A(n_3553),
.B(n_533),
.Y(n_3627)
);

NAND3x1_ASAP7_75t_L g3628 ( 
.A(n_3556),
.B(n_534),
.C(n_535),
.Y(n_3628)
);

OAI211xp5_ASAP7_75t_L g3629 ( 
.A1(n_3581),
.A2(n_537),
.B(n_534),
.C(n_535),
.Y(n_3629)
);

OAI211xp5_ASAP7_75t_SL g3630 ( 
.A1(n_3558),
.A2(n_539),
.B(n_537),
.C(n_538),
.Y(n_3630)
);

OAI221xp5_ASAP7_75t_L g3631 ( 
.A1(n_3541),
.A2(n_541),
.B1(n_539),
.B2(n_540),
.C(n_542),
.Y(n_3631)
);

NOR3xp33_ASAP7_75t_L g3632 ( 
.A(n_3585),
.B(n_541),
.C(n_542),
.Y(n_3632)
);

AOI22xp33_ASAP7_75t_SL g3633 ( 
.A1(n_3544),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_3633)
);

OAI221xp5_ASAP7_75t_L g3634 ( 
.A1(n_3542),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.C(n_546),
.Y(n_3634)
);

NAND4xp25_ASAP7_75t_L g3635 ( 
.A(n_3536),
.B(n_548),
.C(n_546),
.D(n_547),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3579),
.B(n_547),
.Y(n_3636)
);

INVx5_ASAP7_75t_L g3637 ( 
.A(n_3586),
.Y(n_3637)
);

OAI211xp5_ASAP7_75t_L g3638 ( 
.A1(n_3562),
.A2(n_550),
.B(n_548),
.C(n_549),
.Y(n_3638)
);

OAI221xp5_ASAP7_75t_SL g3639 ( 
.A1(n_3575),
.A2(n_551),
.B1(n_549),
.B2(n_550),
.C(n_552),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3570),
.B(n_551),
.Y(n_3640)
);

OAI21xp5_ASAP7_75t_L g3641 ( 
.A1(n_3577),
.A2(n_552),
.B(n_553),
.Y(n_3641)
);

OAI211xp5_ASAP7_75t_SL g3642 ( 
.A1(n_3584),
.A2(n_556),
.B(n_554),
.C(n_555),
.Y(n_3642)
);

AOI221xp5_ASAP7_75t_L g3643 ( 
.A1(n_3590),
.A2(n_556),
.B1(n_554),
.B2(n_555),
.C(n_557),
.Y(n_3643)
);

AOI221xp5_ASAP7_75t_L g3644 ( 
.A1(n_3550),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.C(n_560),
.Y(n_3644)
);

AOI221xp5_ASAP7_75t_L g3645 ( 
.A1(n_3588),
.A2(n_560),
.B1(n_558),
.B2(n_559),
.C(n_561),
.Y(n_3645)
);

NAND3xp33_ASAP7_75t_L g3646 ( 
.A(n_3583),
.B(n_561),
.C(n_562),
.Y(n_3646)
);

AOI221xp5_ASAP7_75t_L g3647 ( 
.A1(n_3546),
.A2(n_564),
.B1(n_562),
.B2(n_563),
.C(n_565),
.Y(n_3647)
);

AOI211xp5_ASAP7_75t_SL g3648 ( 
.A1(n_3589),
.A2(n_566),
.B(n_563),
.C(n_565),
.Y(n_3648)
);

NAND3xp33_ASAP7_75t_L g3649 ( 
.A(n_3587),
.B(n_566),
.C(n_567),
.Y(n_3649)
);

OAI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3566),
.A2(n_567),
.B(n_568),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3564),
.Y(n_3651)
);

AOI221xp5_ASAP7_75t_L g3652 ( 
.A1(n_3547),
.A2(n_570),
.B1(n_568),
.B2(n_569),
.C(n_571),
.Y(n_3652)
);

AOI211xp5_ASAP7_75t_L g3653 ( 
.A1(n_3595),
.A2(n_572),
.B(n_569),
.C(n_571),
.Y(n_3653)
);

NAND2xp33_ASAP7_75t_L g3654 ( 
.A(n_3628),
.B(n_3549),
.Y(n_3654)
);

INVx1_ASAP7_75t_L g3655 ( 
.A(n_3622),
.Y(n_3655)
);

XNOR2xp5_ASAP7_75t_L g3656 ( 
.A(n_3611),
.B(n_3565),
.Y(n_3656)
);

INVx1_ASAP7_75t_L g3657 ( 
.A(n_3609),
.Y(n_3657)
);

AND2x2_ASAP7_75t_SL g3658 ( 
.A(n_3604),
.B(n_3571),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3606),
.A2(n_3576),
.B1(n_3557),
.B2(n_3569),
.Y(n_3659)
);

NAND4xp75_ASAP7_75t_L g3660 ( 
.A(n_3597),
.B(n_3569),
.C(n_3582),
.D(n_3592),
.Y(n_3660)
);

INVx2_ASAP7_75t_SL g3661 ( 
.A(n_3637),
.Y(n_3661)
);

NOR2xp67_ASAP7_75t_L g3662 ( 
.A(n_3637),
.B(n_3552),
.Y(n_3662)
);

AOI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_3599),
.A2(n_3593),
.B1(n_575),
.B2(n_573),
.Y(n_3663)
);

NOR2x1_ASAP7_75t_L g3664 ( 
.A(n_3618),
.B(n_3635),
.Y(n_3664)
);

AND2x2_ASAP7_75t_L g3665 ( 
.A(n_3637),
.B(n_573),
.Y(n_3665)
);

NOR2x1_ASAP7_75t_L g3666 ( 
.A(n_3629),
.B(n_574),
.Y(n_3666)
);

NAND4xp75_ASAP7_75t_L g3667 ( 
.A(n_3603),
.B(n_576),
.C(n_574),
.D(n_575),
.Y(n_3667)
);

AOI22xp5_ASAP7_75t_L g3668 ( 
.A1(n_3626),
.A2(n_580),
.B1(n_577),
.B2(n_579),
.Y(n_3668)
);

NAND4xp75_ASAP7_75t_L g3669 ( 
.A(n_3627),
.B(n_582),
.C(n_579),
.D(n_581),
.Y(n_3669)
);

INVxp33_ASAP7_75t_SL g3670 ( 
.A(n_3607),
.Y(n_3670)
);

AND3x4_ASAP7_75t_L g3671 ( 
.A(n_3632),
.B(n_581),
.C(n_582),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3625),
.B(n_3614),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_L g3673 ( 
.A(n_3605),
.B(n_583),
.Y(n_3673)
);

XNOR2xp5_ASAP7_75t_L g3674 ( 
.A(n_3624),
.B(n_583),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3621),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3651),
.Y(n_3676)
);

NAND2xp5_ASAP7_75t_L g3677 ( 
.A(n_3620),
.B(n_584),
.Y(n_3677)
);

NOR2x1_ASAP7_75t_L g3678 ( 
.A(n_3615),
.B(n_584),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3636),
.Y(n_3679)
);

NOR2x1_ASAP7_75t_L g3680 ( 
.A(n_3646),
.B(n_585),
.Y(n_3680)
);

INVx1_ASAP7_75t_L g3681 ( 
.A(n_3610),
.Y(n_3681)
);

NOR2x1_ASAP7_75t_L g3682 ( 
.A(n_3649),
.B(n_586),
.Y(n_3682)
);

NOR2x1_ASAP7_75t_L g3683 ( 
.A(n_3612),
.B(n_586),
.Y(n_3683)
);

NOR2x1_ASAP7_75t_L g3684 ( 
.A(n_3616),
.B(n_587),
.Y(n_3684)
);

NOR2xp33_ASAP7_75t_L g3685 ( 
.A(n_3640),
.B(n_588),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3661),
.B(n_3648),
.Y(n_3686)
);

NAND2xp5_ASAP7_75t_L g3687 ( 
.A(n_3665),
.B(n_3619),
.Y(n_3687)
);

NOR2xp33_ASAP7_75t_R g3688 ( 
.A(n_3654),
.B(n_3633),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_3658),
.B(n_3662),
.Y(n_3689)
);

XNOR2xp5_ASAP7_75t_L g3690 ( 
.A(n_3656),
.B(n_3653),
.Y(n_3690)
);

NAND2xp33_ASAP7_75t_SL g3691 ( 
.A(n_3672),
.B(n_3641),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_SL g3692 ( 
.A(n_3659),
.B(n_3602),
.Y(n_3692)
);

NAND2xp33_ASAP7_75t_SL g3693 ( 
.A(n_3671),
.B(n_3655),
.Y(n_3693)
);

NOR2xp33_ASAP7_75t_R g3694 ( 
.A(n_3673),
.B(n_3617),
.Y(n_3694)
);

NOR3xp33_ASAP7_75t_SL g3695 ( 
.A(n_3660),
.B(n_3596),
.C(n_3631),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_SL g3696 ( 
.A(n_3666),
.B(n_3643),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_SL g3697 ( 
.A(n_3668),
.B(n_3600),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3683),
.B(n_3647),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_SL g3699 ( 
.A(n_3663),
.B(n_3684),
.Y(n_3699)
);

NAND3xp33_ASAP7_75t_L g3700 ( 
.A(n_3682),
.B(n_3598),
.C(n_3601),
.Y(n_3700)
);

NOR2xp33_ASAP7_75t_R g3701 ( 
.A(n_3674),
.B(n_3657),
.Y(n_3701)
);

BUFx2_ASAP7_75t_L g3702 ( 
.A(n_3688),
.Y(n_3702)
);

BUFx2_ASAP7_75t_L g3703 ( 
.A(n_3689),
.Y(n_3703)
);

CKINVDCx16_ASAP7_75t_R g3704 ( 
.A(n_3694),
.Y(n_3704)
);

AOI31xp33_ASAP7_75t_L g3705 ( 
.A1(n_3690),
.A2(n_3680),
.A3(n_3678),
.B(n_3675),
.Y(n_3705)
);

BUFx2_ASAP7_75t_L g3706 ( 
.A(n_3693),
.Y(n_3706)
);

AOI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_3692),
.A2(n_3670),
.B(n_3677),
.Y(n_3707)
);

INVx1_ASAP7_75t_L g3708 ( 
.A(n_3706),
.Y(n_3708)
);

AOI22xp5_ASAP7_75t_L g3709 ( 
.A1(n_3704),
.A2(n_3691),
.B1(n_3696),
.B2(n_3664),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3703),
.Y(n_3710)
);

OAI22x1_ASAP7_75t_SL g3711 ( 
.A1(n_3708),
.A2(n_3679),
.B1(n_3681),
.B2(n_3676),
.Y(n_3711)
);

XOR2xp5_ASAP7_75t_L g3712 ( 
.A(n_3709),
.B(n_3669),
.Y(n_3712)
);

OAI22xp5_ASAP7_75t_L g3713 ( 
.A1(n_3710),
.A2(n_3700),
.B1(n_3695),
.B2(n_3608),
.Y(n_3713)
);

AOI31xp33_ASAP7_75t_L g3714 ( 
.A1(n_3713),
.A2(n_3686),
.A3(n_3707),
.B(n_3687),
.Y(n_3714)
);

AOI31xp33_ASAP7_75t_L g3715 ( 
.A1(n_3712),
.A2(n_3698),
.A3(n_3699),
.B(n_3697),
.Y(n_3715)
);

AOI31xp33_ASAP7_75t_L g3716 ( 
.A1(n_3711),
.A2(n_3685),
.A3(n_3650),
.B(n_3645),
.Y(n_3716)
);

AOI22xp33_ASAP7_75t_L g3717 ( 
.A1(n_3715),
.A2(n_3702),
.B1(n_3701),
.B2(n_3642),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3716),
.B(n_3705),
.Y(n_3718)
);

OR2x2_ASAP7_75t_L g3719 ( 
.A(n_3714),
.B(n_3667),
.Y(n_3719)
);

AOI222xp33_ASAP7_75t_L g3720 ( 
.A1(n_3718),
.A2(n_3652),
.B1(n_3644),
.B2(n_3634),
.C1(n_3638),
.C2(n_3630),
.Y(n_3720)
);

OAI22xp5_ASAP7_75t_L g3721 ( 
.A1(n_3717),
.A2(n_3639),
.B1(n_3623),
.B2(n_3613),
.Y(n_3721)
);

AO21x2_ASAP7_75t_L g3722 ( 
.A1(n_3719),
.A2(n_588),
.B(n_589),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3722),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3721),
.Y(n_3724)
);

OAI221xp5_ASAP7_75t_R g3725 ( 
.A1(n_3724),
.A2(n_3720),
.B1(n_591),
.B2(n_589),
.C(n_590),
.Y(n_3725)
);

OAI221xp5_ASAP7_75t_R g3726 ( 
.A1(n_3723),
.A2(n_592),
.B1(n_590),
.B2(n_591),
.C(n_593),
.Y(n_3726)
);

AOI211xp5_ASAP7_75t_L g3727 ( 
.A1(n_3726),
.A2(n_3725),
.B(n_596),
.C(n_595),
.Y(n_3727)
);


endmodule