module fake_netlist_1_11088_n_914 (n_117, n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_16, n_13, n_113, n_95, n_120, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_122, n_118, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_914);
input n_117;
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_16;
input n_13;
input n_113;
input n_95;
input n_120;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_122;
input n_118;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_914;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_878;
wire n_814;
wire n_911;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_227;
wire n_384;
wire n_617;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_909;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_638;
wire n_540;
wire n_830;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_769;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_844;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_703;
wire n_331;
wire n_485;
wire n_813;
wire n_442;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_699;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_822;
wire n_706;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_200;
wire n_208;
wire n_573;
wire n_898;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_240;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_493;
wire n_698;
wire n_555;
wire n_418;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_650;
wire n_625;
wire n_521;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g124 ( .A(n_76), .Y(n_124) );
BUFx2_ASAP7_75t_L g125 ( .A(n_59), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_14), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_112), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_40), .Y(n_128) );
HB1xp67_ASAP7_75t_L g129 ( .A(n_3), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_91), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_5), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_120), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_56), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_113), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_39), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_103), .Y(n_136) );
INVxp33_ASAP7_75t_SL g137 ( .A(n_83), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_105), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_45), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_11), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_90), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_115), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_108), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_49), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_123), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_75), .Y(n_146) );
BUFx2_ASAP7_75t_SL g147 ( .A(n_19), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_15), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_29), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_111), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_7), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_69), .Y(n_152) );
INVx2_ASAP7_75t_SL g153 ( .A(n_72), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_63), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_46), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_55), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_77), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_2), .Y(n_158) );
INVxp67_ASAP7_75t_L g159 ( .A(n_35), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_19), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_96), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_100), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_88), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_28), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_14), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_84), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_98), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_102), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_5), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_58), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_30), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_20), .Y(n_172) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_57), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_74), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_27), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_129), .B(n_0), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_124), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_153), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_153), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
INVx5_ASAP7_75t_L g182 ( .A(n_125), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_173), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_139), .B(n_1), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_126), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_136), .B(n_3), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_139), .B(n_4), .Y(n_187) );
OAI21x1_ASAP7_75t_L g188 ( .A1(n_145), .A2(n_60), .B(n_121), .Y(n_188) );
INVx5_ASAP7_75t_L g189 ( .A(n_148), .Y(n_189) );
AND2x6_ASAP7_75t_L g190 ( .A(n_150), .B(n_24), .Y(n_190) );
NOR2x1_ASAP7_75t_L g191 ( .A(n_140), .B(n_25), .Y(n_191) );
OAI22x1_ASAP7_75t_SL g192 ( .A1(n_126), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_148), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_151), .B(n_6), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_160), .B(n_8), .Y(n_195) );
INVxp33_ASAP7_75t_SL g196 ( .A(n_131), .Y(n_196) );
AOI22xp5_ASAP7_75t_SL g197 ( .A1(n_147), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_131), .B(n_9), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_148), .Y(n_199) );
INVx3_ASAP7_75t_L g200 ( .A(n_187), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_187), .Y(n_201) );
INVx2_ASAP7_75t_SL g202 ( .A(n_182), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_189), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_187), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_182), .B(n_128), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_189), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_189), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_189), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
AND2x6_ASAP7_75t_L g211 ( .A(n_195), .B(n_155), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_193), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_193), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_195), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_182), .B(n_159), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_195), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_193), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_195), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_193), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_194), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_194), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_193), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_193), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_194), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_199), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_199), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_199), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_199), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_199), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_177), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_196), .A2(n_169), .B1(n_172), .B2(n_170), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
INVxp67_ASAP7_75t_SL g233 ( .A(n_185), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_179), .B(n_148), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_180), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_182), .B(n_169), .Y(n_236) );
INVx1_ASAP7_75t_SL g237 ( .A(n_185), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_177), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_178), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_230), .B(n_182), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_211), .Y(n_241) );
NAND2xp33_ASAP7_75t_SL g242 ( .A(n_214), .B(n_127), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_211), .Y(n_243) );
HB1xp67_ASAP7_75t_L g244 ( .A(n_237), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_237), .B(n_196), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_218), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_211), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_218), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_239), .B(n_182), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_233), .B(n_176), .Y(n_250) );
NOR3xp33_ASAP7_75t_L g251 ( .A(n_231), .B(n_198), .C(n_183), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_220), .B(n_128), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_230), .B(n_178), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_220), .B(n_164), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g256 ( .A(n_231), .B(n_181), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_224), .B(n_164), .Y(n_257) );
NOR2xp67_ASAP7_75t_SL g258 ( .A(n_214), .B(n_174), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_238), .B(n_181), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_238), .B(n_180), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_239), .B(n_186), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_211), .A2(n_172), .B1(n_167), .B2(n_138), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_201), .A2(n_192), .B1(n_158), .B2(n_165), .C(n_184), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_224), .B(n_174), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_216), .B(n_137), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_211), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_216), .A2(n_188), .B(n_197), .C(n_191), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_211), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_218), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_221), .B(n_137), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_234), .Y(n_271) );
INVx8_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_234), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_221), .B(n_133), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_234), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_221), .B(n_134), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_200), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_232), .B(n_190), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_221), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_232), .B(n_190), .Y(n_281) );
INVxp67_ASAP7_75t_L g282 ( .A(n_236), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_235), .B(n_190), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_235), .B(n_190), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_201), .B(n_190), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_204), .B(n_190), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_204), .B(n_148), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_200), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g289 ( .A(n_200), .B(n_135), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_200), .B(n_141), .Y(n_290) );
INVxp67_ASAP7_75t_SL g291 ( .A(n_202), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_202), .B(n_190), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_215), .A2(n_192), .B1(n_161), .B2(n_166), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_206), .A2(n_171), .B1(n_142), .B2(n_168), .Y(n_294) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_203), .A2(n_143), .B1(n_144), .B2(n_146), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_203), .B(n_149), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_285), .A2(n_188), .B(n_209), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_245), .B(n_152), .Y(n_298) );
AOI22xp33_ASAP7_75t_SL g299 ( .A1(n_244), .A2(n_154), .B1(n_156), .B2(n_157), .Y(n_299) );
INVx11_ASAP7_75t_L g300 ( .A(n_242), .Y(n_300) );
CKINVDCx8_ASAP7_75t_R g301 ( .A(n_272), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_L g302 ( .A1(n_267), .A2(n_217), .B(n_207), .C(n_208), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_286), .A2(n_213), .B(n_205), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_250), .B(n_162), .Y(n_305) );
AOI21xp33_ASAP7_75t_L g306 ( .A1(n_258), .A2(n_163), .B(n_175), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_267), .A2(n_217), .B(n_207), .C(n_208), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_251), .B(n_10), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_256), .B(n_205), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_279), .A2(n_222), .B(n_210), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_242), .A2(n_222), .B1(n_210), .B2(n_212), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_281), .A2(n_223), .B(n_212), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_262), .A2(n_223), .B1(n_213), .B2(n_219), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_246), .Y(n_314) );
CKINVDCx8_ASAP7_75t_R g315 ( .A(n_272), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_247), .B(n_11), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_278), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g318 ( .A(n_241), .B(n_209), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_283), .A2(n_219), .B(n_225), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_246), .Y(n_320) );
INVx3_ASAP7_75t_L g321 ( .A(n_271), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_284), .A2(n_225), .B(n_227), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_292), .A2(n_248), .B(n_254), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_241), .B(n_228), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_248), .A2(n_229), .B(n_227), .Y(n_325) );
NOR2x1_ASAP7_75t_L g326 ( .A(n_270), .B(n_226), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_282), .B(n_12), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_254), .A2(n_229), .B(n_226), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_278), .A2(n_228), .B(n_13), .C(n_15), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_253), .B(n_12), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_241), .B(n_228), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_259), .B(n_13), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_269), .A2(n_228), .B(n_68), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_274), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_276), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_269), .A2(n_228), .B(n_67), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_261), .B(n_16), .Y(n_337) );
INVxp67_ASAP7_75t_L g338 ( .A(n_258), .Y(n_338) );
NOR3xp33_ASAP7_75t_L g339 ( .A(n_263), .B(n_16), .C(n_17), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_280), .A2(n_70), .B(n_119), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_247), .B(n_17), .Y(n_341) );
AO21x1_ASAP7_75t_L g342 ( .A1(n_240), .A2(n_18), .B(n_20), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_265), .B(n_18), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_280), .A2(n_122), .B(n_71), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_260), .A2(n_118), .B(n_66), .Y(n_345) );
OAI222xp33_ASAP7_75t_L g346 ( .A1(n_308), .A2(n_293), .B1(n_266), .B2(n_287), .C1(n_257), .C2(n_252), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_323), .A2(n_288), .B(n_272), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_301), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_322), .A2(n_288), .B(n_272), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_302), .A2(n_249), .B(n_268), .Y(n_350) );
INVx5_ASAP7_75t_L g351 ( .A(n_316), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_303), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_322), .A2(n_290), .B(n_289), .Y(n_353) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_316), .A2(n_266), .B1(n_243), .B2(n_241), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_305), .B(n_255), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_315), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_307), .A2(n_337), .B(n_330), .C(n_332), .Y(n_357) );
O2A1O1Ixp5_ASAP7_75t_L g358 ( .A1(n_297), .A2(n_275), .B(n_277), .C(n_287), .Y(n_358) );
OAI22x1_ASAP7_75t_L g359 ( .A1(n_341), .A2(n_264), .B1(n_273), .B2(n_271), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_297), .A2(n_273), .B(n_296), .Y(n_360) );
INVx3_ASAP7_75t_L g361 ( .A(n_321), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_343), .B(n_243), .Y(n_362) );
AOI21x1_ASAP7_75t_L g363 ( .A1(n_345), .A2(n_294), .B(n_268), .Y(n_363) );
AO21x1_ASAP7_75t_L g364 ( .A1(n_345), .A2(n_344), .B(n_340), .Y(n_364) );
BUFx3_ASAP7_75t_L g365 ( .A(n_341), .Y(n_365) );
O2A1O1Ixp5_ASAP7_75t_L g366 ( .A1(n_324), .A2(n_291), .B(n_295), .C(n_243), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_327), .A2(n_241), .B1(n_243), .B2(n_23), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_312), .A2(n_243), .B(n_73), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_311), .B(n_21), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_338), .A2(n_21), .B1(n_22), .B2(n_23), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_339), .B(n_22), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_298), .A2(n_26), .B(n_31), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g373 ( .A1(n_329), .A2(n_32), .B(n_33), .C(n_34), .Y(n_373) );
AO21x2_ASAP7_75t_L g374 ( .A1(n_340), .A2(n_36), .B(n_37), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_300), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_299), .B(n_38), .Y(n_376) );
AO21x1_ASAP7_75t_L g377 ( .A1(n_344), .A2(n_41), .B(n_42), .Y(n_377) );
AOI21x1_ASAP7_75t_L g378 ( .A1(n_333), .A2(n_43), .B(n_44), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_334), .B(n_47), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_335), .B(n_48), .Y(n_380) );
AO31x2_ASAP7_75t_L g381 ( .A1(n_357), .A2(n_342), .A3(n_336), .B(n_312), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_357), .A2(n_310), .B(n_304), .Y(n_382) );
OAI21x1_ASAP7_75t_L g383 ( .A1(n_364), .A2(n_360), .B(n_363), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_352), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
BUFx2_ASAP7_75t_R g386 ( .A(n_348), .Y(n_386) );
OAI21x1_ASAP7_75t_L g387 ( .A1(n_360), .A2(n_358), .B(n_368), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_365), .A2(n_317), .B1(n_309), .B2(n_321), .Y(n_388) );
INVx2_ASAP7_75t_SL g389 ( .A(n_351), .Y(n_389) );
AO21x1_ASAP7_75t_L g390 ( .A1(n_349), .A2(n_313), .B(n_319), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_331), .B(n_318), .Y(n_391) );
OAI21x1_ASAP7_75t_SL g392 ( .A1(n_377), .A2(n_320), .B(n_314), .Y(n_392) );
BUFx2_ASAP7_75t_R g393 ( .A(n_348), .Y(n_393) );
INVx1_ASAP7_75t_SL g394 ( .A(n_365), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_351), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
OAI21x1_ASAP7_75t_L g397 ( .A1(n_378), .A2(n_325), .B(n_328), .Y(n_397) );
INVx3_ASAP7_75t_L g398 ( .A(n_351), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g399 ( .A(n_373), .B(n_306), .C(n_326), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_356), .B(n_50), .Y(n_400) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_375), .B(n_356), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
OAI21x1_ASAP7_75t_L g403 ( .A1(n_347), .A2(n_51), .B(n_52), .Y(n_403) );
OAI21x1_ASAP7_75t_L g404 ( .A1(n_366), .A2(n_53), .B(n_54), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_354), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_355), .B(n_61), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_356), .Y(n_407) );
OA21x2_ASAP7_75t_L g408 ( .A1(n_350), .A2(n_62), .B(n_64), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_383), .A2(n_353), .B(n_367), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_405), .A2(n_371), .B1(n_370), .B2(n_369), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_402), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_402), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_388), .B(n_361), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_385), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_395), .Y(n_417) );
AOI21x1_ASAP7_75t_L g418 ( .A1(n_392), .A2(n_359), .B(n_379), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_390), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_385), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_405), .A2(n_359), .B1(n_376), .B2(n_361), .Y(n_421) );
BUFx3_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
BUFx3_ASAP7_75t_L g423 ( .A(n_395), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_387), .Y(n_424) );
CKINVDCx8_ASAP7_75t_R g425 ( .A(n_400), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_387), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_384), .A2(n_374), .B1(n_372), .B2(n_375), .Y(n_427) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_375), .B1(n_380), .B2(n_362), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_390), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_396), .Y(n_431) );
OAI21x1_ASAP7_75t_L g432 ( .A1(n_392), .A2(n_374), .B(n_346), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_381), .Y(n_433) );
OA21x2_ASAP7_75t_L g434 ( .A1(n_404), .A2(n_65), .B(n_78), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_381), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_382), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_382), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_396), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_382), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_381), .Y(n_441) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_382), .A2(n_79), .B(n_80), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_425), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_433), .B(n_381), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_411), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_411), .B(n_406), .Y(n_447) );
INVx3_ASAP7_75t_L g448 ( .A(n_425), .Y(n_448) );
BUFx2_ASAP7_75t_SL g449 ( .A(n_425), .Y(n_449) );
AO31x2_ASAP7_75t_L g450 ( .A1(n_419), .A2(n_381), .A3(n_399), .B(n_408), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_423), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_413), .Y(n_452) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_435), .Y(n_453) );
INVx3_ASAP7_75t_L g454 ( .A(n_431), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
AOI21xp5_ASAP7_75t_SL g456 ( .A1(n_423), .A2(n_400), .B(n_408), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_410), .A2(n_407), .B1(n_400), .B2(n_406), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_433), .B(n_381), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_436), .B(n_408), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_410), .A2(n_407), .B1(n_400), .B2(n_394), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_423), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_436), .B(n_396), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_437), .Y(n_463) );
BUFx12f_ASAP7_75t_L g464 ( .A(n_420), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_441), .B(n_408), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_441), .B(n_391), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_437), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_419), .B(n_391), .Y(n_468) );
AOI22xp33_ASAP7_75t_SL g469 ( .A1(n_417), .A2(n_407), .B1(n_396), .B2(n_398), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_428), .A2(n_399), .B1(n_401), .B2(n_389), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_414), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_429), .B(n_437), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_437), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_429), .B(n_391), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_414), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_438), .B(n_391), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_435), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_414), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_438), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_417), .Y(n_480) );
INVx5_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
INVx3_ASAP7_75t_L g482 ( .A(n_431), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_417), .B(n_398), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_423), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_422), .Y(n_485) );
INVx3_ASAP7_75t_L g486 ( .A(n_431), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_438), .B(n_440), .Y(n_487) );
INVxp67_ASAP7_75t_SL g488 ( .A(n_412), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_438), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_420), .B(n_398), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_440), .B(n_412), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g492 ( .A(n_416), .B(n_398), .Y(n_492) );
INVx3_ASAP7_75t_L g493 ( .A(n_431), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_440), .B(n_389), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_440), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_422), .Y(n_496) );
NAND2xp33_ASAP7_75t_L g497 ( .A(n_420), .B(n_393), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_412), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_412), .B(n_403), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_458), .B(n_424), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_458), .B(n_424), .Y(n_501) );
INVx4_ASAP7_75t_L g502 ( .A(n_464), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_463), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_446), .B(n_422), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_452), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_463), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_452), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_481), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_481), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_457), .A2(n_428), .B1(n_421), .B2(n_422), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_458), .B(n_424), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_466), .B(n_426), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_466), .B(n_426), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_466), .B(n_426), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_455), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_481), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_455), .B(n_416), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_472), .B(n_426), .Y(n_520) );
AND2x4_ASAP7_75t_SL g521 ( .A(n_448), .B(n_416), .Y(n_521) );
INVx3_ASAP7_75t_L g522 ( .A(n_481), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_471), .Y(n_523) );
BUFx3_ASAP7_75t_L g524 ( .A(n_464), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_467), .Y(n_525) );
BUFx12f_ASAP7_75t_L g526 ( .A(n_464), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_472), .B(n_430), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_471), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_475), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_477), .B(n_415), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_475), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_497), .B(n_393), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_472), .B(n_430), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_487), .B(n_430), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_451), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_477), .B(n_415), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_467), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_478), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_467), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_473), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_457), .A2(n_421), .B1(n_416), .B2(n_439), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_478), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_460), .A2(n_439), .B1(n_427), .B2(n_443), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_460), .A2(n_439), .B1(n_427), .B2(n_443), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_489), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_483), .B(n_386), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
INVx4_ASAP7_75t_L g549 ( .A(n_481), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_496), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_487), .B(n_430), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_489), .Y(n_552) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_444), .B(n_439), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_480), .B(n_439), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_487), .B(n_443), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_468), .B(n_443), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_451), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_480), .B(n_443), .Y(n_558) );
NAND2x1p5_ASAP7_75t_SL g559 ( .A(n_461), .B(n_468), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_473), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_453), .B(n_409), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_484), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_468), .B(n_432), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_474), .B(n_432), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_479), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_479), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_453), .B(n_409), .Y(n_567) );
INVx3_ASAP7_75t_L g568 ( .A(n_481), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
INVx2_ASAP7_75t_L g570 ( .A(n_495), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_495), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_481), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_474), .B(n_491), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_447), .B(n_401), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_495), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_498), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_498), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_491), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_447), .B(n_432), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_491), .Y(n_580) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_496), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_462), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_573), .B(n_484), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_582), .B(n_462), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_505), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_505), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_573), .B(n_484), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_500), .B(n_461), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_506), .Y(n_589) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_560), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_503), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_582), .B(n_578), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_506), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_500), .B(n_461), .Y(n_595) );
INVx2_ASAP7_75t_L g596 ( .A(n_507), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_578), .B(n_494), .Y(n_597) );
AND2x4_ASAP7_75t_L g598 ( .A(n_549), .B(n_485), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_549), .B(n_485), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_580), .B(n_474), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_501), .B(n_485), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_501), .B(n_482), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_549), .B(n_481), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_508), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_508), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_580), .B(n_512), .Y(n_606) );
AND2x4_ASAP7_75t_L g607 ( .A(n_510), .B(n_518), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_512), .B(n_476), .Y(n_608) );
AND2x4_ASAP7_75t_L g609 ( .A(n_510), .B(n_482), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_513), .B(n_476), .Y(n_610) );
OR2x2_ASAP7_75t_L g611 ( .A(n_530), .B(n_494), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_513), .B(n_476), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_517), .Y(n_613) );
NOR2x1p5_ASAP7_75t_L g614 ( .A(n_526), .B(n_448), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_514), .B(n_445), .Y(n_615) );
INVx3_ASAP7_75t_L g616 ( .A(n_510), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_560), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_517), .B(n_445), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_562), .B(n_486), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_535), .B(n_486), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_566), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_523), .Y(n_622) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_566), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_530), .B(n_445), .Y(n_624) );
BUFx3_ASAP7_75t_L g625 ( .A(n_526), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_502), .A2(n_469), .B1(n_449), .B2(n_448), .Y(n_626) );
NAND2x1_ASAP7_75t_SL g627 ( .A(n_502), .B(n_448), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_571), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_536), .B(n_483), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_535), .B(n_486), .Y(n_630) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_502), .B(n_456), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_523), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_528), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_536), .B(n_483), .Y(n_634) );
NAND4xp75_ASAP7_75t_L g635 ( .A(n_532), .B(n_490), .C(n_465), .D(n_459), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_514), .B(n_459), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_528), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_516), .B(n_459), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_516), .B(n_465), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_529), .Y(n_640) );
INVx4_ASAP7_75t_L g641 ( .A(n_524), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_529), .Y(n_642) );
AND2x2_ASAP7_75t_L g643 ( .A(n_542), .B(n_486), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_559), .B(n_494), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_531), .B(n_469), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_524), .B(n_444), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_507), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_531), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_538), .B(n_470), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_538), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_542), .B(n_482), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_557), .B(n_482), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_515), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_563), .B(n_465), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_543), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_515), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_543), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_525), .Y(n_658) );
AND2x4_ASAP7_75t_L g659 ( .A(n_518), .B(n_454), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_544), .B(n_470), .C(n_493), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_557), .B(n_493), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_534), .B(n_493), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_546), .Y(n_663) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_571), .Y(n_664) );
INVx2_ASAP7_75t_L g665 ( .A(n_525), .Y(n_665) );
OR2x2_ASAP7_75t_L g666 ( .A(n_559), .B(n_493), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_546), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_552), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_552), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_537), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_563), .B(n_499), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_559), .B(n_454), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_519), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_534), .B(n_454), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_518), .B(n_454), .Y(n_675) );
NAND2x1_ASAP7_75t_L g676 ( .A(n_522), .B(n_444), .Y(n_676) );
INVxp67_ASAP7_75t_L g677 ( .A(n_581), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_504), .B(n_488), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_551), .B(n_444), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_537), .Y(n_680) );
NAND4xp75_ASAP7_75t_L g681 ( .A(n_645), .B(n_547), .C(n_509), .D(n_556), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_583), .B(n_550), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_587), .B(n_551), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_608), .B(n_522), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_608), .B(n_522), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_592), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_603), .B(n_568), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_585), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_615), .B(n_568), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_615), .B(n_568), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_606), .B(n_554), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_611), .B(n_554), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_586), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_673), .B(n_577), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_601), .B(n_572), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_654), .B(n_572), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_654), .B(n_572), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_600), .B(n_577), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_589), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_610), .B(n_527), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_593), .Y(n_701) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_590), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_590), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_604), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_605), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_613), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_663), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_667), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_668), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_625), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_669), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_622), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_632), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_633), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_610), .B(n_527), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_637), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_624), .B(n_576), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_640), .Y(n_718) );
AND2x4_ASAP7_75t_SL g719 ( .A(n_641), .B(n_444), .Y(n_719) );
OR2x2_ASAP7_75t_L g720 ( .A(n_629), .B(n_520), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_612), .B(n_520), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_617), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_603), .B(n_509), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_642), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_612), .B(n_564), .Y(n_725) );
NOR2xp67_ASAP7_75t_R g726 ( .A(n_641), .B(n_449), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_648), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_650), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_655), .Y(n_729) );
OR2x6_ASAP7_75t_L g730 ( .A(n_631), .B(n_553), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_657), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_636), .B(n_576), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_634), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_671), .B(n_533), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_617), .Y(n_735) );
NAND2x1p5_ASAP7_75t_L g736 ( .A(n_641), .B(n_565), .Y(n_736) );
AND2x2_ASAP7_75t_L g737 ( .A(n_602), .B(n_564), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_621), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_621), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_636), .B(n_556), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_623), .Y(n_741) );
AND2x4_ASAP7_75t_L g742 ( .A(n_603), .B(n_533), .Y(n_742) );
INVx2_ASAP7_75t_L g743 ( .A(n_591), .Y(n_743) );
AND2x4_ASAP7_75t_L g744 ( .A(n_607), .B(n_533), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_638), .B(n_555), .Y(n_745) );
OR2x2_ASAP7_75t_L g746 ( .A(n_671), .B(n_533), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_588), .B(n_555), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_623), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_626), .A2(n_511), .B1(n_545), .B2(n_574), .C(n_579), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_628), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_628), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_664), .Y(n_752) );
OR2x2_ASAP7_75t_L g753 ( .A(n_638), .B(n_561), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_639), .B(n_575), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_639), .B(n_575), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_625), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_664), .Y(n_757) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_614), .B(n_558), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_618), .B(n_570), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_597), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_595), .B(n_553), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_584), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_677), .B(n_570), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_620), .B(n_553), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_677), .Y(n_765) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_678), .Y(n_766) );
INVx2_ASAP7_75t_SL g767 ( .A(n_598), .Y(n_767) );
NAND2x1p5_ASAP7_75t_L g768 ( .A(n_710), .B(n_598), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_696), .B(n_607), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g770 ( .A1(n_749), .A2(n_660), .B(n_644), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_766), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_766), .Y(n_772) );
A2O1A1Ixp33_ASAP7_75t_L g773 ( .A1(n_756), .A2(n_627), .B(n_598), .C(n_599), .Y(n_773) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_702), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_726), .A2(n_676), .B(n_607), .Y(n_775) );
OAI21xp33_ASAP7_75t_L g776 ( .A1(n_749), .A2(n_649), .B(n_666), .Y(n_776) );
OAI221xp5_ASAP7_75t_L g777 ( .A1(n_758), .A2(n_672), .B1(n_646), .B2(n_616), .C(n_541), .Y(n_777) );
AOI322xp5_ASAP7_75t_L g778 ( .A1(n_740), .A2(n_679), .A3(n_662), .B1(n_674), .B2(n_599), .C1(n_661), .C2(n_643), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_694), .Y(n_779) );
OAI22xp33_ASAP7_75t_L g780 ( .A1(n_730), .A2(n_646), .B1(n_616), .B2(n_599), .Y(n_780) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_765), .B(n_616), .C(n_675), .D(n_609), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_762), .B(n_635), .Y(n_782) );
OA222x2_ASAP7_75t_L g783 ( .A1(n_730), .A2(n_558), .B1(n_561), .B2(n_567), .C1(n_665), .C2(n_591), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_697), .B(n_630), .Y(n_784) );
OAI22xp33_ASAP7_75t_L g785 ( .A1(n_730), .A2(n_492), .B1(n_675), .B2(n_609), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_694), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_702), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_686), .B(n_680), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_732), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_733), .B(n_680), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_732), .Y(n_791) );
AO21x1_ASAP7_75t_L g792 ( .A1(n_736), .A2(n_675), .B(n_609), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_703), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_723), .B(n_659), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_703), .Y(n_795) );
OAI211xp5_ASAP7_75t_L g796 ( .A1(n_722), .A2(n_651), .B(n_652), .C(n_619), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_688), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_717), .B(n_670), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_722), .Y(n_799) );
OR2x2_ASAP7_75t_L g800 ( .A(n_753), .B(n_670), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_693), .Y(n_801) );
O2A1O1Ixp33_ASAP7_75t_L g802 ( .A1(n_735), .A2(n_567), .B(n_665), .C(n_658), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_745), .B(n_596), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_681), .A2(n_659), .B1(n_521), .B2(n_656), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_699), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_745), .B(n_596), .Y(n_806) );
INVx2_ASAP7_75t_SL g807 ( .A(n_767), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_717), .B(n_658), .Y(n_808) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_741), .Y(n_809) );
OR2x6_ASAP7_75t_L g810 ( .A(n_736), .B(n_659), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_701), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_704), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_705), .Y(n_813) );
OR2x2_ASAP7_75t_SL g814 ( .A(n_726), .B(n_656), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_725), .B(n_653), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_698), .B(n_653), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_698), .B(n_647), .Y(n_817) );
INVxp33_ASAP7_75t_L g818 ( .A(n_723), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_719), .A2(n_521), .B1(n_647), .B2(n_594), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_743), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_760), .B(n_594), .Y(n_821) );
AOI31xp33_ASAP7_75t_L g822 ( .A1(n_687), .A2(n_492), .A3(n_386), .B(n_548), .Y(n_822) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_740), .B(n_569), .Y(n_823) );
INVxp67_ASAP7_75t_L g824 ( .A(n_763), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_742), .A2(n_492), .B1(n_569), .B2(n_548), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_754), .B(n_540), .Y(n_826) );
INVx2_ASAP7_75t_L g827 ( .A(n_820), .Y(n_827) );
OAI21xp33_ASAP7_75t_L g828 ( .A1(n_770), .A2(n_684), .B(n_685), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_776), .A2(n_763), .B(n_739), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_779), .Y(n_830) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_822), .A2(n_746), .B1(n_734), .B2(n_687), .Y(n_831) );
AOI22x1_ASAP7_75t_L g832 ( .A1(n_768), .A2(n_742), .B1(n_744), .B2(n_690), .Y(n_832) );
AND2x2_ASAP7_75t_L g833 ( .A(n_794), .B(n_737), .Y(n_833) );
OAI22xp33_ASAP7_75t_SL g834 ( .A1(n_810), .A2(n_744), .B1(n_751), .B2(n_738), .Y(n_834) );
OAI21xp33_ASAP7_75t_L g835 ( .A1(n_776), .A2(n_689), .B(n_754), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_794), .B(n_683), .Y(n_836) );
AOI222xp33_ASAP7_75t_L g837 ( .A1(n_777), .A2(n_752), .B1(n_757), .B2(n_709), .C1(n_724), .C2(n_711), .Y(n_837) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_773), .A2(n_719), .B(n_759), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_818), .B(n_691), .Y(n_839) );
OAI22xp5_ASAP7_75t_L g840 ( .A1(n_814), .A2(n_755), .B1(n_692), .B2(n_695), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_786), .B(n_729), .Y(n_841) );
INVxp67_ASAP7_75t_L g842 ( .A(n_782), .Y(n_842) );
OAI21xp33_ASAP7_75t_SL g843 ( .A1(n_781), .A2(n_700), .B(n_715), .Y(n_843) );
OAI21xp5_ASAP7_75t_SL g844 ( .A1(n_804), .A2(n_761), .B(n_764), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_771), .B(n_747), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_796), .A2(n_682), .B1(n_755), .B2(n_713), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g847 ( .A1(n_775), .A2(n_750), .B(n_748), .Y(n_847) );
AOI321xp33_ASAP7_75t_L g848 ( .A1(n_785), .A2(n_759), .A3(n_707), .B1(n_731), .B2(n_728), .C(n_727), .Y(n_848) );
OA21x2_ASAP7_75t_L g849 ( .A1(n_774), .A2(n_743), .B(n_706), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g850 ( .A1(n_792), .A2(n_718), .B(n_716), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_772), .Y(n_851) );
AO22x1_ASAP7_75t_L g852 ( .A1(n_795), .A2(n_721), .B1(n_708), .B2(n_714), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_807), .A2(n_712), .B1(n_720), .B2(n_492), .Y(n_853) );
OAI32xp33_ASAP7_75t_L g854 ( .A1(n_824), .A2(n_565), .A3(n_540), .B1(n_539), .B2(n_499), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g855 ( .A1(n_810), .A2(n_539), .B1(n_488), .B2(n_499), .Y(n_855) );
O2A1O1Ixp33_ASAP7_75t_SL g856 ( .A1(n_780), .A2(n_418), .B(n_434), .C(n_450), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_789), .B(n_450), .Y(n_857) );
OAI221xp5_ASAP7_75t_SL g858 ( .A1(n_778), .A2(n_450), .B1(n_418), .B2(n_403), .C(n_434), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g859 ( .A1(n_804), .A2(n_403), .B(n_404), .C(n_409), .Y(n_859) );
AOI21xp33_ASAP7_75t_L g860 ( .A1(n_802), .A2(n_434), .B(n_82), .Y(n_860) );
OAI21xp5_ASAP7_75t_L g861 ( .A1(n_842), .A2(n_810), .B(n_819), .Y(n_861) );
INVxp67_ASAP7_75t_L g862 ( .A(n_839), .Y(n_862) );
OAI21xp33_ASAP7_75t_L g863 ( .A1(n_843), .A2(n_791), .B(n_821), .Y(n_863) );
AOI211xp5_ASAP7_75t_L g864 ( .A1(n_831), .A2(n_825), .B(n_819), .C(n_787), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g865 ( .A1(n_828), .A2(n_790), .B1(n_788), .B2(n_797), .C(n_811), .Y(n_865) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_844), .A2(n_805), .B1(n_801), .B2(n_812), .C(n_813), .Y(n_866) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_834), .A2(n_817), .B(n_816), .Y(n_867) );
OAI311xp33_ASAP7_75t_L g868 ( .A1(n_837), .A2(n_783), .A3(n_806), .B1(n_803), .C1(n_800), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_841), .Y(n_869) );
OAI221xp5_ASAP7_75t_L g870 ( .A1(n_848), .A2(n_798), .B1(n_808), .B2(n_793), .C(n_799), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_835), .B(n_840), .Y(n_871) );
AOI221xp5_ASAP7_75t_L g872 ( .A1(n_829), .A2(n_809), .B1(n_823), .B2(n_815), .C(n_826), .Y(n_872) );
AOI221xp5_ASAP7_75t_L g873 ( .A1(n_858), .A2(n_784), .B1(n_769), .B2(n_783), .C(n_442), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_852), .A2(n_434), .B(n_397), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_847), .A2(n_434), .B(n_397), .Y(n_875) );
AOI221xp5_ASAP7_75t_L g876 ( .A1(n_850), .A2(n_442), .B1(n_450), .B2(n_418), .C(n_434), .Y(n_876) );
OAI21xp5_ASAP7_75t_L g877 ( .A1(n_832), .A2(n_397), .B(n_450), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_830), .B(n_450), .Y(n_878) );
OAI321xp33_ASAP7_75t_L g879 ( .A1(n_855), .A2(n_442), .A3(n_450), .B1(n_86), .B2(n_87), .C(n_89), .Y(n_879) );
OAI211xp5_ASAP7_75t_L g880 ( .A1(n_873), .A2(n_838), .B(n_846), .C(n_853), .Y(n_880) );
NAND2xp33_ASAP7_75t_L g881 ( .A(n_863), .B(n_836), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_869), .Y(n_882) );
NAND2x1_ASAP7_75t_L g883 ( .A(n_861), .B(n_849), .Y(n_883) );
AOI211xp5_ASAP7_75t_SL g884 ( .A1(n_868), .A2(n_856), .B(n_860), .C(n_851), .Y(n_884) );
INVx1_ASAP7_75t_SL g885 ( .A(n_871), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_862), .B(n_857), .Y(n_886) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_866), .B(n_860), .C(n_854), .Y(n_887) );
NAND3xp33_ASAP7_75t_L g888 ( .A(n_864), .B(n_857), .C(n_849), .Y(n_888) );
AOI211xp5_ASAP7_75t_L g889 ( .A1(n_865), .A2(n_859), .B(n_841), .C(n_833), .Y(n_889) );
AND5x1_ASAP7_75t_L g890 ( .A(n_889), .B(n_872), .C(n_876), .D(n_867), .E(n_874), .Y(n_890) );
NOR3x1_ASAP7_75t_L g891 ( .A(n_880), .B(n_870), .C(n_878), .Y(n_891) );
A2O1A1Ixp33_ASAP7_75t_L g892 ( .A1(n_884), .A2(n_877), .B(n_879), .C(n_875), .Y(n_892) );
NOR2x1_ASAP7_75t_L g893 ( .A(n_885), .B(n_827), .Y(n_893) );
NAND3xp33_ASAP7_75t_L g894 ( .A(n_888), .B(n_845), .C(n_442), .Y(n_894) );
NOR3xp33_ASAP7_75t_SL g895 ( .A(n_886), .B(n_81), .C(n_85), .Y(n_895) );
OAI211xp5_ASAP7_75t_L g896 ( .A1(n_892), .A2(n_883), .B(n_887), .C(n_882), .Y(n_896) );
NAND4xp75_ASAP7_75t_L g897 ( .A(n_891), .B(n_881), .C(n_93), .D(n_94), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_893), .B(n_92), .Y(n_898) );
NAND3xp33_ASAP7_75t_L g899 ( .A(n_894), .B(n_442), .C(n_97), .Y(n_899) );
AND3x4_ASAP7_75t_L g900 ( .A(n_897), .B(n_895), .C(n_890), .Y(n_900) );
NOR2x1_ASAP7_75t_L g901 ( .A(n_896), .B(n_95), .Y(n_901) );
AOI22xp5_ASAP7_75t_L g902 ( .A1(n_898), .A2(n_442), .B1(n_101), .B2(n_104), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_901), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_900), .Y(n_904) );
NAND2xp5_ASAP7_75t_L g905 ( .A(n_904), .B(n_902), .Y(n_905) );
AO22x2_ASAP7_75t_L g906 ( .A1(n_903), .A2(n_899), .B1(n_106), .B2(n_107), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g907 ( .A1(n_905), .A2(n_903), .B1(n_442), .B2(n_110), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_906), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_908), .B(n_99), .Y(n_909) );
INVx2_ASAP7_75t_L g910 ( .A(n_909), .Y(n_910) );
XOR2xp5_ASAP7_75t_L g911 ( .A(n_910), .B(n_907), .Y(n_911) );
NAND2xp5_ASAP7_75t_SL g912 ( .A(n_911), .B(n_442), .Y(n_912) );
OR2x2_ASAP7_75t_L g913 ( .A(n_912), .B(n_109), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g914 ( .A1(n_913), .A2(n_114), .B1(n_116), .B2(n_117), .Y(n_914) );
endmodule