module fake_jpeg_2172_n_140 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_140);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_34),
.B1(n_48),
.B2(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_54),
.Y(n_57)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_40),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_36),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_36),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_47),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_52),
.B1(n_34),
.B2(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_78),
.Y(n_86)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_71),
.B(n_66),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_59),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_50),
.C(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_76),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22x1_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_54),
.B1(n_42),
.B2(n_39),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_67),
.B(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_92),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_68),
.B1(n_39),
.B2(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_89),
.B(n_90),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_60),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_3),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_3),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_4),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_80),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_100),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_85),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_9),
.C(n_10),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_105),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_72),
.C(n_75),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_6),
.C(n_8),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_70),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_111),
.B(n_19),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_86),
.B1(n_94),
.B2(n_39),
.Y(n_107)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_109),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_18),
.B1(n_33),
.B2(n_26),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_113),
.B1(n_9),
.B2(n_10),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_124),
.C(n_125),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_107),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_123),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_22),
.C(n_25),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_20),
.C(n_24),
.Y(n_125)
);

BUFx12f_ASAP7_75t_SL g128 ( 
.A(n_123),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_113),
.B(n_101),
.Y(n_133)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_97),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_121),
.C(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_120),
.C(n_126),
.Y(n_134)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_99),
.C(n_120),
.Y(n_136)
);

AOI322xp5_ASAP7_75t_L g137 ( 
.A1(n_136),
.A2(n_110),
.A3(n_135),
.B1(n_130),
.B2(n_119),
.C1(n_116),
.C2(n_13),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_130),
.C(n_106),
.Y(n_138)
);

AOI211xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_14),
.B(n_16),
.C(n_17),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_23),
.Y(n_140)
);


endmodule