module fake_jpeg_6503_n_103 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_39),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_0),
.C(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_64),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_0),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_46),
.Y(n_70)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_59),
.Y(n_77)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_51),
.B1(n_43),
.B2(n_57),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_74),
.A2(n_49),
.B1(n_42),
.B2(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_55),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_58),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_56),
.B(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_68),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_67),
.C(n_45),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_50),
.C(n_8),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_4),
.B(n_9),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_2),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_86),
.B(n_16),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_84),
.B1(n_18),
.B2(n_20),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_90),
.Y(n_94)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_87),
.B(n_92),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_17),
.C(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_23),
.C(n_24),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_98),
.A2(n_25),
.B(n_26),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_28),
.Y(n_101)
);

NOR4xp25_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_29),
.C(n_32),
.D(n_33),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_35),
.Y(n_103)
);


endmodule