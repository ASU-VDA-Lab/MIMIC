module fake_aes_12215_n_238 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_238);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_238;
wire n_117;
wire n_219;
wire n_133;
wire n_149;
wire n_220;
wire n_81;
wire n_214;
wire n_204;
wire n_221;
wire n_185;
wire n_203;
wire n_88;
wire n_102;
wire n_119;
wire n_141;
wire n_115;
wire n_97;
wire n_80;
wire n_167;
wire n_107;
wire n_158;
wire n_114;
wire n_121;
wire n_94;
wire n_171;
wire n_196;
wire n_125;
wire n_192;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_103;
wire n_137;
wire n_87;
wire n_180;
wire n_104;
wire n_160;
wire n_98;
wire n_206;
wire n_154;
wire n_195;
wire n_165;
wire n_146;
wire n_85;
wire n_237;
wire n_181;
wire n_101;
wire n_215;
wire n_108;
wire n_116;
wire n_155;
wire n_91;
wire n_209;
wire n_217;
wire n_139;
wire n_229;
wire n_230;
wire n_198;
wire n_169;
wire n_193;
wire n_152;
wire n_113;
wire n_95;
wire n_156;
wire n_124;
wire n_128;
wire n_129;
wire n_120;
wire n_90;
wire n_135;
wire n_188;
wire n_78;
wire n_201;
wire n_197;
wire n_127;
wire n_170;
wire n_111;
wire n_157;
wire n_79;
wire n_202;
wire n_210;
wire n_142;
wire n_184;
wire n_191;
wire n_232;
wire n_200;
wire n_208;
wire n_211;
wire n_122;
wire n_187;
wire n_138;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_84;
wire n_131;
wire n_112;
wire n_205;
wire n_86;
wire n_143;
wire n_213;
wire n_235;
wire n_182;
wire n_166;
wire n_162;
wire n_186;
wire n_75;
wire n_163;
wire n_226;
wire n_105;
wire n_159;
wire n_174;
wire n_227;
wire n_231;
wire n_136;
wire n_76;
wire n_89;
wire n_176;
wire n_144;
wire n_183;
wire n_77;
wire n_216;
wire n_147;
wire n_199;
wire n_148;
wire n_123;
wire n_83;
wire n_172;
wire n_100;
wire n_212;
wire n_228;
wire n_92;
wire n_223;
wire n_236;
wire n_150;
wire n_218;
wire n_168;
wire n_194;
wire n_110;
wire n_134;
wire n_222;
wire n_234;
wire n_164;
wire n_233;
wire n_82;
wire n_106;
wire n_175;
wire n_173;
wire n_190;
wire n_145;
wire n_153;
wire n_132;
wire n_99;
wire n_93;
wire n_109;
wire n_151;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_225;
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_21), .Y(n_75) );
BUFx5_ASAP7_75t_L g76 ( .A(n_7), .Y(n_76) );
BUFx2_ASAP7_75t_L g77 ( .A(n_56), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_48), .Y(n_78) );
INVxp67_ASAP7_75t_L g79 ( .A(n_52), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_67), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_26), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_47), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_71), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_6), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_70), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_32), .Y(n_88) );
INVx2_ASAP7_75t_SL g89 ( .A(n_43), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_5), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_33), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_66), .Y(n_92) );
BUFx2_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_58), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_14), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_25), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_62), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_31), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_7), .Y(n_101) );
BUFx8_ASAP7_75t_SL g102 ( .A(n_17), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_68), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_44), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_42), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_34), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_69), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_63), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_35), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_39), .B(n_22), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
INVx3_ASAP7_75t_L g114 ( .A(n_95), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_93), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_89), .B(n_0), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_76), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_102), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_106), .Y(n_120) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_85), .A2(n_16), .B(n_15), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_106), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_76), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_101), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_115), .B(n_79), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_114), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_117), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_119), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_125), .B(n_101), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_116), .B(n_79), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_118), .Y(n_132) );
INVx4_ASAP7_75t_L g133 ( .A(n_117), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_113), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_114), .B(n_110), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_114), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_127), .Y(n_137) );
AND2x6_ASAP7_75t_SL g138 ( .A(n_126), .B(n_86), .Y(n_138) );
AND2x6_ASAP7_75t_SL g139 ( .A(n_131), .B(n_90), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g140 ( .A(n_128), .B(n_113), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_128), .A2(n_123), .B1(n_96), .B2(n_98), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_127), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_136), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_128), .B(n_121), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_135), .B(n_75), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_130), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_133), .B(n_111), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_133), .B(n_78), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_147), .B(n_129), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_148), .B(n_132), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_145), .A2(n_134), .B(n_80), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_140), .A2(n_82), .B(n_81), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_149), .A2(n_84), .B(n_83), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_143), .Y(n_155) );
AOI21x1_ASAP7_75t_L g156 ( .A1(n_137), .A2(n_112), .B(n_87), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
OAI22xp5_ASAP7_75t_L g158 ( .A1(n_151), .A2(n_141), .B1(n_146), .B2(n_144), .Y(n_158) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_152), .A2(n_144), .B(n_88), .Y(n_159) );
AOI221xp5_ASAP7_75t_L g160 ( .A1(n_150), .A2(n_139), .B1(n_138), .B2(n_99), .C(n_100), .Y(n_160) );
AO31x2_ASAP7_75t_L g161 ( .A1(n_157), .A2(n_104), .A3(n_105), .B(n_103), .Y(n_161) );
AO31x2_ASAP7_75t_L g162 ( .A1(n_153), .A2(n_108), .A3(n_109), .B(n_107), .Y(n_162) );
BUFx5_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
AO21x1_ASAP7_75t_L g165 ( .A1(n_154), .A2(n_97), .B(n_91), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_161), .Y(n_166) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_164), .A2(n_94), .B(n_92), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_161), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_162), .Y(n_170) );
AO31x2_ASAP7_75t_L g171 ( .A1(n_165), .A2(n_122), .A3(n_124), .B(n_120), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_162), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_158), .A2(n_124), .B(n_19), .Y(n_173) );
AO21x2_ASAP7_75t_L g174 ( .A1(n_159), .A2(n_20), .B(n_18), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_163), .B(n_1), .Y(n_175) );
OAI211xp5_ASAP7_75t_L g176 ( .A1(n_160), .A2(n_4), .B(n_2), .C(n_3), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_170), .Y(n_177) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_172), .A2(n_24), .B(n_23), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_166), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_175), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_171), .Y(n_181) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_168), .A2(n_9), .B(n_10), .Y(n_182) );
OA21x2_ASAP7_75t_L g183 ( .A1(n_169), .A2(n_28), .B(n_27), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_171), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_174), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_174), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_176), .Y(n_187) );
BUFx2_ASAP7_75t_L g188 ( .A(n_167), .Y(n_188) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_12), .B(n_13), .Y(n_189) );
OA21x2_ASAP7_75t_L g190 ( .A1(n_170), .A2(n_30), .B(n_29), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_177), .Y(n_191) );
AO31x2_ASAP7_75t_L g192 ( .A1(n_185), .A2(n_36), .A3(n_37), .B(n_38), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_179), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_182), .Y(n_195) );
INVx1_ASAP7_75t_SL g196 ( .A(n_180), .Y(n_196) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_186), .A2(n_45), .B(n_46), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_180), .B(n_49), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_187), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_180), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_188), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_189), .Y(n_202) );
AO21x2_ASAP7_75t_L g203 ( .A1(n_184), .A2(n_50), .B(n_51), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_178), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_178), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_190), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_199), .B(n_183), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_191), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_193), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_191), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_200), .B(n_53), .Y(n_211) );
AND2x4_ASAP7_75t_L g212 ( .A(n_196), .B(n_54), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_201), .Y(n_213) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_194), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_195), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_196), .B(n_55), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_213), .B(n_202), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_209), .B(n_204), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_215), .B(n_205), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_214), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_208), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_207), .B(n_206), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_210), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_221), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_223), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_217), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_226), .B(n_220), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_227), .Y(n_228) );
AOI222xp33_ASAP7_75t_L g229 ( .A1(n_228), .A2(n_224), .B1(n_225), .B2(n_218), .C1(n_222), .C2(n_219), .Y(n_229) );
AOI22x1_ASAP7_75t_L g230 ( .A1(n_229), .A2(n_212), .B1(n_216), .B2(n_211), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_230), .Y(n_231) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_231), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_232), .Y(n_233) );
AOI22x1_ASAP7_75t_L g234 ( .A1(n_233), .A2(n_198), .B1(n_192), .B2(n_203), .Y(n_234) );
XNOR2xp5_ASAP7_75t_L g235 ( .A(n_234), .B(n_57), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_235), .A2(n_197), .B(n_59), .Y(n_236) );
OAI21xp5_ASAP7_75t_SL g237 ( .A1(n_236), .A2(n_60), .B(n_61), .Y(n_237) );
AOI21xp33_ASAP7_75t_SL g238 ( .A1(n_237), .A2(n_64), .B(n_65), .Y(n_238) );
endmodule