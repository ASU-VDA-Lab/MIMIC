module fake_jpeg_29916_n_131 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_7),
.B(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_51),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_61),
.B(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_21),
.C(n_39),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_1),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_1),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_55),
.B1(n_42),
.B2(n_43),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_70),
.B1(n_74),
.B2(n_47),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_71),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_55),
.B1(n_42),
.B2(n_43),
.Y(n_70)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_42),
.B1(n_54),
.B2(n_53),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_52),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_3),
.Y(n_88)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_6),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_49),
.B1(n_54),
.B2(n_46),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_79),
.A2(n_11),
.B1(n_17),
.B2(n_18),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_58),
.Y(n_80)
);

OAI32xp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_89),
.A3(n_11),
.B1(n_15),
.B2(n_16),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_58),
.B(n_61),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_65),
.C(n_66),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_2),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_3),
.B(n_4),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_88),
.C(n_10),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_23),
.B(n_38),
.C(n_37),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_6),
.Y(n_91)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_8),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_22),
.C(n_24),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_8),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_102),
.Y(n_109)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_66),
.B1(n_13),
.B2(n_14),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_105),
.B(n_41),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_19),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_106),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.C(n_113),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_96),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_26),
.C(n_28),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_29),
.C(n_30),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_31),
.B(n_34),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_120),
.C(n_122),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_95),
.C(n_104),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_101),
.B(n_103),
.C(n_93),
.D(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_112),
.C(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_108),
.C(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_126),
.Y(n_127)
);

OAI21x1_ASAP7_75t_L g128 ( 
.A1(n_127),
.A2(n_123),
.B(n_107),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_122),
.B(n_115),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_92),
.C(n_35),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_36),
.Y(n_131)
);


endmodule