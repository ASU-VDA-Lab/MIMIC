module real_aes_9755_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_2003;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_1034;
wire n_1328;
wire n_549;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_1346;
wire n_1383;
wire n_552;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_2004;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1914;
wire n_1648;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1812;
wire n_1769;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1638;
wire n_1078;
wire n_1072;
wire n_495;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1799;
wire n_1691;
wire n_640;
wire n_1931;
wire n_1176;
wire n_1721;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_892;
wire n_578;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_1252;
wire n_430;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_1705;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g921 ( .A1(n_0), .A2(n_539), .B1(n_922), .B2(n_924), .C(n_931), .Y(n_921) );
AOI21xp33_ASAP7_75t_L g956 ( .A1(n_0), .A2(n_744), .B(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_1), .A2(n_373), .B1(n_460), .B2(n_951), .Y(n_1385) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1), .Y(n_1408) );
INVx1_ASAP7_75t_L g1420 ( .A(n_2), .Y(n_1420) );
OAI221xp5_ASAP7_75t_L g1447 ( .A1(n_2), .A2(n_210), .B1(n_474), .B2(n_1448), .C(n_1449), .Y(n_1447) );
INVxp67_ASAP7_75t_L g1218 ( .A(n_3), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1251 ( .A1(n_3), .A2(n_223), .B1(n_722), .B2(n_1238), .C(n_1252), .Y(n_1251) );
INVx1_ASAP7_75t_L g882 ( .A(n_4), .Y(n_882) );
XNOR2x2_ASAP7_75t_L g1082 ( .A(n_5), .B(n_1083), .Y(n_1082) );
INVxp33_ASAP7_75t_L g1159 ( .A(n_6), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_6), .A2(n_119), .B1(n_1190), .B2(n_1191), .C(n_1192), .Y(n_1189) );
CKINVDCx5p33_ASAP7_75t_R g1581 ( .A(n_7), .Y(n_1581) );
OAI22xp5_ASAP7_75t_L g1974 ( .A1(n_8), .A2(n_84), .B1(n_1131), .B2(n_1975), .Y(n_1974) );
INVx1_ASAP7_75t_L g1986 ( .A(n_8), .Y(n_1986) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_9), .A2(n_284), .B1(n_1202), .B2(n_1204), .C(n_1206), .Y(n_1201) );
INVx1_ASAP7_75t_L g1247 ( .A(n_9), .Y(n_1247) );
INVx1_ASAP7_75t_L g1174 ( .A(n_10), .Y(n_1174) );
OAI221xp5_ASAP7_75t_L g934 ( .A1(n_11), .A2(n_206), .B1(n_526), .B2(n_532), .C(n_536), .Y(n_934) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_11), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g987 ( .A1(n_12), .A2(n_349), .B1(n_988), .B2(n_989), .C(n_991), .Y(n_987) );
INVx1_ASAP7_75t_L g1000 ( .A(n_12), .Y(n_1000) );
INVx1_ASAP7_75t_L g1737 ( .A(n_13), .Y(n_1737) );
CKINVDCx5p33_ASAP7_75t_R g1229 ( .A(n_14), .Y(n_1229) );
OAI22xp33_ASAP7_75t_L g1634 ( .A1(n_15), .A2(n_344), .B1(n_1129), .B2(n_1131), .Y(n_1634) );
INVx1_ASAP7_75t_L g1657 ( .A(n_15), .Y(n_1657) );
INVx1_ASAP7_75t_L g1982 ( .A(n_16), .Y(n_1982) );
OAI22xp5_ASAP7_75t_L g1996 ( .A1(n_16), .A2(n_105), .B1(n_910), .B2(n_915), .Y(n_1996) );
INVx1_ASAP7_75t_L g972 ( .A(n_17), .Y(n_972) );
AOI221xp5_ASAP7_75t_L g1917 ( .A1(n_18), .A2(n_38), .B1(n_828), .B2(n_1067), .C(n_1116), .Y(n_1917) );
INVx1_ASAP7_75t_L g1943 ( .A(n_18), .Y(n_1943) );
AOI22xp33_ASAP7_75t_SL g1040 ( .A1(n_19), .A2(n_175), .B1(n_782), .B2(n_1041), .Y(n_1040) );
AOI221xp5_ASAP7_75t_L g1064 ( .A1(n_19), .A2(n_279), .B1(n_835), .B2(n_1065), .C(n_1067), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_20), .A2(n_183), .B1(n_442), .B2(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g545 ( .A(n_20), .Y(n_545) );
OAI221xp5_ASAP7_75t_L g1211 ( .A1(n_21), .A2(n_136), .B1(n_524), .B2(n_536), .C(n_1212), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_21), .A2(n_136), .B1(n_791), .B2(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1971 ( .A(n_22), .Y(n_1971) );
OAI221xp5_ASAP7_75t_L g1988 ( .A1(n_22), .A2(n_899), .B1(n_1109), .B2(n_1989), .C(n_1990), .Y(n_1988) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_23), .A2(n_27), .B1(n_989), .B2(n_1088), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_23), .A2(n_312), .B1(n_915), .B2(n_1137), .Y(n_1136) );
CKINVDCx5p33_ASAP7_75t_R g845 ( .A(n_24), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_25), .A2(n_661), .B1(n_751), .B2(n_752), .Y(n_660) );
INVx1_ASAP7_75t_L g752 ( .A(n_25), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_26), .A2(n_225), .B1(n_810), .B2(n_1239), .Y(n_1632) );
OAI22xp5_ASAP7_75t_L g1636 ( .A1(n_26), .A2(n_225), .B1(n_1637), .B2(n_1638), .Y(n_1636) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_27), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1622 ( .A1(n_28), .A2(n_245), .B1(n_1623), .B2(n_1625), .Y(n_1622) );
INVxp67_ASAP7_75t_SL g1643 ( .A(n_28), .Y(n_1643) );
AOI22xp5_ASAP7_75t_L g1726 ( .A1(n_29), .A2(n_154), .B1(n_1675), .B2(n_1683), .Y(n_1726) );
INVx1_ASAP7_75t_L g699 ( .A(n_30), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g750 ( .A1(n_30), .A2(n_360), .B1(n_407), .B2(n_417), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_31), .A2(n_59), .B1(n_879), .B2(n_975), .C(n_976), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_31), .A2(n_320), .B1(n_1007), .B2(n_1008), .Y(n_1006) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_32), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1911 ( .A1(n_33), .A2(n_160), .B1(n_1623), .B2(n_1912), .Y(n_1911) );
INVx1_ASAP7_75t_L g1927 ( .A(n_33), .Y(n_1927) );
INVx1_ASAP7_75t_L g978 ( .A(n_34), .Y(n_978) );
AOI221xp5_ASAP7_75t_L g1002 ( .A1(n_34), .A2(n_59), .B1(n_718), .B2(n_1003), .C(n_1005), .Y(n_1002) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_35), .A2(n_357), .B1(n_1286), .B2(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g1313 ( .A(n_35), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_36), .A2(n_366), .B1(n_442), .B2(n_1013), .Y(n_1516) );
INVx1_ASAP7_75t_L g1549 ( .A(n_36), .Y(n_1549) );
CKINVDCx5p33_ASAP7_75t_R g1914 ( .A(n_37), .Y(n_1914) );
INVx1_ASAP7_75t_L g1938 ( .A(n_38), .Y(n_1938) );
OAI22xp5_ASAP7_75t_L g936 ( .A1(n_39), .A2(n_86), .B1(n_656), .B2(n_937), .Y(n_936) );
INVx1_ASAP7_75t_L g953 ( .A(n_39), .Y(n_953) );
INVx1_ASAP7_75t_L g1107 ( .A(n_40), .Y(n_1107) );
AOI221xp5_ASAP7_75t_L g1115 ( .A1(n_40), .A2(n_199), .B1(n_1116), .B2(n_1118), .C(n_1119), .Y(n_1115) );
INVx1_ASAP7_75t_L g993 ( .A(n_41), .Y(n_993) );
INVxp33_ASAP7_75t_L g1564 ( .A(n_42), .Y(n_1564) );
AOI221xp5_ASAP7_75t_L g1586 ( .A1(n_42), .A2(n_117), .B1(n_1587), .B2(n_1588), .C(n_1589), .Y(n_1586) );
AOI221xp5_ASAP7_75t_L g1327 ( .A1(n_43), .A2(n_269), .B1(n_433), .B2(n_602), .C(n_1328), .Y(n_1327) );
INVx1_ASAP7_75t_L g1353 ( .A(n_43), .Y(n_1353) );
AOI22xp33_ASAP7_75t_SL g1571 ( .A1(n_44), .A2(n_193), .B1(n_1572), .B2(n_1573), .Y(n_1571) );
AOI22xp33_ASAP7_75t_L g1599 ( .A1(n_44), .A2(n_193), .B1(n_1600), .B2(n_1601), .Y(n_1599) );
INVx1_ASAP7_75t_L g705 ( .A(n_45), .Y(n_705) );
OAI211xp5_ASAP7_75t_SL g709 ( .A1(n_45), .A2(n_710), .B(n_712), .C(n_723), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g1650 ( .A1(n_46), .A2(n_155), .B1(n_780), .B2(n_782), .C(n_1651), .Y(n_1650) );
OAI22xp5_ASAP7_75t_L g1660 ( .A1(n_46), .A2(n_180), .B1(n_1661), .B2(n_1663), .Y(n_1660) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_47), .A2(n_252), .B1(n_780), .B2(n_782), .Y(n_779) );
INVxp33_ASAP7_75t_SL g813 ( .A(n_47), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_48), .A2(n_334), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_48), .A2(n_152), .B1(n_807), .B2(n_809), .Y(n_806) );
INVx1_ASAP7_75t_L g380 ( .A(n_49), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g1747 ( .A1(n_50), .A2(n_146), .B1(n_1675), .B2(n_1683), .Y(n_1747) );
INVx1_ASAP7_75t_L g1146 ( .A(n_51), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_52), .A2(n_257), .B1(n_774), .B2(n_775), .Y(n_778) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_52), .Y(n_788) );
INVx1_ASAP7_75t_L g1508 ( .A(n_53), .Y(n_1508) );
CKINVDCx5p33_ASAP7_75t_R g1196 ( .A(n_54), .Y(n_1196) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_55), .A2(n_133), .B1(n_1281), .B2(n_1283), .Y(n_1280) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_55), .A2(n_236), .B1(n_742), .B2(n_1310), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1969 ( .A1(n_56), .A2(n_209), .B1(n_1587), .B2(n_1912), .Y(n_1969) );
INVx1_ASAP7_75t_L g1992 ( .A(n_56), .Y(n_1992) );
INVx1_ASAP7_75t_L g670 ( .A(n_57), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_57), .A2(n_311), .B1(n_742), .B2(n_745), .C(n_748), .Y(n_741) );
INVx1_ASAP7_75t_L g1111 ( .A(n_58), .Y(n_1111) );
CKINVDCx5p33_ASAP7_75t_R g1437 ( .A(n_60), .Y(n_1437) );
AOI22xp33_ASAP7_75t_SL g1575 ( .A1(n_61), .A2(n_338), .B1(n_1043), .B2(n_1576), .Y(n_1575) );
AOI221xp5_ASAP7_75t_L g1596 ( .A1(n_61), .A2(n_338), .B1(n_1328), .B2(n_1383), .C(n_1597), .Y(n_1596) );
INVx1_ASAP7_75t_L g1292 ( .A(n_62), .Y(n_1292) );
CKINVDCx5p33_ASAP7_75t_R g1485 ( .A(n_63), .Y(n_1485) );
INVx1_ASAP7_75t_L g1631 ( .A(n_64), .Y(n_1631) );
OAI211xp5_ASAP7_75t_SL g1645 ( .A1(n_64), .A2(n_859), .B(n_1646), .C(n_1652), .Y(n_1645) );
CKINVDCx5p33_ASAP7_75t_R g1275 ( .A(n_65), .Y(n_1275) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_66), .Y(n_1049) );
INVx1_ASAP7_75t_L g591 ( .A(n_67), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_67), .A2(n_318), .B1(n_624), .B2(n_625), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_68), .Y(n_1226) );
XOR2x2_ASAP7_75t_L g1020 ( .A(n_69), .B(n_1021), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_70), .A2(n_371), .B1(n_830), .B2(n_831), .Y(n_833) );
OAI22xp33_ASAP7_75t_L g898 ( .A1(n_70), .A2(n_353), .B1(n_899), .B2(n_901), .Y(n_898) );
AOI22xp33_ASAP7_75t_SL g1577 ( .A1(n_71), .A2(n_159), .B1(n_1043), .B2(n_1573), .Y(n_1577) );
INVxp67_ASAP7_75t_SL g1584 ( .A(n_71), .Y(n_1584) );
AOI22xp33_ASAP7_75t_L g1727 ( .A1(n_72), .A2(n_101), .B1(n_1691), .B2(n_1705), .Y(n_1727) );
INVx1_ASAP7_75t_L g1903 ( .A(n_72), .Y(n_1903) );
AOI22xp33_ASAP7_75t_L g1953 ( .A1(n_72), .A2(n_1954), .B1(n_1958), .B2(n_2000), .Y(n_1953) );
INVxp33_ASAP7_75t_L g1144 ( .A(n_73), .Y(n_1144) );
AOI221xp5_ASAP7_75t_L g1181 ( .A1(n_73), .A2(n_143), .B1(n_1182), .B2(n_1184), .C(n_1186), .Y(n_1181) );
CKINVDCx5p33_ASAP7_75t_R g1034 ( .A(n_74), .Y(n_1034) );
INVx1_ASAP7_75t_L g971 ( .A(n_75), .Y(n_971) );
INVxp33_ASAP7_75t_SL g1035 ( .A(n_76), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_76), .A2(n_274), .B1(n_1056), .B2(n_1058), .C(n_1059), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g1230 ( .A(n_77), .Y(n_1230) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_78), .A2(n_198), .B1(n_894), .B2(n_930), .Y(n_933) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_78), .A2(n_198), .B1(n_407), .B2(n_423), .Y(n_941) );
INVxp33_ASAP7_75t_L g1156 ( .A(n_79), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1193 ( .A1(n_79), .A2(n_310), .B1(n_716), .B2(n_1194), .Y(n_1193) );
OAI221xp5_ASAP7_75t_L g1150 ( .A1(n_80), .A2(n_254), .B1(n_535), .B2(n_677), .C(n_1151), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1179 ( .A1(n_80), .A2(n_254), .B1(n_791), .B2(n_1180), .Y(n_1179) );
OAI221xp5_ASAP7_75t_L g1102 ( .A1(n_81), .A2(n_899), .B1(n_1103), .B2(n_1106), .C(n_1109), .Y(n_1102) );
AOI221xp5_ASAP7_75t_L g1121 ( .A1(n_81), .A2(n_261), .B1(n_830), .B2(n_1065), .C(n_1122), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1699 ( .A1(n_82), .A2(n_232), .B1(n_1675), .B2(n_1683), .Y(n_1699) );
AOI22xp33_ASAP7_75t_SL g1042 ( .A1(n_83), .A2(n_279), .B1(n_1043), .B2(n_1044), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_83), .A2(n_175), .B1(n_1013), .B2(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1987 ( .A(n_84), .Y(n_1987) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_85), .A2(n_122), .B1(n_524), .B2(n_677), .C(n_678), .Y(n_676) );
INVx1_ASAP7_75t_L g737 ( .A(n_85), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_86), .A2(n_145), .B1(n_432), .B2(n_951), .Y(n_955) );
AO22x1_ASAP7_75t_SL g1717 ( .A1(n_87), .A2(n_156), .B1(n_1675), .B2(n_1683), .Y(n_1717) );
CKINVDCx5p33_ASAP7_75t_R g1519 ( .A(n_88), .Y(n_1519) );
INVxp67_ASAP7_75t_SL g1028 ( .A(n_89), .Y(n_1028) );
OAI22xp33_ASAP7_75t_L g1053 ( .A1(n_89), .A2(n_321), .B1(n_735), .B2(n_1054), .Y(n_1053) );
XOR2xp5_ASAP7_75t_L g820 ( .A(n_90), .B(n_821), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_91), .Y(n_1388) );
CKINVDCx5p33_ASAP7_75t_R g1324 ( .A(n_92), .Y(n_1324) );
INVx1_ASAP7_75t_L g1032 ( .A(n_93), .Y(n_1032) );
INVx1_ASAP7_75t_L g880 ( .A(n_94), .Y(n_880) );
AOI22xp33_ASAP7_75t_SL g1578 ( .A1(n_95), .A2(n_140), .B1(n_1572), .B2(n_1576), .Y(n_1578) );
INVxp67_ASAP7_75t_L g1595 ( .A(n_95), .Y(n_1595) );
INVx1_ASAP7_75t_L g1440 ( .A(n_96), .Y(n_1440) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_96), .A2(n_339), .B1(n_432), .B2(n_449), .Y(n_1450) );
CKINVDCx5p33_ASAP7_75t_R g1227 ( .A(n_97), .Y(n_1227) );
AOI22xp33_ASAP7_75t_SL g1423 ( .A1(n_98), .A2(n_207), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
AOI22xp33_ASAP7_75t_L g1456 ( .A1(n_98), .A2(n_208), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
INVx1_ASAP7_75t_L g1522 ( .A(n_99), .Y(n_1522) );
OAI221xp5_ASAP7_75t_L g1538 ( .A1(n_99), .A2(n_164), .B1(n_532), .B2(n_1151), .C(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1531 ( .A(n_100), .Y(n_1531) );
CKINVDCx5p33_ASAP7_75t_R g1919 ( .A(n_102), .Y(n_1919) );
CKINVDCx5p33_ASAP7_75t_R g1527 ( .A(n_103), .Y(n_1527) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_104), .A2(n_337), .B1(n_809), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g863 ( .A(n_104), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g1983 ( .A1(n_105), .A2(n_364), .B1(n_770), .B2(n_1651), .C(n_1984), .Y(n_1983) );
AOI22xp5_ASAP7_75t_L g1700 ( .A1(n_106), .A2(n_248), .B1(n_1687), .B2(n_1691), .Y(n_1700) );
INVx1_ASAP7_75t_L g1269 ( .A(n_107), .Y(n_1269) );
OAI22xp5_ASAP7_75t_L g1296 ( .A1(n_107), .A2(n_192), .B1(n_1054), .B2(n_1297), .Y(n_1296) );
OAI22xp5_ASAP7_75t_L g1915 ( .A1(n_108), .A2(n_271), .B1(n_1054), .B2(n_1297), .Y(n_1915) );
OAI221xp5_ASAP7_75t_L g1933 ( .A1(n_108), .A2(n_271), .B1(n_677), .B2(n_678), .C(n_1151), .Y(n_1933) );
INVx1_ASAP7_75t_L g1972 ( .A(n_109), .Y(n_1972) );
OAI211xp5_ASAP7_75t_L g1978 ( .A1(n_109), .A2(n_859), .B(n_1979), .C(n_1985), .Y(n_1978) );
INVx1_ASAP7_75t_L g1487 ( .A(n_110), .Y(n_1487) );
OAI211xp5_ASAP7_75t_SL g604 ( .A1(n_111), .A2(n_605), .B(n_606), .C(n_609), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_111), .A2(n_216), .B1(n_628), .B2(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g1528 ( .A1(n_112), .A2(n_243), .B1(n_462), .B2(n_1011), .C(n_1473), .Y(n_1528) );
INVx1_ASAP7_75t_L g1537 ( .A(n_112), .Y(n_1537) );
AOI22xp33_ASAP7_75t_L g1973 ( .A1(n_113), .A2(n_251), .B1(n_810), .B2(n_1239), .Y(n_1973) );
OAI22xp5_ASAP7_75t_L g1993 ( .A1(n_113), .A2(n_251), .B1(n_1637), .B2(n_1638), .Y(n_1993) );
CKINVDCx5p33_ASAP7_75t_R g674 ( .A(n_114), .Y(n_674) );
INVx1_ASAP7_75t_L g1377 ( .A(n_115), .Y(n_1377) );
OAI221xp5_ASAP7_75t_L g1400 ( .A1(n_115), .A2(n_137), .B1(n_531), .B2(n_535), .C(n_1344), .Y(n_1400) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_116), .Y(n_688) );
INVxp33_ASAP7_75t_SL g1568 ( .A(n_117), .Y(n_1568) );
AOI22xp5_ASAP7_75t_L g1686 ( .A1(n_118), .A2(n_135), .B1(n_1687), .B2(n_1691), .Y(n_1686) );
INVxp67_ASAP7_75t_L g1161 ( .A(n_119), .Y(n_1161) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_120), .A2(n_270), .B1(n_433), .B2(n_462), .C(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1494 ( .A(n_120), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_121), .A2(n_363), .B1(n_469), .B2(n_474), .Y(n_468) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_121), .A2(n_363), .B1(n_524), .B2(n_531), .C(n_535), .Y(n_523) );
INVx1_ASAP7_75t_L g733 ( .A(n_122), .Y(n_733) );
BUFx2_ASAP7_75t_L g481 ( .A(n_123), .Y(n_481) );
OR2x2_ASAP7_75t_L g486 ( .A(n_123), .B(n_487), .Y(n_486) );
BUFx2_ASAP7_75t_L g490 ( .A(n_123), .Y(n_490) );
INVx1_ASAP7_75t_L g502 ( .A(n_123), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g929 ( .A1(n_124), .A2(n_168), .B1(n_894), .B2(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g947 ( .A(n_124), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_125), .Y(n_1387) );
INVx1_ASAP7_75t_L g1712 ( .A(n_126), .Y(n_1712) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_127), .A2(n_130), .B1(n_1432), .B2(n_1434), .Y(n_1431) );
INVx1_ASAP7_75t_L g1460 ( .A(n_127), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1695 ( .A1(n_128), .A2(n_325), .B1(n_1675), .B2(n_1683), .Y(n_1695) );
AOI22xp33_ASAP7_75t_SL g1046 ( .A1(n_129), .A2(n_231), .B1(n_1043), .B2(n_1044), .Y(n_1046) );
INVxp33_ASAP7_75t_SL g1073 ( .A(n_129), .Y(n_1073) );
INVx1_ASAP7_75t_L g1454 ( .A(n_130), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g1748 ( .A1(n_131), .A2(n_293), .B1(n_1691), .B2(n_1705), .Y(n_1748) );
AOI22xp33_ASAP7_75t_L g1918 ( .A1(n_132), .A2(n_294), .B1(n_1058), .B2(n_1070), .Y(n_1918) );
INVx1_ASAP7_75t_L g1944 ( .A(n_132), .Y(n_1944) );
AOI221xp5_ASAP7_75t_L g1305 ( .A1(n_133), .A2(n_306), .B1(n_602), .B2(n_1306), .C(n_1308), .Y(n_1305) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_134), .A2(n_218), .B1(n_431), .B2(n_433), .C(n_436), .Y(n_430) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_134), .Y(n_558) );
INVx1_ASAP7_75t_L g1378 ( .A(n_137), .Y(n_1378) );
AOI22xp33_ASAP7_75t_SL g1047 ( .A1(n_138), .A2(n_292), .B1(n_782), .B2(n_1041), .Y(n_1047) );
INVxp33_ASAP7_75t_L g1072 ( .A(n_138), .Y(n_1072) );
INVx1_ASAP7_75t_L g1276 ( .A(n_139), .Y(n_1276) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_139), .A2(n_149), .B1(n_1058), .B2(n_1300), .C(n_1302), .Y(n_1299) );
INVxp33_ASAP7_75t_L g1603 ( .A(n_140), .Y(n_1603) );
INVx1_ASAP7_75t_L g1628 ( .A(n_141), .Y(n_1628) );
OAI221xp5_ASAP7_75t_L g1639 ( .A1(n_141), .A2(n_899), .B1(n_1109), .B2(n_1640), .C(n_1642), .Y(n_1639) );
INVx1_ASAP7_75t_L g992 ( .A(n_142), .Y(n_992) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_142), .A2(n_349), .B1(n_467), .B2(n_997), .C(n_999), .Y(n_996) );
INVxp33_ASAP7_75t_L g1149 ( .A(n_143), .Y(n_1149) );
NAND2xp33_ASAP7_75t_SL g1375 ( .A(n_144), .B(n_1254), .Y(n_1375) );
INVx1_ASAP7_75t_L g1396 ( .A(n_144), .Y(n_1396) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_145), .A2(n_165), .B1(n_485), .B2(n_655), .Y(n_938) );
INVx1_ASAP7_75t_L g1265 ( .A(n_146), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1959 ( .A1(n_147), .A2(n_1960), .B1(n_1998), .B2(n_1999), .Y(n_1959) );
CKINVDCx14_ASAP7_75t_R g1998 ( .A(n_147), .Y(n_1998) );
INVx1_ASAP7_75t_L g1720 ( .A(n_148), .Y(n_1720) );
INVx1_ASAP7_75t_L g1272 ( .A(n_149), .Y(n_1272) );
INVx1_ASAP7_75t_L g1567 ( .A(n_150), .Y(n_1567) );
INVx1_ASAP7_75t_L g1207 ( .A(n_151), .Y(n_1207) );
AOI22xp33_ASAP7_75t_SL g768 ( .A1(n_152), .A2(n_308), .B1(n_769), .B2(n_771), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_153), .A2(n_187), .B1(n_433), .B2(n_460), .C(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g511 ( .A(n_153), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g1659 ( .A1(n_155), .A2(n_229), .B1(n_910), .B2(n_915), .Y(n_1659) );
INVx1_ASAP7_75t_L g816 ( .A(n_156), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g1334 ( .A(n_157), .Y(n_1334) );
CKINVDCx5p33_ASAP7_75t_R g1486 ( .A(n_158), .Y(n_1486) );
INVxp33_ASAP7_75t_L g1604 ( .A(n_159), .Y(n_1604) );
INVx1_ASAP7_75t_L g1932 ( .A(n_160), .Y(n_1932) );
CKINVDCx5p33_ASAP7_75t_R g1333 ( .A(n_161), .Y(n_1333) );
INVx1_ASAP7_75t_L g1464 ( .A(n_162), .Y(n_1464) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_163), .Y(n_608) );
INVx1_ASAP7_75t_L g1521 ( .A(n_164), .Y(n_1521) );
INVx1_ASAP7_75t_L g959 ( .A(n_165), .Y(n_959) );
INVxp67_ASAP7_75t_SL g1561 ( .A(n_166), .Y(n_1561) );
OAI22xp33_ASAP7_75t_L g1585 ( .A1(n_166), .A2(n_196), .B1(n_791), .B2(n_1236), .Y(n_1585) );
INVx1_ASAP7_75t_L g429 ( .A(n_167), .Y(n_429) );
INVx1_ASAP7_75t_L g944 ( .A(n_168), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g1480 ( .A1(n_169), .A2(n_273), .B1(n_436), .B2(n_1124), .C(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1503 ( .A(n_169), .Y(n_1503) );
AOI21xp33_ASAP7_75t_L g600 ( .A1(n_170), .A2(n_601), .B(n_602), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_170), .A2(n_195), .B1(n_628), .B2(n_630), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g1612 ( .A(n_171), .Y(n_1612) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_172), .A2(n_216), .B1(n_407), .B2(n_417), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_172), .A2(n_299), .B1(n_625), .B2(n_637), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g1330 ( .A(n_173), .Y(n_1330) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_174), .Y(n_607) );
INVx1_ASAP7_75t_L g1104 ( .A(n_176), .Y(n_1104) );
INVx1_ASAP7_75t_L g1679 ( .A(n_177), .Y(n_1679) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_178), .A2(n_312), .B1(n_887), .B2(n_1091), .C(n_1093), .Y(n_1090) );
INVxp67_ASAP7_75t_SL g1135 ( .A(n_178), .Y(n_1135) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_179), .Y(n_684) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_179), .A2(n_343), .B1(n_718), .B2(n_720), .C(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g1648 ( .A(n_180), .Y(n_1648) );
CKINVDCx5p33_ASAP7_75t_R g1471 ( .A(n_181), .Y(n_1471) );
INVx1_ASAP7_75t_L g1148 ( .A(n_182), .Y(n_1148) );
INVx1_ASAP7_75t_L g561 ( .A(n_183), .Y(n_561) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_184), .A2(n_401), .B1(n_581), .B2(n_582), .Y(n_400) );
INVx1_ASAP7_75t_L g582 ( .A(n_184), .Y(n_582) );
INVx1_ASAP7_75t_L g1439 ( .A(n_185), .Y(n_1439) );
AOI21xp33_ASAP7_75t_L g1451 ( .A1(n_185), .A2(n_797), .B(n_957), .Y(n_1451) );
AOI221xp5_ASAP7_75t_L g1703 ( .A1(n_186), .A2(n_266), .B1(n_1704), .B2(n_1706), .C(n_1708), .Y(n_1703) );
INVx1_ASAP7_75t_L g505 ( .A(n_187), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g1374 ( .A1(n_188), .A2(n_332), .B1(n_810), .B2(n_1240), .Y(n_1374) );
INVx1_ASAP7_75t_L g1395 ( .A(n_188), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_189), .A2(n_237), .B1(n_465), .B2(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g495 ( .A(n_189), .Y(n_495) );
INVx1_ASAP7_75t_L g1680 ( .A(n_190), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1685 ( .A(n_190), .B(n_1678), .Y(n_1685) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_191), .A2(n_224), .B1(n_457), .B2(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1338 ( .A(n_191), .Y(n_1338) );
INVx1_ASAP7_75t_L g1270 ( .A(n_192), .Y(n_1270) );
INVx2_ASAP7_75t_L g392 ( .A(n_194), .Y(n_392) );
INVx1_ASAP7_75t_L g594 ( .A(n_195), .Y(n_594) );
INVxp67_ASAP7_75t_SL g1562 ( .A(n_196), .Y(n_1562) );
AO221x2_ASAP7_75t_L g1733 ( .A1(n_197), .A2(n_239), .B1(n_1705), .B2(n_1734), .C(n_1735), .Y(n_1733) );
AOI21xp33_ASAP7_75t_L g1108 ( .A1(n_199), .A2(n_540), .B(n_1091), .Y(n_1108) );
CKINVDCx5p33_ASAP7_75t_R g1273 ( .A(n_200), .Y(n_1273) );
INVx1_ASAP7_75t_L g412 ( .A(n_201), .Y(n_412) );
BUFx3_ASAP7_75t_L g427 ( .A(n_201), .Y(n_427) );
XNOR2x2_ASAP7_75t_L g1198 ( .A(n_202), .B(n_1199), .Y(n_1198) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_203), .A2(n_662), .B(n_664), .C(n_708), .Y(n_661) );
INVx1_ASAP7_75t_L g877 ( .A(n_204), .Y(n_877) );
INVxp67_ASAP7_75t_L g1224 ( .A(n_205), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_205), .A2(n_290), .B1(n_830), .B2(n_1256), .Y(n_1255) );
CKINVDCx5p33_ASAP7_75t_R g964 ( .A(n_206), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g1455 ( .A1(n_207), .A2(n_313), .B1(n_431), .B2(n_433), .C(n_1005), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_208), .A2(n_313), .B1(n_1427), .B2(n_1428), .Y(n_1426) );
INVx1_ASAP7_75t_L g1991 ( .A(n_209), .Y(n_1991) );
INVx1_ASAP7_75t_L g1419 ( .A(n_210), .Y(n_1419) );
AOI221xp5_ASAP7_75t_L g1381 ( .A1(n_211), .A2(n_297), .B1(n_431), .B2(n_1382), .C(n_1383), .Y(n_1381) );
INVx1_ASAP7_75t_L g1403 ( .A(n_211), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g1475 ( .A1(n_212), .A2(n_314), .B1(n_790), .B2(n_1476), .Y(n_1475) );
OAI221xp5_ASAP7_75t_L g1496 ( .A1(n_212), .A2(n_314), .B1(n_531), .B2(n_536), .C(n_1344), .Y(n_1496) );
INVx1_ASAP7_75t_L g1167 ( .A(n_213), .Y(n_1167) );
INVx1_ASAP7_75t_L g979 ( .A(n_214), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g1908 ( .A1(n_215), .A2(n_226), .B1(n_748), .B2(n_1909), .C(n_1910), .Y(n_1908) );
INVx1_ASAP7_75t_L g1931 ( .A(n_215), .Y(n_1931) );
INVx1_ASAP7_75t_L g1105 ( .A(n_217), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g552 ( .A(n_218), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_219), .A2(n_353), .B1(n_835), .B2(n_836), .Y(n_834) );
OAI22xp33_ASAP7_75t_L g854 ( .A1(n_219), .A2(n_371), .B1(n_855), .B2(n_859), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_220), .Y(n_850) );
INVxp33_ASAP7_75t_SL g761 ( .A(n_221), .Y(n_761) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_221), .A2(n_264), .B1(n_593), .B2(n_601), .Y(n_795) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_222), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_222), .A2(n_265), .B1(n_790), .B2(n_791), .C(n_793), .Y(n_789) );
INVxp67_ASAP7_75t_L g1222 ( .A(n_223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1342 ( .A(n_224), .Y(n_1342) );
INVx1_ASAP7_75t_L g1929 ( .A(n_226), .Y(n_1929) );
INVx1_ASAP7_75t_L g409 ( .A(n_227), .Y(n_409) );
INVx1_ASAP7_75t_L g439 ( .A(n_227), .Y(n_439) );
INVx1_ASAP7_75t_L g415 ( .A(n_228), .Y(n_415) );
INVx1_ASAP7_75t_L g1649 ( .A(n_229), .Y(n_1649) );
INVx1_ASAP7_75t_L g1565 ( .A(n_230), .Y(n_1565) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_231), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_233), .Y(n_1332) );
CKINVDCx20_ASAP7_75t_R g1369 ( .A(n_234), .Y(n_1369) );
OAI21xp33_ASAP7_75t_L g968 ( .A1(n_235), .A2(n_969), .B(n_994), .Y(n_968) );
INVx1_ASAP7_75t_L g1019 ( .A(n_235), .Y(n_1019) );
AOI22xp33_ASAP7_75t_SL g1284 ( .A1(n_236), .A2(n_306), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
INVx1_ASAP7_75t_L g516 ( .A(n_237), .Y(n_516) );
OA22x2_ASAP7_75t_L g1314 ( .A1(n_238), .A2(n_1315), .B1(n_1360), .B2(n_1361), .Y(n_1314) );
INVx1_ASAP7_75t_L g1361 ( .A(n_238), .Y(n_1361) );
XOR2xp5_ASAP7_75t_L g918 ( .A(n_240), .B(n_919), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g1674 ( .A1(n_240), .A2(n_301), .B1(n_1675), .B2(n_1683), .Y(n_1674) );
INVx1_ASAP7_75t_L g1139 ( .A(n_241), .Y(n_1139) );
AOI22xp5_ASAP7_75t_L g1696 ( .A1(n_242), .A2(n_324), .B1(n_1687), .B2(n_1691), .Y(n_1696) );
INVx1_ASAP7_75t_L g1535 ( .A(n_243), .Y(n_1535) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_244), .A2(n_304), .B1(n_593), .B2(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g654 ( .A1(n_244), .A2(n_367), .B1(n_655), .B2(n_656), .Y(n_654) );
INVxp67_ASAP7_75t_SL g1644 ( .A(n_245), .Y(n_1644) );
INVx1_ASAP7_75t_L g986 ( .A(n_246), .Y(n_986) );
AOI221xp5_ASAP7_75t_L g1010 ( .A1(n_246), .A2(n_322), .B1(n_808), .B2(n_957), .C(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g1981 ( .A(n_247), .Y(n_1981) );
OAI22xp5_ASAP7_75t_L g1997 ( .A1(n_247), .A2(n_364), .B1(n_1661), .B2(n_1663), .Y(n_1997) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_249), .Y(n_1514) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_250), .Y(n_885) );
INVxp67_ASAP7_75t_SL g799 ( .A(n_252), .Y(n_799) );
INVx1_ASAP7_75t_L g1175 ( .A(n_253), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_255), .A2(n_340), .B1(n_1096), .B2(n_1098), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g1128 ( .A1(n_255), .A2(n_340), .B1(n_1129), .B2(n_1131), .C(n_1132), .Y(n_1128) );
INVx1_ASAP7_75t_L g482 ( .A(n_256), .Y(n_482) );
INVxp33_ASAP7_75t_SL g814 ( .A(n_257), .Y(n_814) );
INVx1_ASAP7_75t_L g1721 ( .A(n_258), .Y(n_1721) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_259), .A2(n_278), .B1(n_830), .B2(n_831), .Y(n_829) );
INVx1_ASAP7_75t_L g872 ( .A(n_259), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g1462 ( .A(n_260), .Y(n_1462) );
OAI211xp5_ASAP7_75t_L g1085 ( .A1(n_261), .A2(n_859), .B(n_1086), .C(n_1099), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g1736 ( .A(n_262), .Y(n_1736) );
INVx1_ASAP7_75t_L g1100 ( .A(n_263), .Y(n_1100) );
INVxp33_ASAP7_75t_SL g766 ( .A(n_264), .Y(n_766) );
INVxp67_ASAP7_75t_SL g758 ( .A(n_265), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g1518 ( .A(n_267), .Y(n_1518) );
INVx1_ASAP7_75t_L g690 ( .A(n_268), .Y(n_690) );
INVx1_ASAP7_75t_L g1349 ( .A(n_269), .Y(n_1349) );
INVx1_ASAP7_75t_L g1492 ( .A(n_270), .Y(n_1492) );
OAI22xp5_ASAP7_75t_L g1325 ( .A1(n_272), .A2(n_276), .B1(n_474), .B2(n_790), .Y(n_1325) );
OAI221xp5_ASAP7_75t_L g1343 ( .A1(n_272), .A2(n_276), .B1(n_531), .B2(n_535), .C(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1500 ( .A(n_273), .Y(n_1500) );
INVxp33_ASAP7_75t_SL g1030 ( .A(n_274), .Y(n_1030) );
INVx1_ASAP7_75t_L g695 ( .A(n_275), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g728 ( .A1(n_275), .A2(n_729), .B(n_731), .C(n_738), .Y(n_728) );
INVx1_ASAP7_75t_L g1923 ( .A(n_277), .Y(n_1923) );
INVx1_ASAP7_75t_L g868 ( .A(n_278), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g1921 ( .A(n_280), .Y(n_1921) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_281), .Y(n_667) );
INVx1_ASAP7_75t_L g1101 ( .A(n_282), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g1319 ( .A1(n_283), .A2(n_298), .B1(n_433), .B2(n_1320), .C(n_1321), .Y(n_1319) );
INVx1_ASAP7_75t_L g1339 ( .A(n_283), .Y(n_1339) );
AOI221xp5_ASAP7_75t_L g1237 ( .A1(n_284), .A2(n_369), .B1(n_1238), .B2(n_1241), .C(n_1244), .Y(n_1237) );
AOI22xp33_ASAP7_75t_L g1483 ( .A1(n_285), .A2(n_315), .B1(n_951), .B2(n_1457), .Y(n_1483) );
INVx1_ASAP7_75t_L g1504 ( .A(n_285), .Y(n_1504) );
CKINVDCx20_ASAP7_75t_R g1605 ( .A(n_286), .Y(n_1605) );
INVx1_ASAP7_75t_L g1621 ( .A(n_287), .Y(n_1621) );
INVx1_ASAP7_75t_L g414 ( .A(n_288), .Y(n_414) );
BUFx3_ASAP7_75t_L g420 ( .A(n_288), .Y(n_420) );
INVx1_ASAP7_75t_L g785 ( .A(n_289), .Y(n_785) );
INVxp67_ASAP7_75t_L g1216 ( .A(n_290), .Y(n_1216) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_291), .A2(n_460), .B(n_462), .Y(n_614) );
INVx1_ASAP7_75t_L g651 ( .A(n_291), .Y(n_651) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_292), .Y(n_1063) );
INVx1_ASAP7_75t_L g1936 ( .A(n_294), .Y(n_1936) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_295), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_295), .B(n_354), .Y(n_487) );
AND2x2_ASAP7_75t_L g503 ( .A(n_295), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g580 ( .A(n_295), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g1515 ( .A1(n_296), .A2(n_342), .B1(n_601), .B2(n_1011), .C(n_1383), .Y(n_1515) );
INVx1_ASAP7_75t_L g1544 ( .A(n_296), .Y(n_1544) );
INVx1_ASAP7_75t_L g1409 ( .A(n_297), .Y(n_1409) );
INVx1_ASAP7_75t_L g1341 ( .A(n_298), .Y(n_1341) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_299), .A2(n_423), .B1(n_588), .B2(n_595), .C(n_603), .Y(n_587) );
OR2x2_ASAP7_75t_L g408 ( .A(n_300), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g440 ( .A(n_300), .Y(n_440) );
INVx1_ASAP7_75t_L g1554 ( .A(n_302), .Y(n_1554) );
CKINVDCx5p33_ASAP7_75t_R g1922 ( .A(n_303), .Y(n_1922) );
INVx1_ASAP7_75t_L g653 ( .A(n_304), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_305), .A2(n_319), .B1(n_519), .B2(n_567), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_305), .A2(n_319), .B1(n_417), .B2(n_605), .Y(n_940) );
INVx1_ASAP7_75t_L g926 ( .A(n_307), .Y(n_926) );
AOI21xp33_ASAP7_75t_L g945 ( .A1(n_307), .A2(n_431), .B(n_602), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_308), .A2(n_334), .B1(n_602), .B2(n_801), .C(n_803), .Y(n_800) );
CKINVDCx5p33_ASAP7_75t_R g1525 ( .A(n_309), .Y(n_1525) );
INVxp67_ASAP7_75t_L g1164 ( .A(n_310), .Y(n_1164) );
INVx1_ASAP7_75t_L g673 ( .A(n_311), .Y(n_673) );
INVx1_ASAP7_75t_L g1499 ( .A(n_315), .Y(n_1499) );
AOI22xp33_ASAP7_75t_SL g1290 ( .A1(n_316), .A2(n_317), .B1(n_782), .B2(n_1041), .Y(n_1290) );
INVx1_ASAP7_75t_L g1304 ( .A(n_316), .Y(n_1304) );
INVx1_ASAP7_75t_L g1312 ( .A(n_317), .Y(n_1312) );
INVx1_ASAP7_75t_L g596 ( .A(n_318), .Y(n_596) );
INVxp67_ASAP7_75t_SL g977 ( .A(n_320), .Y(n_977) );
INVxp67_ASAP7_75t_SL g1025 ( .A(n_321), .Y(n_1025) );
INVx1_ASAP7_75t_L g985 ( .A(n_322), .Y(n_985) );
INVxp33_ASAP7_75t_SL g765 ( .A(n_323), .Y(n_765) );
AOI21xp33_ASAP7_75t_L g796 ( .A1(n_323), .A2(n_749), .B(n_797), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_325), .A2(n_584), .B1(n_657), .B2(n_658), .Y(n_583) );
INVxp67_ASAP7_75t_SL g657 ( .A(n_325), .Y(n_657) );
CKINVDCx5p33_ASAP7_75t_R g1390 ( .A(n_326), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g1261 ( .A(n_327), .Y(n_1261) );
INVx1_ASAP7_75t_L g1391 ( .A(n_328), .Y(n_1391) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_329), .A2(n_350), .B1(n_1088), .B2(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g1461 ( .A(n_329), .Y(n_1461) );
OAI221xp5_ASAP7_75t_SL g982 ( .A1(n_330), .A2(n_361), .B1(n_559), .B2(n_983), .C(n_984), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_330), .A2(n_361), .B1(n_601), .B2(n_1013), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_331), .A2(n_351), .B1(n_1190), .B2(n_1458), .Y(n_1474) );
INVx1_ASAP7_75t_L g1491 ( .A(n_331), .Y(n_1491) );
INVx1_ASAP7_75t_L g1399 ( .A(n_332), .Y(n_1399) );
INVx1_ASAP7_75t_L g763 ( .A(n_333), .Y(n_763) );
CKINVDCx5p33_ASAP7_75t_R g1530 ( .A(n_335), .Y(n_1530) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_336), .Y(n_1380) );
INVx1_ASAP7_75t_L g864 ( .A(n_337), .Y(n_864) );
INVx1_ASAP7_75t_L g1436 ( .A(n_339), .Y(n_1436) );
CKINVDCx5p33_ASAP7_75t_R g1479 ( .A(n_341), .Y(n_1479) );
INVx1_ASAP7_75t_L g1546 ( .A(n_342), .Y(n_1546) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_343), .Y(n_693) );
INVx1_ASAP7_75t_L g1655 ( .A(n_344), .Y(n_1655) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_345), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_345), .B(n_380), .Y(n_1682) );
AND3x2_ASAP7_75t_L g1688 ( .A(n_345), .B(n_380), .C(n_1679), .Y(n_1688) );
CKINVDCx5p33_ASAP7_75t_R g1963 ( .A(n_346), .Y(n_1963) );
INVx2_ASAP7_75t_L g393 ( .A(n_347), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_348), .A2(n_365), .B1(n_1241), .B2(n_1320), .Y(n_1329) );
INVx1_ASAP7_75t_L g1348 ( .A(n_348), .Y(n_1348) );
INVx1_ASAP7_75t_L g1446 ( .A(n_350), .Y(n_1446) );
INVx1_ASAP7_75t_L g1495 ( .A(n_351), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g1968 ( .A(n_352), .Y(n_1968) );
INVx1_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
INVx2_ASAP7_75t_L g504 ( .A(n_354), .Y(n_504) );
OR2x2_ASAP7_75t_L g585 ( .A(n_355), .B(n_484), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g1967 ( .A(n_356), .Y(n_1967) );
INVx1_ASAP7_75t_L g1295 ( .A(n_357), .Y(n_1295) );
INVx1_ASAP7_75t_L g895 ( .A(n_358), .Y(n_895) );
INVx1_ASAP7_75t_L g458 ( .A(n_359), .Y(n_458) );
INVx1_ASAP7_75t_L g701 ( .A(n_360), .Y(n_701) );
INVx1_ASAP7_75t_L g1609 ( .A(n_362), .Y(n_1609) );
INVx1_ASAP7_75t_L g1355 ( .A(n_365), .Y(n_1355) );
INVx1_ASAP7_75t_L g1542 ( .A(n_366), .Y(n_1542) );
INVx1_ASAP7_75t_L g610 ( .A(n_367), .Y(n_610) );
AOI21xp33_ASAP7_75t_L g1376 ( .A1(n_368), .A2(n_460), .B(n_957), .Y(n_1376) );
INVx1_ASAP7_75t_L g1398 ( .A(n_368), .Y(n_1398) );
INVxp33_ASAP7_75t_SL g1209 ( .A(n_369), .Y(n_1209) );
INVx1_ASAP7_75t_L g1617 ( .A(n_370), .Y(n_1617) );
INVx1_ASAP7_75t_L g405 ( .A(n_372), .Y(n_405) );
INVx1_ASAP7_75t_L g1405 ( .A(n_373), .Y(n_1405) );
INVx1_ASAP7_75t_L g1170 ( .A(n_374), .Y(n_1170) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_396), .B(n_1667), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_383), .Y(n_377) );
AND2x4_ASAP7_75t_L g1952 ( .A(n_378), .B(n_384), .Y(n_1952) );
NOR2xp33_ASAP7_75t_SL g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_SL g1957 ( .A(n_379), .Y(n_1957) );
NAND2xp5_ASAP7_75t_L g2005 ( .A(n_379), .B(n_381), .Y(n_2005) );
HB1xp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g1956 ( .A(n_381), .B(n_1957), .Y(n_1956) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_389), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g622 ( .A(n_387), .B(n_395), .Y(n_622) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g540 ( .A(n_388), .B(n_541), .Y(n_540) );
OR2x6_ASAP7_75t_L g389 ( .A(n_390), .B(n_394), .Y(n_389) );
OR2x2_ASAP7_75t_L g485 ( .A(n_390), .B(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g544 ( .A(n_390), .Y(n_544) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_390), .Y(n_570) );
BUFx2_ASAP7_75t_L g871 ( .A(n_390), .Y(n_871) );
INVx1_ASAP7_75t_L g884 ( .A(n_390), .Y(n_884) );
OAI22xp33_ASAP7_75t_L g976 ( .A1(n_390), .A2(n_572), .B1(n_977), .B2(n_978), .Y(n_976) );
OAI22xp33_ASAP7_75t_L g991 ( .A1(n_390), .A2(n_572), .B1(n_992), .B2(n_993), .Y(n_991) );
INVx2_ASAP7_75t_SL g1158 ( .A(n_390), .Y(n_1158) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
AND2x4_ASAP7_75t_L g499 ( .A(n_392), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g509 ( .A(n_392), .Y(n_509) );
AND2x2_ASAP7_75t_L g515 ( .A(n_392), .B(n_393), .Y(n_515) );
INVx2_ASAP7_75t_L g520 ( .A(n_392), .Y(n_520) );
INVx1_ASAP7_75t_L g551 ( .A(n_392), .Y(n_551) );
INVx2_ASAP7_75t_L g500 ( .A(n_393), .Y(n_500) );
INVx1_ASAP7_75t_L g522 ( .A(n_393), .Y(n_522) );
INVx1_ASAP7_75t_L g529 ( .A(n_393), .Y(n_529) );
INVx1_ASAP7_75t_L g550 ( .A(n_393), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_393), .B(n_520), .Y(n_557) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_1078), .B1(n_1665), .B2(n_1666), .Y(n_396) );
INVx1_ASAP7_75t_SL g1666 ( .A(n_397), .Y(n_1666) );
XNOR2x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_818), .Y(n_397) );
XNOR2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_659), .Y(n_398) );
XOR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_583), .Y(n_399) );
INVx1_ASAP7_75t_L g581 ( .A(n_401), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_492), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_478), .B1(n_482), .B2(n_483), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_404), .B(n_421), .C(n_455), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_415), .B2(n_416), .Y(n_404) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_405), .A2(n_429), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_406), .A2(n_416), .B1(n_813), .B2(n_814), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_406), .A2(n_416), .B1(n_1072), .B2(n_1073), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1195 ( .A1(n_406), .A2(n_730), .B1(n_1167), .B2(n_1174), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1258 ( .A1(n_406), .A2(n_416), .B1(n_1226), .B2(n_1229), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_406), .A2(n_416), .B1(n_1312), .B2(n_1313), .Y(n_1311) );
AOI22xp33_ASAP7_75t_L g1331 ( .A1(n_406), .A2(n_416), .B1(n_1332), .B2(n_1333), .Y(n_1331) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_406), .A2(n_416), .B1(n_1387), .B2(n_1388), .Y(n_1386) );
AOI22xp33_ASAP7_75t_L g1459 ( .A1(n_406), .A2(n_416), .B1(n_1460), .B2(n_1461), .Y(n_1459) );
AOI22xp33_ASAP7_75t_L g1484 ( .A1(n_406), .A2(n_416), .B1(n_1485), .B2(n_1486), .Y(n_1484) );
AOI22xp33_ASAP7_75t_L g1517 ( .A1(n_406), .A2(n_416), .B1(n_1518), .B2(n_1519), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g1602 ( .A1(n_406), .A2(n_416), .B1(n_1603), .B2(n_1604), .Y(n_1602) );
AOI22xp33_ASAP7_75t_L g1920 ( .A1(n_406), .A2(n_416), .B1(n_1921), .B2(n_1922), .Y(n_1920) );
INVx6_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_410), .Y(n_407) );
OR2x2_ASAP7_75t_L g417 ( .A(n_408), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g428 ( .A(n_408), .Y(n_428) );
OR2x2_ASAP7_75t_L g908 ( .A(n_408), .B(n_502), .Y(n_908) );
INVx1_ASAP7_75t_L g453 ( .A(n_409), .Y(n_453) );
INVx2_ASAP7_75t_L g590 ( .A(n_410), .Y(n_590) );
INVx1_ASAP7_75t_L g949 ( .A(n_410), .Y(n_949) );
INVx1_ASAP7_75t_L g998 ( .A(n_410), .Y(n_998) );
BUFx2_ASAP7_75t_L g1592 ( .A(n_410), .Y(n_1592) );
OR2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
AND2x2_ASAP7_75t_L g599 ( .A(n_411), .B(n_413), .Y(n_599) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g419 ( .A(n_412), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AND2x4_ASAP7_75t_L g432 ( .A(n_414), .B(n_427), .Y(n_432) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_415), .A2(n_458), .B1(n_563), .B2(n_566), .Y(n_562) );
AOI211xp5_ASAP7_75t_L g1178 ( .A1(n_416), .A2(n_1170), .B(n_1179), .C(n_1181), .Y(n_1178) );
INVx4_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g951 ( .A(n_418), .Y(n_951) );
INVx2_ASAP7_75t_L g1243 ( .A(n_418), .Y(n_1243) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_419), .Y(n_449) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_419), .Y(n_593) );
INVx1_ASAP7_75t_L g811 ( .A(n_419), .Y(n_811) );
INVx1_ASAP7_75t_L g1185 ( .A(n_419), .Y(n_1185) );
AND2x2_ASAP7_75t_L g426 ( .A(n_420), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g447 ( .A(n_420), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_429), .B1(n_430), .B2(n_441), .C(n_450), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
BUFx6f_ASAP7_75t_L g711 ( .A(n_424), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_424), .A2(n_450), .B1(n_1327), .B2(n_1329), .C(n_1330), .Y(n_1326) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_424), .A2(n_450), .B1(n_1380), .B2(n_1381), .C(n_1385), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g1453 ( .A(n_424), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g1478 ( .A(n_424), .Y(n_1478) );
AOI221xp5_ASAP7_75t_L g1513 ( .A1(n_424), .A2(n_450), .B1(n_1514), .B2(n_1515), .C(n_1516), .Y(n_1513) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
AND2x4_ASAP7_75t_L g450 ( .A(n_425), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g721 ( .A(n_425), .Y(n_721) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_425), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_425), .A2(n_457), .B1(n_993), .B2(n_1000), .Y(n_999) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_425), .Y(n_1004) );
BUFx4f_ASAP7_75t_L g1382 ( .A(n_425), .Y(n_1382) );
INVx1_ASAP7_75t_L g1482 ( .A(n_425), .Y(n_1482) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_426), .Y(n_435) );
INVx2_ASAP7_75t_L g446 ( .A(n_427), .Y(n_446) );
AND2x2_ASAP7_75t_L g456 ( .A(n_428), .B(n_457), .Y(n_456) );
AND2x4_ASAP7_75t_L g730 ( .A(n_428), .B(n_613), .Y(n_730) );
AOI222xp33_ASAP7_75t_L g995 ( .A1(n_428), .A2(n_470), .B1(n_475), .B2(n_971), .C1(n_972), .C2(n_996), .Y(n_995) );
INVx2_ASAP7_75t_L g802 ( .A(n_431), .Y(n_802) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_432), .Y(n_457) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_432), .Y(n_465) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_432), .Y(n_601) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_432), .Y(n_613) );
INVx2_ASAP7_75t_SL g719 ( .A(n_432), .Y(n_719) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_432), .Y(n_740) );
BUFx2_ASAP7_75t_L g1190 ( .A(n_432), .Y(n_1190) );
BUFx3_ASAP7_75t_L g1240 ( .A(n_432), .Y(n_1240) );
BUFx2_ASAP7_75t_L g1328 ( .A(n_432), .Y(n_1328) );
INVx1_ASAP7_75t_L g1598 ( .A(n_433), .Y(n_1598) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g1254 ( .A(n_434), .Y(n_1254) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx6f_ASAP7_75t_L g727 ( .A(n_435), .Y(n_727) );
INVx1_ASAP7_75t_L g805 ( .A(n_435), .Y(n_805) );
BUFx6f_ASAP7_75t_L g1011 ( .A(n_435), .Y(n_1011) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g1005 ( .A(n_437), .Y(n_1005) );
INVx1_ASAP7_75t_L g1192 ( .A(n_437), .Y(n_1192) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_SL g602 ( .A(n_438), .Y(n_602) );
INVx2_ASAP7_75t_L g826 ( .A(n_438), .Y(n_826) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
AND2x4_ASAP7_75t_L g463 ( .A(n_439), .B(n_454), .Y(n_463) );
INVx2_ASAP7_75t_L g454 ( .A(n_440), .Y(n_454) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx4_ASAP7_75t_L g1194 ( .A(n_443), .Y(n_1194) );
INVx1_ASAP7_75t_L g1473 ( .A(n_443), .Y(n_1473) );
INVx1_ASAP7_75t_L g1910 ( .A(n_443), .Y(n_1910) );
BUFx6f_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g744 ( .A(n_444), .Y(n_744) );
INVx2_ASAP7_75t_SL g797 ( .A(n_444), .Y(n_797) );
INVx2_ASAP7_75t_L g808 ( .A(n_444), .Y(n_808) );
INVx1_ASAP7_75t_L g1320 ( .A(n_444), .Y(n_1320) );
INVx6_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g461 ( .A(n_445), .Y(n_461) );
AND2x2_ASAP7_75t_L g491 ( .A(n_445), .B(n_452), .Y(n_491) );
BUFx2_ASAP7_75t_L g1457 ( .A(n_445), .Y(n_1457) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g477 ( .A(n_446), .Y(n_477) );
INVx1_ASAP7_75t_L g473 ( .A(n_447), .Y(n_473) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g467 ( .A(n_449), .Y(n_467) );
BUFx6f_ASAP7_75t_L g716 ( .A(n_449), .Y(n_716) );
INVx2_ASAP7_75t_L g837 ( .A(n_449), .Y(n_837) );
BUFx6f_ASAP7_75t_L g1013 ( .A(n_449), .Y(n_1013) );
INVx1_ASAP7_75t_L g1127 ( .A(n_449), .Y(n_1127) );
INVx1_ASAP7_75t_L g603 ( .A(n_450), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g1001 ( .A1(n_450), .A2(n_1002), .B(n_1006), .Y(n_1001) );
AOI221xp5_ASAP7_75t_L g1452 ( .A1(n_450), .A2(n_1453), .B1(n_1454), .B2(n_1455), .C(n_1456), .Y(n_1452) );
AOI221xp5_ASAP7_75t_L g1477 ( .A1(n_450), .A2(n_1478), .B1(n_1479), .B2(n_1480), .C(n_1483), .Y(n_1477) );
BUFx3_ASAP7_75t_L g965 ( .A(n_451), .Y(n_965) );
BUFx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g470 ( .A(n_452), .B(n_471), .Y(n_470) );
AND2x4_ASAP7_75t_L g475 ( .A(n_452), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g726 ( .A(n_452), .Y(n_726) );
AND2x4_ASAP7_75t_L g732 ( .A(n_452), .B(n_471), .Y(n_732) );
AND2x2_ASAP7_75t_L g792 ( .A(n_452), .B(n_476), .Y(n_792) );
NAND2x1p5_ASAP7_75t_L g844 ( .A(n_452), .B(n_577), .Y(n_844) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_452), .B(n_476), .Y(n_1298) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_458), .B1(n_459), .B2(n_464), .C(n_468), .Y(n_455) );
INVx1_ASAP7_75t_L g605 ( .A(n_456), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g1318 ( .A1(n_456), .A2(n_1319), .B1(n_1322), .B2(n_1324), .C(n_1325), .Y(n_1318) );
BUFx4f_ASAP7_75t_L g1124 ( .A(n_457), .Y(n_1124) );
INVx1_ASAP7_75t_L g1301 ( .A(n_457), .Y(n_1301) );
INVx1_ASAP7_75t_L g1307 ( .A(n_457), .Y(n_1307) );
BUFx2_ASAP7_75t_L g830 ( .A(n_460), .Y(n_830) );
AND2x2_ASAP7_75t_L g906 ( .A(n_460), .B(n_907), .Y(n_906) );
A2O1A1Ixp33_ASAP7_75t_L g958 ( .A1(n_460), .A2(n_959), .B(n_960), .C(n_965), .Y(n_958) );
INVx2_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g1070 ( .A(n_461), .Y(n_1070) );
INVx1_ASAP7_75t_L g1187 ( .A(n_462), .Y(n_1187) );
INVx2_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g749 ( .A(n_463), .Y(n_749) );
AND2x4_ASAP7_75t_L g840 ( .A(n_463), .B(n_490), .Y(n_840) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_463), .Y(n_957) );
HB1xp67_ASAP7_75t_L g1061 ( .A(n_463), .Y(n_1061) );
OAI221xp5_ASAP7_75t_L g1244 ( .A1(n_463), .A2(n_1207), .B1(n_1245), .B2(n_1247), .C(n_1248), .Y(n_1244) );
INVx1_ASAP7_75t_L g1321 ( .A(n_463), .Y(n_1321) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g1008 ( .A(n_467), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1119 ( .A1(n_467), .A2(n_719), .B1(n_1104), .B2(n_1105), .Y(n_1119) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_470), .A2(n_475), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx2_ASAP7_75t_L g790 ( .A(n_470), .Y(n_790) );
INVx4_ASAP7_75t_L g1448 ( .A(n_470), .Y(n_1448) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_471), .A2(n_476), .B1(n_963), .B2(n_964), .Y(n_962) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g848 ( .A(n_472), .Y(n_848) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AOI322xp5_ASAP7_75t_L g1373 ( .A1(n_475), .A2(n_732), .A3(n_1374), .B1(n_1375), .B2(n_1376), .C1(n_1377), .C2(n_1378), .Y(n_1373) );
INVx2_ASAP7_75t_L g1476 ( .A(n_475), .Y(n_1476) );
INVx2_ASAP7_75t_L g736 ( .A(n_476), .Y(n_736) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g815 ( .A(n_478), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g1371 ( .A1(n_478), .A2(n_483), .B1(n_1372), .B2(n_1391), .Y(n_1371) );
CKINVDCx8_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g1084 ( .A1(n_479), .A2(n_1085), .B(n_1102), .Y(n_1084) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g618 ( .A(n_480), .Y(n_618) );
AND2x4_ASAP7_75t_L g621 ( .A(n_480), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g640 ( .A(n_480), .B(n_641), .Y(n_640) );
OR2x6_ASAP7_75t_L g825 ( .A(n_480), .B(n_826), .Y(n_825) );
AND2x4_ASAP7_75t_L g1039 ( .A(n_480), .B(n_622), .Y(n_1039) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OR2x6_ASAP7_75t_L g539 ( .A(n_481), .B(n_540), .Y(n_539) );
BUFx2_ASAP7_75t_L g904 ( .A(n_481), .Y(n_904) );
AOI22xp5_ASAP7_75t_L g1316 ( .A1(n_483), .A2(n_618), .B1(n_1317), .B2(n_1334), .Y(n_1316) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
INVx5_ASAP7_75t_L g663 ( .A(n_484), .Y(n_663) );
INVx2_ASAP7_75t_L g1463 ( .A(n_484), .Y(n_1463) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_488), .Y(n_484) );
INVx2_ASAP7_75t_L g980 ( .A(n_485), .Y(n_980) );
INVx3_ASAP7_75t_L g530 ( .A(n_486), .Y(n_530) );
INVx1_ASAP7_75t_L g893 ( .A(n_487), .Y(n_893) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI222xp33_ASAP7_75t_L g905 ( .A1(n_489), .A2(n_880), .B1(n_885), .B2(n_895), .C1(n_906), .C2(n_909), .Y(n_905) );
OR2x6_ASAP7_75t_L g1112 ( .A(n_489), .B(n_1113), .Y(n_1112) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g1015 ( .A(n_491), .Y(n_1015) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_523), .C(n_538), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_494), .B(n_510), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B1(n_505), .B2(n_506), .Y(n_494) );
INVx2_ASAP7_75t_L g655 ( .A(n_496), .Y(n_655) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .Y(n_496) );
INVx2_ASAP7_75t_L g631 ( .A(n_497), .Y(n_631) );
INVx1_ASAP7_75t_L g687 ( .A(n_497), .Y(n_687) );
INVx2_ASAP7_75t_L g990 ( .A(n_497), .Y(n_990) );
INVx2_ASAP7_75t_L g1354 ( .A(n_497), .Y(n_1354) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g560 ( .A(n_498), .Y(n_560) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_498), .Y(n_698) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g568 ( .A(n_499), .Y(n_568) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_499), .Y(n_777) );
AND2x4_ASAP7_75t_L g508 ( .A(n_500), .B(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g506 ( .A(n_501), .B(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g512 ( .A(n_501), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g517 ( .A(n_501), .B(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g652 ( .A(n_501), .B(n_518), .Y(n_652) );
AND2x4_ASAP7_75t_L g669 ( .A(n_501), .B(n_560), .Y(n_669) );
AND2x6_ASAP7_75t_L g671 ( .A(n_501), .B(n_537), .Y(n_671) );
AND2x2_ASAP7_75t_L g675 ( .A(n_501), .B(n_518), .Y(n_675) );
AND2x2_ASAP7_75t_L g923 ( .A(n_501), .B(n_894), .Y(n_923) );
AOI22xp5_ASAP7_75t_L g981 ( .A1(n_501), .A2(n_640), .B1(n_982), .B2(n_987), .Y(n_981) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_501), .B(n_518), .Y(n_1203) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_501), .B(n_518), .Y(n_1277) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
INVx2_ASAP7_75t_L g858 ( .A(n_503), .Y(n_858) );
AND2x4_ASAP7_75t_L g900 ( .A(n_503), .B(n_639), .Y(n_900) );
AND2x2_ASAP7_75t_L g902 ( .A(n_503), .B(n_519), .Y(n_902) );
INVx1_ASAP7_75t_L g541 ( .A(n_504), .Y(n_541) );
INVx1_ASAP7_75t_L g579 ( .A(n_504), .Y(n_579) );
INVx1_ASAP7_75t_L g656 ( .A(n_506), .Y(n_656) );
INVx2_ASAP7_75t_SL g783 ( .A(n_507), .Y(n_783) );
BUFx6f_ASAP7_75t_L g1425 ( .A(n_507), .Y(n_1425) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g537 ( .A(n_508), .Y(n_537) );
BUFx3_ASAP7_75t_L g626 ( .A(n_508), .Y(n_626) );
BUFx2_ASAP7_75t_L g649 ( .A(n_508), .Y(n_649) );
BUFx6f_ASAP7_75t_L g930 ( .A(n_508), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_516), .B2(n_517), .Y(n_510) );
AOI221xp5_ASAP7_75t_L g650 ( .A1(n_512), .A2(n_651), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_512), .A2(n_673), .B1(n_674), .B2(n_675), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_512), .A2(n_675), .B1(n_765), .B2(n_766), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_512), .A2(n_675), .B1(n_1034), .B2(n_1035), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_512), .A2(n_652), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
BUFx2_ASAP7_75t_L g1208 ( .A(n_512), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_512), .A2(n_1275), .B1(n_1276), .B2(n_1277), .Y(n_1274) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_512), .A2(n_675), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1397 ( .A1(n_512), .A2(n_517), .B1(n_1398), .B2(n_1399), .Y(n_1397) );
AOI22xp33_ASAP7_75t_L g1438 ( .A1(n_512), .A2(n_1203), .B1(n_1439), .B2(n_1440), .Y(n_1438) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_512), .A2(n_675), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g1536 ( .A1(n_512), .A2(n_652), .B1(n_1525), .B2(n_1537), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1930 ( .A1(n_512), .A2(n_1277), .B1(n_1931), .B2(n_1932), .Y(n_1930) );
BUFx2_ASAP7_75t_L g624 ( .A(n_513), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_513), .A2(n_649), .B1(n_985), .B2(n_986), .Y(n_984) );
BUFx3_ASAP7_75t_L g1041 ( .A(n_513), .Y(n_1041) );
INVx1_ASAP7_75t_L g1092 ( .A(n_513), .Y(n_1092) );
INVx1_ASAP7_75t_L g1433 ( .A(n_513), .Y(n_1433) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_SL g894 ( .A(n_514), .Y(n_894) );
INVx2_ASAP7_75t_L g1424 ( .A(n_514), .Y(n_1424) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_515), .Y(n_639) );
INVx1_ASAP7_75t_L g937 ( .A(n_517), .Y(n_937) );
INVx2_ASAP7_75t_SL g1287 ( .A(n_518), .Y(n_1287) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g629 ( .A(n_519), .Y(n_629) );
BUFx2_ASAP7_75t_L g774 ( .A(n_519), .Y(n_774) );
BUFx6f_ASAP7_75t_L g975 ( .A(n_519), .Y(n_975) );
BUFx6f_ASAP7_75t_L g988 ( .A(n_519), .Y(n_988) );
INVx1_ASAP7_75t_L g1089 ( .A(n_519), .Y(n_1089) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g534 ( .A(n_520), .Y(n_534) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_SL g1151 ( .A(n_525), .Y(n_1151) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g1344 ( .A(n_526), .Y(n_1344) );
NAND2x1_ASAP7_75t_SL g526 ( .A(n_527), .B(n_530), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_527), .A2(n_533), .B1(n_845), .B2(n_850), .Y(n_897) );
NAND2x1p5_ASAP7_75t_L g1096 ( .A(n_527), .B(n_1097), .Y(n_1096) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_529), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_530), .B(n_533), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_530), .B(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_L g643 ( .A(n_530), .B(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g645 ( .A(n_530), .B(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g648 ( .A(n_530), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_531), .Y(n_1212) );
BUFx4f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx4f_ASAP7_75t_L g677 ( .A(n_532), .Y(n_677) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OR2x6_ASAP7_75t_L g1098 ( .A(n_534), .B(n_892), .Y(n_1098) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g678 ( .A(n_536), .Y(n_678) );
BUFx2_ASAP7_75t_L g1539 ( .A(n_536), .Y(n_1539) );
BUFx2_ASAP7_75t_L g1984 ( .A(n_537), .Y(n_1984) );
OAI33xp33_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_542), .A3(n_553), .B1(n_562), .B2(n_569), .B3(n_574), .Y(n_538) );
OAI33xp33_ASAP7_75t_L g679 ( .A1(n_539), .A2(n_680), .A3(n_689), .B1(n_694), .B2(n_700), .B3(n_706), .Y(n_679) );
INVx1_ASAP7_75t_L g1154 ( .A(n_539), .Y(n_1154) );
HB1xp67_ASAP7_75t_L g1214 ( .A(n_539), .Y(n_1214) );
OAI33xp33_ASAP7_75t_L g1345 ( .A1(n_539), .A2(n_706), .A3(n_1346), .B1(n_1350), .B2(n_1356), .B3(n_1359), .Y(n_1345) );
OAI33xp33_ASAP7_75t_L g1401 ( .A1(n_539), .A2(n_706), .A3(n_1402), .B1(n_1406), .B2(n_1410), .B3(n_1413), .Y(n_1401) );
OAI33xp33_ASAP7_75t_L g1497 ( .A1(n_539), .A2(n_576), .A3(n_1498), .B1(n_1501), .B2(n_1505), .B3(n_1507), .Y(n_1497) );
OAI33xp33_ASAP7_75t_L g1540 ( .A1(n_539), .A2(n_706), .A3(n_1541), .B1(n_1545), .B2(n_1550), .B3(n_1551), .Y(n_1540) );
OAI22xp33_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .B1(n_546), .B2(n_552), .Y(n_542) );
BUFx2_ASAP7_75t_L g1947 ( .A(n_543), .Y(n_1947) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI22xp33_ASAP7_75t_L g1359 ( .A1(n_546), .A2(n_1330), .B1(n_1332), .B2(n_1347), .Y(n_1359) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_548), .B(n_892), .Y(n_1109) );
OAI22xp33_ASAP7_75t_L g1507 ( .A1(n_548), .A2(n_1347), .B1(n_1479), .B2(n_1485), .Y(n_1507) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx3_ASAP7_75t_L g704 ( .A(n_549), .Y(n_704) );
INVx2_ASAP7_75t_L g867 ( .A(n_549), .Y(n_867) );
BUFx2_ASAP7_75t_L g1412 ( .A(n_549), .Y(n_1412) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_550), .B(n_551), .Y(n_573) );
INVx1_ASAP7_75t_L g647 ( .A(n_551), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_558), .B1(n_559), .B2(n_561), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g862 ( .A1(n_554), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_862) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g876 ( .A(n_555), .Y(n_876) );
INVx2_ASAP7_75t_L g1942 ( .A(n_555), .Y(n_1942) );
BUFx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g983 ( .A(n_556), .Y(n_983) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g565 ( .A(n_557), .Y(n_565) );
BUFx2_ASAP7_75t_L g683 ( .A(n_557), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_559), .A2(n_563), .B1(n_1104), .B2(n_1105), .Y(n_1103) );
INVx1_ASAP7_75t_L g1430 ( .A(n_559), .Y(n_1430) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_SL g927 ( .A(n_560), .Y(n_927) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_560), .Y(n_1172) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g925 ( .A(n_565), .Y(n_925) );
INVx1_ASAP7_75t_L g1352 ( .A(n_565), .Y(n_1352) );
INVx2_ASAP7_75t_L g1980 ( .A(n_565), .Y(n_1980) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g1404 ( .A(n_567), .Y(n_1404) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_567), .Y(n_1428) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g635 ( .A(n_568), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_570), .A2(n_690), .B1(n_691), .B2(n_693), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_570), .A2(n_701), .B1(n_702), .B2(n_705), .Y(n_700) );
INVx1_ASAP7_75t_L g1553 ( .A(n_570), .Y(n_1553) );
OAI22xp33_ASAP7_75t_L g1155 ( .A1(n_571), .A2(n_1156), .B1(n_1157), .B2(n_1159), .Y(n_1155) );
OAI22xp33_ASAP7_75t_L g1173 ( .A1(n_571), .A2(n_1157), .B1(n_1174), .B2(n_1175), .Y(n_1173) );
OAI22xp33_ASAP7_75t_L g1946 ( .A1(n_571), .A2(n_1919), .B1(n_1921), .B2(n_1947), .Y(n_1946) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g692 ( .A(n_572), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g881 ( .A1(n_572), .A2(n_882), .B1(n_883), .B2(n_885), .C(n_886), .Y(n_881) );
INVx2_ASAP7_75t_L g1220 ( .A(n_572), .Y(n_1220) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI33xp33_ASAP7_75t_L g767 ( .A1(n_575), .A2(n_621), .A3(n_768), .B1(n_773), .B2(n_778), .B3(n_779), .Y(n_767) );
AOI33xp33_ASAP7_75t_L g1036 ( .A1(n_575), .A2(n_1037), .A3(n_1040), .B1(n_1042), .B2(n_1046), .B3(n_1047), .Y(n_1036) );
AOI33xp33_ASAP7_75t_L g1278 ( .A1(n_575), .A2(n_1279), .A3(n_1280), .B1(n_1284), .B2(n_1288), .B3(n_1290), .Y(n_1278) );
AOI33xp33_ASAP7_75t_L g1421 ( .A1(n_575), .A2(n_1422), .A3(n_1423), .B1(n_1426), .B2(n_1429), .B3(n_1431), .Y(n_1421) );
INVx6_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx5_ASAP7_75t_L g707 ( .A(n_576), .Y(n_707) );
OR2x6_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVx2_ASAP7_75t_L g641 ( .A(n_578), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g658 ( .A(n_584), .Y(n_658) );
NAND4xp75_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .C(n_619), .D(n_650), .Y(n_584) );
OAI31xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_604), .A3(n_615), .B(n_616), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B1(n_592), .B2(n_594), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_590), .Y(n_714) );
INVx2_ASAP7_75t_L g1060 ( .A(n_590), .Y(n_1060) );
INVx2_ASAP7_75t_L g1248 ( .A(n_590), .Y(n_1248) );
INVx1_ASAP7_75t_L g1662 ( .A(n_590), .Y(n_1662) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_593), .Y(n_1058) );
BUFx6f_ASAP7_75t_L g1323 ( .A(n_593), .Y(n_1323) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_600), .Y(n_595) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g611 ( .A(n_598), .Y(n_611) );
INVx2_ASAP7_75t_L g794 ( .A(n_598), .Y(n_794) );
BUFx4f_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g916 ( .A(n_599), .Y(n_916) );
INVx1_ASAP7_75t_L g954 ( .A(n_599), .Y(n_954) );
INVx1_ASAP7_75t_L g961 ( .A(n_599), .Y(n_961) );
BUFx2_ASAP7_75t_L g1246 ( .A(n_599), .Y(n_1246) );
INVx1_ASAP7_75t_L g1620 ( .A(n_599), .Y(n_1620) );
BUFx2_ASAP7_75t_L g828 ( .A(n_601), .Y(n_828) );
BUFx3_ASAP7_75t_L g835 ( .A(n_601), .Y(n_835) );
INVx1_ASAP7_75t_L g1057 ( .A(n_601), .Y(n_1057) );
INVx2_ASAP7_75t_L g1183 ( .A(n_601), .Y(n_1183) );
BUFx2_ASAP7_75t_L g722 ( .A(n_602), .Y(n_722) );
INVx1_ASAP7_75t_L g1068 ( .A(n_602), .Y(n_1068) );
INVx1_ASAP7_75t_L g1445 ( .A(n_605), .Y(n_1445) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_607), .A2(n_608), .B1(n_643), .B2(n_645), .C(n_648), .Y(n_642) );
OAI211xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_612), .C(n_614), .Y(n_609) );
INVx2_ASAP7_75t_SL g1624 ( .A(n_613), .Y(n_1624) );
OAI31xp33_ASAP7_75t_L g708 ( .A1(n_616), .A2(n_709), .A3(n_728), .B(n_750), .Y(n_708) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI31xp33_ASAP7_75t_SL g994 ( .A1(n_617), .A2(n_995), .A3(n_1001), .B(n_1009), .Y(n_994) );
OAI31xp33_ASAP7_75t_SL g1635 ( .A1(n_617), .A2(n_1636), .A3(n_1639), .B(n_1645), .Y(n_1635) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp67_ASAP7_75t_L g1113 ( .A(n_618), .B(n_890), .Y(n_1113) );
AND2x2_ASAP7_75t_SL g619 ( .A(n_620), .B(n_642), .Y(n_619) );
AOI33xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_623), .A3(n_627), .B1(n_632), .B2(n_636), .B3(n_640), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g973 ( .A1(n_621), .A2(n_974), .B1(n_979), .B2(n_980), .Y(n_973) );
BUFx2_ASAP7_75t_L g1422 ( .A(n_621), .Y(n_1422) );
INVx1_ASAP7_75t_L g874 ( .A(n_622), .Y(n_874) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x4_ASAP7_75t_L g860 ( .A(n_626), .B(n_857), .Y(n_860) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g1427 ( .A(n_629), .Y(n_1427) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g1358 ( .A(n_631), .Y(n_1358) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g856 ( .A(n_635), .B(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_SL g1285 ( .A(n_638), .Y(n_1285) );
INVx3_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_639), .Y(n_770) );
NAND3xp33_ASAP7_75t_L g931 ( .A(n_640), .B(n_932), .C(n_933), .Y(n_931) );
INVx2_ASAP7_75t_SL g887 ( .A(n_641), .Y(n_887) );
INVx1_ASAP7_75t_L g1651 ( .A(n_641), .Y(n_1651) );
AOI221xp5_ASAP7_75t_L g757 ( .A1(n_643), .A2(n_645), .B1(n_648), .B2(n_758), .C(n_759), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_643), .A2(n_645), .B1(n_648), .B2(n_971), .C(n_972), .Y(n_970) );
INVx1_ASAP7_75t_L g1027 ( .A(n_643), .Y(n_1027) );
AOI221xp5_ASAP7_75t_L g1418 ( .A1(n_643), .A2(n_645), .B1(n_648), .B2(n_1419), .C(n_1420), .Y(n_1418) );
AOI221xp5_ASAP7_75t_L g1560 ( .A1(n_643), .A2(n_645), .B1(n_648), .B2(n_1561), .C(n_1562), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1654 ( .A(n_644), .B(n_891), .Y(n_1654) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_645), .Y(n_1024) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_648), .A2(n_1024), .B1(n_1025), .B2(n_1026), .C(n_1028), .Y(n_1023) );
AOI221xp5_ASAP7_75t_L g1268 ( .A1(n_648), .A2(n_1024), .B1(n_1026), .B2(n_1269), .C(n_1270), .Y(n_1268) );
INVx1_ASAP7_75t_L g772 ( .A(n_649), .Y(n_772) );
HB1xp67_ASAP7_75t_L g1576 ( .A(n_649), .Y(n_1576) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_753), .B1(n_754), .B2(n_817), .Y(n_659) );
INVx1_ASAP7_75t_L g817 ( .A(n_660), .Y(n_817) );
INVx1_ASAP7_75t_L g751 ( .A(n_661), .Y(n_751) );
INVx1_ASAP7_75t_L g1262 ( .A(n_662), .Y(n_1262) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_663), .A2(n_785), .B(n_786), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g1048 ( .A1(n_663), .A2(n_1049), .B(n_1050), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_663), .A2(n_1075), .B1(n_1177), .B2(n_1196), .Y(n_1176) );
AOI21xp5_ASAP7_75t_L g1291 ( .A1(n_663), .A2(n_1292), .B(n_1293), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_663), .A2(n_1442), .B1(n_1512), .B2(n_1531), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1905 ( .A1(n_663), .A2(n_966), .B1(n_1906), .B2(n_1923), .Y(n_1905) );
NOR3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .C(n_679), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_672), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_670), .B2(n_671), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g738 ( .A1(n_667), .A2(n_674), .B1(n_715), .B2(n_739), .C(n_741), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g1435 ( .A1(n_668), .A2(n_671), .B1(n_1436), .B2(n_1437), .Y(n_1435) );
BUFx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g762 ( .A(n_669), .Y(n_762) );
BUFx2_ASAP7_75t_L g1031 ( .A(n_669), .Y(n_1031) );
BUFx2_ASAP7_75t_L g1145 ( .A(n_669), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_669), .A2(n_671), .B1(n_1338), .B2(n_1339), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1490 ( .A1(n_669), .A2(n_671), .B1(n_1491), .B2(n_1492), .Y(n_1490) );
BUFx2_ASAP7_75t_L g1569 ( .A(n_669), .Y(n_1569) );
BUFx2_ASAP7_75t_L g1928 ( .A(n_669), .Y(n_1928) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_671), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_671), .A2(n_1030), .B1(n_1031), .B2(n_1032), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_671), .A2(n_1144), .B1(n_1145), .B2(n_1146), .Y(n_1143) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_671), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g1271 ( .A1(n_671), .A2(n_1031), .B1(n_1272), .B2(n_1273), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1394 ( .A1(n_671), .A2(n_1145), .B1(n_1395), .B2(n_1396), .Y(n_1394) );
AOI22xp33_ASAP7_75t_L g1534 ( .A1(n_671), .A2(n_1031), .B1(n_1527), .B2(n_1535), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1926 ( .A1(n_671), .A2(n_1927), .B1(n_1928), .B2(n_1929), .Y(n_1926) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B1(n_685), .B2(n_688), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_681), .A2(n_695), .B1(n_696), .B2(n_699), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g1990 ( .A1(n_681), .A2(n_685), .B1(n_1991), .B2(n_1992), .Y(n_1990) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g1642 ( .A1(n_685), .A2(n_1223), .B1(n_1643), .B2(n_1644), .Y(n_1642) );
INVx2_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g712 ( .A1(n_688), .A2(n_690), .B1(n_713), .B2(n_715), .C(n_717), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g1228 ( .A1(n_691), .A2(n_1171), .B1(n_1229), .B2(n_1230), .Y(n_1228) );
BUFx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OAI22xp33_ASAP7_75t_L g1346 ( .A1(n_692), .A2(n_1347), .B1(n_1348), .B2(n_1349), .Y(n_1346) );
OAI22xp33_ASAP7_75t_L g1406 ( .A1(n_692), .A2(n_1407), .B1(n_1408), .B2(n_1409), .Y(n_1406) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g1165 ( .A(n_697), .Y(n_1165) );
INVx3_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g879 ( .A(n_698), .Y(n_879) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_704), .A2(n_892), .B(n_897), .Y(n_896) );
BUFx2_ASAP7_75t_L g1641 ( .A(n_704), .Y(n_1641) );
OAI33xp33_ASAP7_75t_L g1152 ( .A1(n_706), .A2(n_1153), .A3(n_1155), .B1(n_1160), .B2(n_1166), .B3(n_1173), .Y(n_1152) );
OAI33xp33_ASAP7_75t_L g1213 ( .A1(n_706), .A2(n_1214), .A3(n_1215), .B1(n_1221), .B2(n_1225), .B3(n_1228), .Y(n_1213) );
INVx1_ASAP7_75t_L g1579 ( .A(n_706), .Y(n_1579) );
OAI33xp33_ASAP7_75t_L g1934 ( .A1(n_706), .A2(n_1153), .A3(n_1935), .B1(n_1939), .B2(n_1945), .B3(n_1946), .Y(n_1934) );
CKINVDCx8_ASAP7_75t_R g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g1250 ( .A(n_710), .Y(n_1250) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_711), .A2(n_724), .B1(n_799), .B2(n_800), .C(n_806), .Y(n_798) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_711), .A2(n_724), .B1(n_1063), .B2(n_1064), .C(n_1069), .Y(n_1062) );
AOI221xp5_ASAP7_75t_L g1188 ( .A1(n_711), .A2(n_724), .B1(n_1175), .B2(n_1189), .C(n_1193), .Y(n_1188) );
AOI221xp5_ASAP7_75t_L g1303 ( .A1(n_711), .A2(n_724), .B1(n_1304), .B2(n_1305), .C(n_1309), .Y(n_1303) );
AOI221xp5_ASAP7_75t_L g1916 ( .A1(n_711), .A2(n_724), .B1(n_1917), .B2(n_1918), .C(n_1919), .Y(n_1916) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g913 ( .A(n_719), .Y(n_913) );
INVx2_ASAP7_75t_SL g1587 ( .A(n_719), .Y(n_1587) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g1257 ( .A(n_723), .Y(n_1257) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g1594 ( .A1(n_724), .A2(n_1478), .B1(n_1595), .B2(n_1596), .C(n_1599), .Y(n_1594) );
AND2x4_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g735 ( .A(n_726), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g832 ( .A(n_727), .Y(n_832) );
INVx1_ASAP7_75t_L g1117 ( .A(n_727), .Y(n_1117) );
BUFx6f_ASAP7_75t_L g1191 ( .A(n_727), .Y(n_1191) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_SL g787 ( .A1(n_730), .A2(n_788), .B(n_789), .Y(n_787) );
AOI211xp5_ASAP7_75t_L g1051 ( .A1(n_730), .A2(n_1052), .B(n_1053), .C(n_1055), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1234 ( .A(n_730), .Y(n_1234) );
AOI211xp5_ASAP7_75t_SL g1294 ( .A1(n_730), .A2(n_1295), .B(n_1296), .C(n_1299), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1389 ( .A(n_730), .B(n_1390), .Y(n_1389) );
AOI221xp5_ASAP7_75t_L g1470 ( .A1(n_730), .A2(n_1471), .B1(n_1472), .B2(n_1474), .C(n_1475), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1529 ( .A(n_730), .B(n_1530), .Y(n_1529) );
AOI211xp5_ASAP7_75t_L g1583 ( .A1(n_730), .A2(n_1584), .B(n_1585), .C(n_1586), .Y(n_1583) );
AOI221xp5_ASAP7_75t_L g1907 ( .A1(n_730), .A2(n_1908), .B1(n_1911), .B2(n_1914), .C(n_1915), .Y(n_1907) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_734), .B2(n_737), .Y(n_731) );
INVx2_ASAP7_75t_L g1054 ( .A(n_732), .Y(n_1054) );
INVx1_ASAP7_75t_L g1180 ( .A(n_732), .Y(n_1180) );
INVx2_ASAP7_75t_SL g1236 ( .A(n_732), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1520 ( .A1(n_732), .A2(n_1298), .B1(n_1521), .B2(n_1522), .Y(n_1520) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OR2x6_ASAP7_75t_L g843 ( .A(n_736), .B(n_844), .Y(n_843) );
OR2x2_ASAP7_75t_L g1131 ( .A(n_736), .B(n_844), .Y(n_1131) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
BUFx6f_ASAP7_75t_L g1007 ( .A(n_744), .Y(n_1007) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g1066 ( .A(n_747), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1132 ( .A(n_747), .B(n_852), .Y(n_1132) );
BUFx2_ASAP7_75t_SL g1308 ( .A(n_747), .Y(n_1308) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
XNOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_816), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_784), .Y(n_755) );
AND4x1_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .C(n_764), .D(n_767), .Y(n_756) );
OAI211xp5_ASAP7_75t_L g793 ( .A1(n_763), .A2(n_794), .B(n_795), .C(n_796), .Y(n_793) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g781 ( .A(n_770), .Y(n_781) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g1939 ( .A1(n_776), .A2(n_1940), .B1(n_1943), .B2(n_1944), .Y(n_1939) );
INVx2_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_SL g865 ( .A(n_777), .Y(n_865) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_777), .Y(n_1045) );
INVx4_ASAP7_75t_L g1282 ( .A(n_777), .Y(n_1282) );
BUFx3_ASAP7_75t_L g1289 ( .A(n_777), .Y(n_1289) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_783), .Y(n_1283) );
AOI31xp33_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_798), .A3(n_812), .B(n_815), .Y(n_786) );
INVx3_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
AND2x2_ASAP7_75t_L g851 ( .A(n_804), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g1909 ( .A(n_805), .Y(n_1909) );
BUFx3_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
HB1xp67_ASAP7_75t_L g1118 ( .A(n_808), .Y(n_1118) );
BUFx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OR2x6_ASAP7_75t_L g910 ( .A(n_811), .B(n_908), .Y(n_910) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_811), .B(n_908), .Y(n_1137) );
AO22x2_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_1020), .B1(n_1076), .B2(n_1077), .Y(n_818) );
INVx1_ASAP7_75t_L g1076 ( .A(n_819), .Y(n_1076) );
XNOR2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_917), .Y(n_819) );
NAND4xp75_ASAP7_75t_L g821 ( .A(n_822), .B(n_853), .C(n_905), .D(n_911), .Y(n_821) );
AND2x2_ASAP7_75t_SL g822 ( .A(n_823), .B(n_841), .Y(n_822) );
AOI33xp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_827), .A3(n_829), .B1(n_833), .B2(n_834), .B3(n_838), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g1120 ( .A(n_825), .Y(n_1120) );
INVx1_ASAP7_75t_L g1384 ( .A(n_826), .Y(n_1384) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g1614 ( .A1(n_839), .A2(n_1615), .B1(n_1616), .B2(n_1627), .Y(n_1614) );
OAI22xp5_ASAP7_75t_L g1965 ( .A1(n_839), .A2(n_1615), .B1(n_1966), .B2(n_1970), .Y(n_1965) );
INVx4_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_840), .A2(n_1115), .B1(n_1120), .B2(n_1121), .C(n_1128), .Y(n_1114) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_845), .B1(n_846), .B2(n_850), .C(n_851), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_SL g849 ( .A(n_844), .Y(n_849) );
INVx1_ASAP7_75t_L g852 ( .A(n_844), .Y(n_852) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx2_ASAP7_75t_L g1130 ( .A(n_847), .Y(n_1130) );
INVx2_ASAP7_75t_L g1976 ( .A(n_847), .Y(n_1976) );
NAND2x1p5_ASAP7_75t_L g847 ( .A(n_848), .B(n_849), .Y(n_847) );
BUFx2_ASAP7_75t_L g1633 ( .A(n_851), .Y(n_1633) );
OAI31xp33_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_861), .A3(n_898), .B(n_903), .Y(n_853) );
INVx3_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_856), .A2(n_902), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
INVx3_ASAP7_75t_L g1638 ( .A(n_856), .Y(n_1638) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx8_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_866), .B1(n_875), .B2(n_881), .C(n_888), .Y(n_861) );
OAI221xp5_ASAP7_75t_L g1646 ( .A1(n_865), .A2(n_1647), .B1(n_1648), .B2(n_1649), .C(n_1650), .Y(n_1646) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B1(n_869), .B2(n_872), .C(n_873), .Y(n_866) );
OAI21xp5_ASAP7_75t_SL g1106 ( .A1(n_867), .A2(n_1107), .B(n_1108), .Y(n_1106) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_SL g1347 ( .A(n_870), .Y(n_1347) );
INVx1_ASAP7_75t_L g1407 ( .A(n_870), .Y(n_1407) );
INVx2_ASAP7_75t_SL g870 ( .A(n_871), .Y(n_870) );
OAI221xp5_ASAP7_75t_L g1640 ( .A1(n_873), .A2(n_1157), .B1(n_1617), .B2(n_1621), .C(n_1641), .Y(n_1640) );
OAI221xp5_ASAP7_75t_L g1989 ( .A1(n_873), .A2(n_1157), .B1(n_1937), .B2(n_1967), .C(n_1968), .Y(n_1989) );
INVx2_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_877), .B1(n_878), .B2(n_880), .Y(n_875) );
BUFx2_ASAP7_75t_L g1223 ( .A(n_876), .Y(n_1223) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_877), .A2(n_882), .B1(n_912), .B2(n_914), .Y(n_911) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
OAI22xp33_ASAP7_75t_L g1935 ( .A1(n_883), .A2(n_1936), .B1(n_1937), .B2(n_1938), .Y(n_1935) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g1217 ( .A(n_884), .Y(n_1217) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_895), .B(n_896), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_891), .B(n_894), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g1097 ( .A(n_892), .Y(n_1097) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
CKINVDCx6p67_ASAP7_75t_R g899 ( .A(n_900), .Y(n_899) );
INVx3_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx3_ASAP7_75t_L g1637 ( .A(n_902), .Y(n_1637) );
INVx2_ASAP7_75t_L g966 ( .A(n_903), .Y(n_966) );
BUFx8_ASAP7_75t_SL g1260 ( .A(n_903), .Y(n_1260) );
AOI31xp33_ASAP7_75t_L g1582 ( .A1(n_903), .A2(n_1583), .A3(n_1594), .B(n_1602), .Y(n_1582) );
INVx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
BUFx2_ASAP7_75t_L g1075 ( .A(n_904), .Y(n_1075) );
AOI221xp5_ASAP7_75t_L g1133 ( .A1(n_906), .A2(n_912), .B1(n_1134), .B2(n_1135), .C(n_1136), .Y(n_1133) );
AND2x2_ASAP7_75t_L g912 ( .A(n_907), .B(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OR2x6_ASAP7_75t_L g915 ( .A(n_908), .B(n_916), .Y(n_915) );
OR2x2_ASAP7_75t_L g1661 ( .A(n_908), .B(n_1662), .Y(n_1661) );
OR2x2_ASAP7_75t_L g1663 ( .A(n_908), .B(n_1301), .Y(n_1663) );
CKINVDCx6p67_ASAP7_75t_R g909 ( .A(n_910), .Y(n_909) );
CKINVDCx6p67_ASAP7_75t_R g914 ( .A(n_915), .Y(n_914) );
OAI21xp33_ASAP7_75t_L g943 ( .A1(n_916), .A2(n_944), .B(n_945), .Y(n_943) );
OAI221xp5_ASAP7_75t_L g1059 ( .A1(n_916), .A2(n_1032), .B1(n_1034), .B2(n_1060), .C(n_1061), .Y(n_1059) );
INVx1_ASAP7_75t_L g1630 ( .A(n_916), .Y(n_1630) );
XNOR2xp5_ASAP7_75t_L g917 ( .A(n_918), .B(n_967), .Y(n_917) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_935), .C(n_939), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_934), .Y(n_920) );
INVx1_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B1(n_927), .B2(n_928), .C(n_929), .Y(n_924) );
INVx1_ASAP7_75t_L g1169 ( .A(n_925), .Y(n_1169) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_928), .A2(n_947), .B1(n_948), .B2(n_950), .Y(n_946) );
INVx2_ASAP7_75t_SL g1094 ( .A(n_930), .Y(n_1094) );
BUFx2_ASAP7_75t_L g1434 ( .A(n_930), .Y(n_1434) );
NOR2xp33_ASAP7_75t_SL g935 ( .A(n_936), .B(n_938), .Y(n_935) );
OAI31xp33_ASAP7_75t_SL g939 ( .A1(n_940), .A2(n_941), .A3(n_942), .B(n_966), .Y(n_939) );
OAI211xp5_ASAP7_75t_SL g942 ( .A1(n_943), .A2(n_946), .B(n_952), .C(n_958), .Y(n_942) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_948), .A2(n_954), .B1(n_1061), .B2(n_1273), .C(n_1275), .Y(n_1302) );
INVx2_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OAI211xp5_ASAP7_75t_L g952 ( .A1(n_953), .A2(n_954), .B(n_955), .C(n_956), .Y(n_952) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_954), .A2(n_1060), .B1(n_1146), .B2(n_1148), .C(n_1187), .Y(n_1186) );
OAI211xp5_ASAP7_75t_L g1449 ( .A1(n_954), .A2(n_1437), .B(n_1450), .C(n_1451), .Y(n_1449) );
NAND2xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_962), .Y(n_960) );
INVx1_ASAP7_75t_L g1591 ( .A(n_961), .Y(n_1591) );
NAND2xp5_ASAP7_75t_SL g967 ( .A(n_968), .B(n_1016), .Y(n_967) );
INVx1_ASAP7_75t_L g1018 ( .A(n_969), .Y(n_1018) );
NAND3xp33_ASAP7_75t_SL g969 ( .A(n_970), .B(n_973), .C(n_981), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g1009 ( .A1(n_979), .A2(n_1010), .B1(n_1012), .B2(n_1014), .Y(n_1009) );
INVx2_ASAP7_75t_L g1163 ( .A(n_983), .Y(n_1163) );
BUFx3_ASAP7_75t_L g1043 ( .A(n_988), .Y(n_1043) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1017 ( .A(n_994), .Y(n_1017) );
INVx2_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
HB1xp67_ASAP7_75t_L g1310 ( .A(n_1013), .Y(n_1310) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1013), .Y(n_1526) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1013), .Y(n_1626) );
INVx2_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
NAND3xp33_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1018), .C(n_1019), .Y(n_1016) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1020), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1048), .Y(n_1021) );
AND4x1_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1029), .C(n_1033), .D(n_1036), .Y(n_1022) );
INVx1_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
AOI33xp33_ASAP7_75t_L g1570 ( .A1(n_1037), .A2(n_1571), .A3(n_1575), .B1(n_1577), .B2(n_1578), .B3(n_1579), .Y(n_1570) );
INVx2_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
BUFx3_ASAP7_75t_L g1279 ( .A(n_1039), .Y(n_1279) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AOI31xp33_ASAP7_75t_L g1050 ( .A1(n_1051), .A2(n_1062), .A3(n_1071), .B(n_1074), .Y(n_1050) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
AOI31xp33_ASAP7_75t_L g1293 ( .A1(n_1074), .A2(n_1294), .A3(n_1303), .B(n_1311), .Y(n_1293) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1074), .Y(n_1442) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1078), .Y(n_1665) );
XNOR2xp5_ASAP7_75t_L g1078 ( .A(n_1079), .B(n_1364), .Y(n_1078) );
XOR2xp5_ASAP7_75t_L g1079 ( .A(n_1080), .B(n_1197), .Y(n_1079) );
HB1xp67_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
XNOR2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1138), .Y(n_1081) );
NAND4xp25_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1110), .C(n_1114), .D(n_1133), .Y(n_1083) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1090), .B(n_1095), .Y(n_1086) );
INVx2_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
CKINVDCx11_ASAP7_75t_R g1656 ( .A(n_1098), .Y(n_1656) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_1100), .A2(n_1101), .B1(n_1123), .B2(n_1125), .Y(n_1122) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1611 ( .A(n_1112), .B(n_1612), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1962 ( .A(n_1112), .B(n_1963), .Y(n_1962) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1117), .Y(n_1116) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1120), .Y(n_1615) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1127), .Y(n_1256) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
XNOR2x1_ASAP7_75t_SL g1138 ( .A(n_1139), .B(n_1140), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1176), .Y(n_1140) );
NOR3xp33_ASAP7_75t_SL g1141 ( .A(n_1142), .B(n_1150), .C(n_1152), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1147), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1210 ( .A(n_1145), .Y(n_1210) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
INVx3_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1162), .B1(n_1164), .B2(n_1165), .Y(n_1160) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1163), .Y(n_1502) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1163), .Y(n_1506) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1163), .Y(n_1647) );
OAI22xp5_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1168), .B1(n_1170), .B2(n_1171), .Y(n_1166) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1171), .A2(n_1222), .B1(n_1223), .B2(n_1224), .Y(n_1221) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1172), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g1574 ( .A(n_1172), .Y(n_1574) );
NAND3xp33_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1188), .C(n_1195), .Y(n_1177) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1185), .Y(n_1588) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1185), .Y(n_1601) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1190), .Y(n_1524) );
XNOR2x1_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1263), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1231), .Y(n_1199) );
NOR3xp33_ASAP7_75t_SL g1200 ( .A(n_1201), .B(n_1211), .C(n_1213), .Y(n_1200) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1563 ( .A1(n_1203), .A2(n_1205), .B1(n_1564), .B2(n_1565), .Y(n_1563) );
INVxp67_ASAP7_75t_SL g1204 ( .A(n_1205), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1208), .B1(n_1209), .B2(n_1210), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1566 ( .A1(n_1208), .A2(n_1567), .B1(n_1568), .B2(n_1569), .Y(n_1566) );
OAI22xp5_ASAP7_75t_SL g1215 ( .A1(n_1216), .A2(n_1217), .B1(n_1218), .B2(n_1219), .Y(n_1215) );
OAI22xp33_ASAP7_75t_L g1225 ( .A1(n_1217), .A2(n_1223), .B1(n_1226), .B2(n_1227), .Y(n_1225) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_1219), .A2(n_1347), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
OAI22xp33_ASAP7_75t_L g1551 ( .A1(n_1219), .A2(n_1514), .B1(n_1518), .B2(n_1552), .Y(n_1551) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
INVx1_ASAP7_75t_L g1937 ( .A(n_1220), .Y(n_1937) );
AOI211xp5_ASAP7_75t_L g1233 ( .A1(n_1227), .A2(n_1234), .B(n_1235), .C(n_1237), .Y(n_1233) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_1230), .A2(n_1250), .B1(n_1251), .B2(n_1255), .C(n_1257), .Y(n_1249) );
AOI22xp33_ASAP7_75t_SL g1231 ( .A1(n_1232), .A2(n_1259), .B1(n_1261), .B2(n_1262), .Y(n_1231) );
NAND3xp33_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1249), .C(n_1258), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
BUFx3_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx2_ASAP7_75t_SL g1241 ( .A(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1242), .Y(n_1458) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1243), .Y(n_1242) );
BUFx2_ASAP7_75t_L g1913 ( .A(n_1243), .Y(n_1913) );
INVx2_ASAP7_75t_SL g1245 ( .A(n_1246), .Y(n_1245) );
OAI221xp5_ASAP7_75t_L g1627 ( .A1(n_1248), .A2(n_1628), .B1(n_1629), .B2(n_1631), .C(n_1632), .Y(n_1627) );
OAI221xp5_ASAP7_75t_L g1966 ( .A1(n_1248), .A2(n_1618), .B1(n_1967), .B2(n_1968), .C(n_1969), .Y(n_1966) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_SL g1994 ( .A(n_1259), .Y(n_1994) );
INVx5_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
AO22x2_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1314), .B1(n_1362), .B2(n_1363), .Y(n_1263) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1264), .Y(n_1363) );
XNOR2x1_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1266), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1291), .Y(n_1266) );
AND4x1_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1271), .C(n_1274), .D(n_1278), .Y(n_1267) );
INVx2_ASAP7_75t_SL g1281 ( .A(n_1282), .Y(n_1281) );
OAI22xp5_ASAP7_75t_L g1945 ( .A1(n_1282), .A2(n_1914), .B1(n_1922), .B2(n_1940), .Y(n_1945) );
OAI221xp5_ASAP7_75t_L g1979 ( .A1(n_1282), .A2(n_1980), .B1(n_1981), .B2(n_1982), .C(n_1983), .Y(n_1979) );
INVx3_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
INVx2_ASAP7_75t_SL g1297 ( .A(n_1298), .Y(n_1297) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx3_ASAP7_75t_L g1362 ( .A(n_1314), .Y(n_1362) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1315), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1316), .B(n_1335), .Y(n_1315) );
NAND3xp33_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1326), .C(n_1331), .Y(n_1317) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1321), .Y(n_1593) );
OAI22xp5_ASAP7_75t_L g1356 ( .A1(n_1324), .A2(n_1333), .B1(n_1351), .B2(n_1357), .Y(n_1356) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1343), .C(n_1345), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1340), .Y(n_1336) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_1347), .A2(n_1380), .B1(n_1387), .B2(n_1411), .Y(n_1410) );
OAI22xp33_ASAP7_75t_L g1541 ( .A1(n_1347), .A2(n_1542), .B1(n_1543), .B2(n_1544), .Y(n_1541) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_1351), .A2(n_1353), .B1(n_1354), .B2(n_1355), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1351), .A2(n_1403), .B1(n_1404), .B2(n_1405), .Y(n_1402) );
OAI22xp5_ASAP7_75t_L g1413 ( .A1(n_1351), .A2(n_1388), .B1(n_1390), .B2(n_1414), .Y(n_1413) );
BUFx2_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx2_ASAP7_75t_SL g1548 ( .A(n_1354), .Y(n_1548) );
OAI22xp5_ASAP7_75t_L g1550 ( .A1(n_1354), .A2(n_1506), .B1(n_1519), .B2(n_1530), .Y(n_1550) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
AOI22xp33_ASAP7_75t_L g1364 ( .A1(n_1365), .A2(n_1366), .B1(n_1555), .B2(n_1664), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1366), .Y(n_1365) );
XNOR2x2_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1465), .Y(n_1366) );
XNOR2xp5_ASAP7_75t_L g1367 ( .A(n_1368), .B(n_1415), .Y(n_1367) );
XNOR2xp5_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1370), .Y(n_1368) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1392), .Y(n_1370) );
NAND4xp25_ASAP7_75t_L g1372 ( .A(n_1373), .B(n_1379), .C(n_1386), .D(n_1389), .Y(n_1372) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
NOR3xp33_ASAP7_75t_SL g1392 ( .A(n_1393), .B(n_1400), .C(n_1401), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1397), .Y(n_1393) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_1404), .A2(n_1502), .B1(n_1503), .B2(n_1504), .Y(n_1501) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1412), .Y(n_1543) );
OAI22xp5_ASAP7_75t_L g1505 ( .A1(n_1414), .A2(n_1471), .B1(n_1486), .B2(n_1506), .Y(n_1505) );
XNOR2x1_ASAP7_75t_L g1415 ( .A(n_1416), .B(n_1464), .Y(n_1415) );
NAND2x1_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1441), .Y(n_1416) );
AND4x1_ASAP7_75t_L g1417 ( .A(n_1418), .B(n_1421), .C(n_1435), .D(n_1438), .Y(n_1417) );
BUFx3_ASAP7_75t_L g1572 ( .A(n_1424), .Y(n_1572) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1433), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1443), .B1(n_1462), .B2(n_1463), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1468 ( .A1(n_1442), .A2(n_1463), .B1(n_1469), .B2(n_1487), .Y(n_1468) );
NAND3xp33_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1452), .C(n_1459), .Y(n_1443) );
AOI21xp5_ASAP7_75t_SL g1444 ( .A1(n_1445), .A2(n_1446), .B(n_1447), .Y(n_1444) );
HB1xp67_ASAP7_75t_L g1600 ( .A(n_1457), .Y(n_1600) );
AOI21xp5_ASAP7_75t_L g1580 ( .A1(n_1463), .A2(n_1581), .B(n_1582), .Y(n_1580) );
XNOR2xp5_ASAP7_75t_L g1465 ( .A(n_1466), .B(n_1509), .Y(n_1465) );
XOR2x2_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1508), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1488), .Y(n_1467) );
NAND3xp33_ASAP7_75t_L g1469 ( .A(n_1470), .B(n_1477), .C(n_1484), .Y(n_1469) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
NOR3xp33_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1496), .C(n_1497), .Y(n_1488) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1493), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1545 ( .A1(n_1502), .A2(n_1546), .B1(n_1547), .B2(n_1549), .Y(n_1545) );
OAI22xp33_ASAP7_75t_L g1708 ( .A1(n_1508), .A2(n_1709), .B1(n_1712), .B2(n_1713), .Y(n_1708) );
XNOR2x1_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1554), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1510 ( .A(n_1511), .B(n_1532), .Y(n_1510) );
NAND5xp2_ASAP7_75t_L g1512 ( .A(n_1513), .B(n_1517), .C(n_1520), .D(n_1523), .E(n_1529), .Y(n_1512) );
OAI221xp5_ASAP7_75t_SL g1523 ( .A1(n_1524), .A2(n_1525), .B1(n_1526), .B2(n_1527), .C(n_1528), .Y(n_1523) );
NOR3xp33_ASAP7_75t_L g1532 ( .A(n_1533), .B(n_1538), .C(n_1540), .Y(n_1532) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1534), .B(n_1536), .Y(n_1533) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
INVx1_ASAP7_75t_L g1664 ( .A(n_1555), .Y(n_1664) );
AOI22xp5_ASAP7_75t_L g1555 ( .A1(n_1556), .A2(n_1557), .B1(n_1606), .B2(n_1607), .Y(n_1555) );
INVx2_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
XOR2x2_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1605), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1559), .B(n_1580), .Y(n_1558) );
AND4x1_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1563), .C(n_1566), .D(n_1570), .Y(n_1559) );
OAI221xp5_ASAP7_75t_L g1589 ( .A1(n_1565), .A2(n_1567), .B1(n_1590), .B2(n_1592), .C(n_1593), .Y(n_1589) );
INVx1_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
OAI221xp5_ASAP7_75t_L g1616 ( .A1(n_1592), .A2(n_1617), .B1(n_1618), .B2(n_1621), .C(n_1622), .Y(n_1616) );
OAI221xp5_ASAP7_75t_L g1970 ( .A1(n_1592), .A2(n_1629), .B1(n_1971), .B2(n_1972), .C(n_1973), .Y(n_1970) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1598), .Y(n_1597) );
INVx1_ASAP7_75t_L g1606 ( .A(n_1607), .Y(n_1606) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
XNOR2xp5_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1610), .Y(n_1608) );
AND4x1_ASAP7_75t_L g1610 ( .A(n_1611), .B(n_1613), .C(n_1635), .D(n_1658), .Y(n_1610) );
NOR3xp33_ASAP7_75t_L g1613 ( .A(n_1614), .B(n_1633), .C(n_1634), .Y(n_1613) );
INVx2_ASAP7_75t_L g1618 ( .A(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1624), .Y(n_1623) );
INVx1_ASAP7_75t_L g1625 ( .A(n_1626), .Y(n_1625) );
INVx2_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
NOR3xp33_ASAP7_75t_SL g1964 ( .A(n_1633), .B(n_1965), .C(n_1974), .Y(n_1964) );
AOI22xp33_ASAP7_75t_L g1652 ( .A1(n_1653), .A2(n_1655), .B1(n_1656), .B2(n_1657), .Y(n_1652) );
AOI22xp33_ASAP7_75t_L g1985 ( .A1(n_1653), .A2(n_1656), .B1(n_1986), .B2(n_1987), .Y(n_1985) );
HB1xp67_ASAP7_75t_L g1653 ( .A(n_1654), .Y(n_1653) );
NOR2xp33_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1660), .Y(n_1658) );
OAI221xp5_ASAP7_75t_L g1667 ( .A1(n_1668), .A2(n_1900), .B1(n_1901), .B2(n_1948), .C(n_1953), .Y(n_1667) );
HB1xp67_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
NOR4xp25_ASAP7_75t_L g1669 ( .A(n_1670), .B(n_1764), .C(n_1850), .D(n_1877), .Y(n_1669) );
O2A1O1Ixp33_ASAP7_75t_L g1670 ( .A1(n_1671), .A2(n_1701), .B(n_1722), .C(n_1756), .Y(n_1670) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
OAI211xp5_ASAP7_75t_L g1848 ( .A1(n_1672), .A2(n_1743), .B(n_1780), .C(n_1849), .Y(n_1848) );
AOI21xp5_ASAP7_75t_L g1875 ( .A1(n_1672), .A2(n_1728), .B(n_1795), .Y(n_1875) );
NAND2xp5_ASAP7_75t_L g1880 ( .A(n_1672), .B(n_1881), .Y(n_1880) );
AND2x2_ASAP7_75t_L g1672 ( .A(n_1673), .B(n_1692), .Y(n_1672) );
CKINVDCx5p33_ASAP7_75t_R g1729 ( .A(n_1673), .Y(n_1729) );
NAND2xp5_ASAP7_75t_L g1788 ( .A(n_1673), .B(n_1698), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1809 ( .A(n_1673), .B(n_1732), .Y(n_1809) );
NOR2xp33_ASAP7_75t_L g1819 ( .A(n_1673), .B(n_1820), .Y(n_1819) );
OR2x2_ASAP7_75t_L g1823 ( .A(n_1673), .B(n_1824), .Y(n_1823) );
AND2x2_ASAP7_75t_L g1836 ( .A(n_1673), .B(n_1820), .Y(n_1836) );
NOR2xp33_ASAP7_75t_L g1846 ( .A(n_1673), .B(n_1782), .Y(n_1846) );
AND2x2_ASAP7_75t_L g1852 ( .A(n_1673), .B(n_1760), .Y(n_1852) );
AND2x2_ASAP7_75t_L g1858 ( .A(n_1673), .B(n_1792), .Y(n_1858) );
AND2x2_ASAP7_75t_L g1888 ( .A(n_1673), .B(n_1783), .Y(n_1888) );
AND2x4_ASAP7_75t_SL g1673 ( .A(n_1674), .B(n_1686), .Y(n_1673) );
AND2x4_ASAP7_75t_L g1675 ( .A(n_1676), .B(n_1681), .Y(n_1675) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
OR2x2_ASAP7_75t_L g1711 ( .A(n_1677), .B(n_1682), .Y(n_1711) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1680), .Y(n_1677) );
HB1xp67_ASAP7_75t_L g2003 ( .A(n_1678), .Y(n_2003) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1680), .Y(n_1690) );
AND2x4_ASAP7_75t_L g1683 ( .A(n_1681), .B(n_1684), .Y(n_1683) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
OR2x2_ASAP7_75t_L g1715 ( .A(n_1682), .B(n_1685), .Y(n_1715) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
AND2x2_ASAP7_75t_L g1687 ( .A(n_1688), .B(n_1689), .Y(n_1687) );
AND2x4_ASAP7_75t_L g1691 ( .A(n_1688), .B(n_1690), .Y(n_1691) );
AND2x4_ASAP7_75t_L g1705 ( .A(n_1688), .B(n_1689), .Y(n_1705) );
HB1xp67_ASAP7_75t_L g2004 ( .A(n_1689), .Y(n_2004) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
INVx2_ASAP7_75t_L g1707 ( .A(n_1691), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1753 ( .A(n_1692), .B(n_1729), .Y(n_1753) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1692), .Y(n_1808) );
AND2x2_ASAP7_75t_L g1833 ( .A(n_1692), .B(n_1809), .Y(n_1833) );
AOI22xp33_ASAP7_75t_L g1898 ( .A1(n_1692), .A2(n_1757), .B1(n_1816), .B2(n_1899), .Y(n_1898) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1697), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1760 ( .A(n_1693), .B(n_1698), .Y(n_1760) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1693), .Y(n_1820) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1694), .B(n_1741), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1694), .B(n_1698), .Y(n_1792) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1695), .B(n_1696), .Y(n_1694) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
INVxp67_ASAP7_75t_SL g1741 ( .A(n_1698), .Y(n_1741) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1698), .Y(n_1783) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1700), .Y(n_1698) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1701), .Y(n_1826) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_1702), .B(n_1716), .Y(n_1701) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1702), .Y(n_1767) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1703), .Y(n_1702) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1704), .Y(n_1900) );
BUFx3_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1705), .Y(n_1719) );
INVx1_ASAP7_75t_L g1706 ( .A(n_1707), .Y(n_1706) );
OAI22xp5_ASAP7_75t_SL g1718 ( .A1(n_1707), .A2(n_1719), .B1(n_1720), .B2(n_1721), .Y(n_1718) );
INVx2_ASAP7_75t_L g1734 ( .A(n_1707), .Y(n_1734) );
BUFx3_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
OAI22xp33_ASAP7_75t_L g1735 ( .A1(n_1710), .A2(n_1736), .B1(n_1737), .B2(n_1738), .Y(n_1735) );
BUFx6f_ASAP7_75t_L g1710 ( .A(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1713 ( .A(n_1714), .Y(n_1713) );
INVx1_ASAP7_75t_L g1714 ( .A(n_1715), .Y(n_1714) );
HB1xp67_ASAP7_75t_L g1738 ( .A(n_1715), .Y(n_1738) );
CKINVDCx6p67_ASAP7_75t_R g1776 ( .A(n_1716), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1790 ( .A(n_1716), .B(n_1786), .Y(n_1790) );
OR2x2_ASAP7_75t_L g1817 ( .A(n_1716), .B(n_1786), .Y(n_1817) );
AND2x2_ASAP7_75t_L g1840 ( .A(n_1716), .B(n_1746), .Y(n_1840) );
OR2x2_ASAP7_75t_L g1847 ( .A(n_1716), .B(n_1761), .Y(n_1847) );
OR2x6_ASAP7_75t_L g1716 ( .A(n_1717), .B(n_1718), .Y(n_1716) );
OR2x2_ASAP7_75t_L g1780 ( .A(n_1717), .B(n_1718), .Y(n_1780) );
OAI22xp5_ASAP7_75t_L g1722 ( .A1(n_1723), .A2(n_1742), .B1(n_1749), .B2(n_1754), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1723 ( .A(n_1724), .B(n_1728), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1825 ( .A(n_1724), .B(n_1732), .Y(n_1825) );
A2O1A1Ixp33_ASAP7_75t_L g1872 ( .A1(n_1724), .A2(n_1786), .B(n_1873), .C(n_1875), .Y(n_1872) );
INVx1_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1725), .Y(n_1744) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1725), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1725), .B(n_1745), .Y(n_1761) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1725), .B(n_1746), .Y(n_1763) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1725), .B(n_1776), .Y(n_1775) );
OAI321xp33_ASAP7_75t_L g1811 ( .A1(n_1725), .A2(n_1765), .A3(n_1812), .B1(n_1814), .B2(n_1815), .C(n_1821), .Y(n_1811) );
NAND3xp33_ASAP7_75t_L g1832 ( .A(n_1725), .B(n_1816), .C(n_1833), .Y(n_1832) );
AND2x2_ASAP7_75t_L g1725 ( .A(n_1726), .B(n_1727), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1728 ( .A(n_1729), .B(n_1730), .Y(n_1728) );
OR2x2_ASAP7_75t_L g1758 ( .A(n_1729), .B(n_1759), .Y(n_1758) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1729), .B(n_1771), .Y(n_1770) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1729), .B(n_1733), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1813 ( .A(n_1729), .B(n_1740), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1843 ( .A(n_1729), .B(n_1760), .Y(n_1843) );
AND2x2_ASAP7_75t_L g1866 ( .A(n_1729), .B(n_1792), .Y(n_1866) );
AND2x2_ASAP7_75t_L g1874 ( .A(n_1729), .B(n_1773), .Y(n_1874) );
NOR2xp33_ASAP7_75t_L g1730 ( .A(n_1731), .B(n_1739), .Y(n_1730) );
NAND2xp5_ASAP7_75t_L g1759 ( .A(n_1731), .B(n_1760), .Y(n_1759) );
NOR2x1p5_ASAP7_75t_L g1773 ( .A(n_1731), .B(n_1774), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1818 ( .A(n_1731), .B(n_1819), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1837 ( .A(n_1731), .B(n_1743), .Y(n_1837) );
HB1xp67_ASAP7_75t_L g1881 ( .A(n_1731), .Y(n_1881) );
INVx2_ASAP7_75t_SL g1731 ( .A(n_1732), .Y(n_1731) );
BUFx3_ASAP7_75t_L g1752 ( .A(n_1732), .Y(n_1752) );
BUFx2_ASAP7_75t_L g1772 ( .A(n_1732), .Y(n_1772) );
NOR2xp33_ASAP7_75t_L g1895 ( .A(n_1732), .B(n_1744), .Y(n_1895) );
INVx2_ASAP7_75t_SL g1732 ( .A(n_1733), .Y(n_1732) );
AND2x2_ASAP7_75t_L g1795 ( .A(n_1733), .B(n_1744), .Y(n_1795) );
OR2x2_ASAP7_75t_L g1771 ( .A(n_1739), .B(n_1772), .Y(n_1771) );
NOR2xp33_ASAP7_75t_L g1882 ( .A(n_1739), .B(n_1883), .Y(n_1882) );
INVx1_ASAP7_75t_L g1739 ( .A(n_1740), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1800 ( .A(n_1740), .B(n_1801), .Y(n_1800) );
AND2x2_ASAP7_75t_L g1831 ( .A(n_1740), .B(n_1809), .Y(n_1831) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
NAND2xp5_ASAP7_75t_SL g1891 ( .A(n_1743), .B(n_1776), .Y(n_1891) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1745), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1802 ( .A(n_1744), .B(n_1776), .Y(n_1802) );
AND2x2_ASAP7_75t_L g1810 ( .A(n_1744), .B(n_1746), .Y(n_1810) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
BUFx6f_ASAP7_75t_L g1755 ( .A(n_1746), .Y(n_1755) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1746), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1748), .Y(n_1746) );
INVxp67_ASAP7_75t_L g1854 ( .A(n_1749), .Y(n_1854) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1751), .Y(n_1749) );
INVx3_ASAP7_75t_L g1830 ( .A(n_1750), .Y(n_1830) );
AOI221xp5_ASAP7_75t_L g1863 ( .A1(n_1750), .A2(n_1765), .B1(n_1810), .B2(n_1864), .C(n_1867), .Y(n_1863) );
O2A1O1Ixp33_ASAP7_75t_L g1838 ( .A1(n_1751), .A2(n_1839), .B(n_1840), .C(n_1841), .Y(n_1838) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1752), .B(n_1753), .Y(n_1751) );
NAND2xp5_ASAP7_75t_L g1868 ( .A(n_1752), .B(n_1866), .Y(n_1868) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1752), .Y(n_1890) );
A2O1A1Ixp33_ASAP7_75t_L g1869 ( .A1(n_1754), .A2(n_1818), .B(n_1870), .C(n_1872), .Y(n_1869) );
CKINVDCx14_ASAP7_75t_R g1754 ( .A(n_1755), .Y(n_1754) );
AOI32xp33_ASAP7_75t_L g1859 ( .A1(n_1755), .A2(n_1759), .A3(n_1765), .B1(n_1860), .B2(n_1861), .Y(n_1859) );
OAI21xp5_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1761), .B(n_1762), .Y(n_1756) );
INVx2_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
INVx2_ASAP7_75t_L g1774 ( .A(n_1760), .Y(n_1774) );
INVx2_ASAP7_75t_L g1853 ( .A(n_1761), .Y(n_1853) );
AOI21xp33_ASAP7_75t_L g1896 ( .A1(n_1762), .A2(n_1799), .B(n_1897), .Y(n_1896) );
INVx1_ASAP7_75t_L g1762 ( .A(n_1763), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1763), .B(n_1772), .Y(n_1779) );
AOI21xp33_ASAP7_75t_L g1855 ( .A1(n_1763), .A2(n_1856), .B(n_1859), .Y(n_1855) );
OAI211xp5_ASAP7_75t_L g1764 ( .A1(n_1765), .A2(n_1768), .B(n_1797), .C(n_1838), .Y(n_1764) );
INVx3_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
AOI31xp33_ASAP7_75t_L g1877 ( .A1(n_1766), .A2(n_1878), .A3(n_1884), .B(n_1898), .Y(n_1877) );
INVx2_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
NAND2xp5_ASAP7_75t_L g1814 ( .A(n_1767), .B(n_1776), .Y(n_1814) );
NAND2xp5_ASAP7_75t_L g1862 ( .A(n_1767), .B(n_1786), .Y(n_1862) );
O2A1O1Ixp33_ASAP7_75t_L g1768 ( .A1(n_1769), .A2(n_1773), .B(n_1775), .C(n_1777), .Y(n_1768) );
INVx1_ASAP7_75t_L g1769 ( .A(n_1770), .Y(n_1769) );
NAND2xp5_ASAP7_75t_L g1864 ( .A(n_1771), .B(n_1865), .Y(n_1864) );
OR2x2_ASAP7_75t_L g1787 ( .A(n_1772), .B(n_1788), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_1772), .B(n_1792), .Y(n_1791) );
NAND2xp5_ASAP7_75t_L g1845 ( .A(n_1772), .B(n_1846), .Y(n_1845) );
INVx2_ASAP7_75t_L g1849 ( .A(n_1772), .Y(n_1849) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1773), .Y(n_1892) );
AOI221xp5_ASAP7_75t_L g1798 ( .A1(n_1775), .A2(n_1799), .B1(n_1802), .B2(n_1803), .C(n_1805), .Y(n_1798) );
CKINVDCx5p33_ASAP7_75t_R g1889 ( .A(n_1775), .Y(n_1889) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1776), .B(n_1786), .Y(n_1785) );
AOI31xp33_ASAP7_75t_L g1805 ( .A1(n_1776), .A2(n_1806), .A3(n_1809), .B(n_1810), .Y(n_1805) );
AND2x2_ASAP7_75t_L g1885 ( .A(n_1776), .B(n_1810), .Y(n_1885) );
OAI321xp33_ASAP7_75t_L g1777 ( .A1(n_1778), .A2(n_1780), .A3(n_1781), .B1(n_1784), .B2(n_1787), .C(n_1789), .Y(n_1777) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
NOR3xp33_ASAP7_75t_L g1793 ( .A(n_1780), .B(n_1794), .C(n_1796), .Y(n_1793) );
OAI211xp5_ASAP7_75t_L g1834 ( .A1(n_1780), .A2(n_1835), .B(n_1836), .C(n_1837), .Y(n_1834) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1783), .Y(n_1782) );
OAI221xp5_ASAP7_75t_SL g1841 ( .A1(n_1784), .A2(n_1803), .B1(n_1842), .B2(n_1847), .C(n_1848), .Y(n_1841) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
INVx1_ASAP7_75t_L g1894 ( .A(n_1788), .Y(n_1894) );
AOI21xp5_ASAP7_75t_L g1789 ( .A1(n_1790), .A2(n_1791), .B(n_1793), .Y(n_1789) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1790), .Y(n_1828) );
AOI211xp5_ASAP7_75t_L g1884 ( .A1(n_1791), .A2(n_1885), .B(n_1886), .C(n_1896), .Y(n_1884) );
INVx1_ASAP7_75t_L g1796 ( .A(n_1792), .Y(n_1796) );
OAI211xp5_ASAP7_75t_L g1821 ( .A1(n_1792), .A2(n_1822), .B(n_1825), .C(n_1826), .Y(n_1821) );
INVx1_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
OR2x2_ASAP7_75t_L g1803 ( .A(n_1796), .B(n_1804), .Y(n_1803) );
NAND2xp5_ASAP7_75t_L g1807 ( .A(n_1796), .B(n_1808), .Y(n_1807) );
NOR3xp33_ASAP7_75t_SL g1797 ( .A(n_1798), .B(n_1811), .C(n_1827), .Y(n_1797) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
AND2x2_ASAP7_75t_L g1839 ( .A(n_1800), .B(n_1830), .Y(n_1839) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1801), .Y(n_1804) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
AOI21xp5_ASAP7_75t_L g1878 ( .A1(n_1810), .A2(n_1879), .B(n_1882), .Y(n_1878) );
NAND2xp5_ASAP7_75t_L g1856 ( .A(n_1812), .B(n_1857), .Y(n_1856) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1814), .Y(n_1876) );
NAND2xp5_ASAP7_75t_L g1815 ( .A(n_1816), .B(n_1818), .Y(n_1815) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
HB1xp67_ASAP7_75t_L g1835 ( .A(n_1819), .Y(n_1835) );
INVx1_ASAP7_75t_L g1824 ( .A(n_1820), .Y(n_1824) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
OAI211xp5_ASAP7_75t_L g1827 ( .A1(n_1828), .A2(n_1829), .B(n_1832), .C(n_1834), .Y(n_1827) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1830), .B(n_1831), .Y(n_1829) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1830), .Y(n_1871) );
INVx1_ASAP7_75t_L g1897 ( .A(n_1833), .Y(n_1897) );
INVx1_ASAP7_75t_L g1883 ( .A(n_1837), .Y(n_1883) );
AOI21xp5_ASAP7_75t_L g1851 ( .A1(n_1839), .A2(n_1852), .B(n_1853), .Y(n_1851) );
NOR2xp33_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1844), .Y(n_1842) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1843), .Y(n_1860) );
INVx1_ASAP7_75t_L g1844 ( .A(n_1845), .Y(n_1844) );
INVx1_ASAP7_75t_L g1899 ( .A(n_1847), .Y(n_1899) );
AOI321xp33_ASAP7_75t_L g1850 ( .A1(n_1851), .A2(n_1854), .A3(n_1855), .B1(n_1863), .B2(n_1869), .C(n_1876), .Y(n_1850) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1862), .Y(n_1861) );
INVx1_ASAP7_75t_L g1865 ( .A(n_1866), .Y(n_1865) );
INVx1_ASAP7_75t_L g1867 ( .A(n_1868), .Y(n_1867) );
INVx1_ASAP7_75t_L g1870 ( .A(n_1871), .Y(n_1870) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1874), .Y(n_1873) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
OAI321xp33_ASAP7_75t_L g1886 ( .A1(n_1887), .A2(n_1889), .A3(n_1890), .B1(n_1891), .B2(n_1892), .C(n_1893), .Y(n_1886) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1888), .Y(n_1887) );
NAND2xp5_ASAP7_75t_L g1893 ( .A(n_1894), .B(n_1895), .Y(n_1893) );
INVx2_ASAP7_75t_L g1901 ( .A(n_1902), .Y(n_1901) );
XNOR2x1_ASAP7_75t_L g1902 ( .A(n_1903), .B(n_1904), .Y(n_1902) );
AND2x2_ASAP7_75t_L g1904 ( .A(n_1905), .B(n_1924), .Y(n_1904) );
NAND3xp33_ASAP7_75t_L g1906 ( .A(n_1907), .B(n_1916), .C(n_1920), .Y(n_1906) );
HB1xp67_ASAP7_75t_L g1912 ( .A(n_1913), .Y(n_1912) );
NOR3xp33_ASAP7_75t_SL g1924 ( .A(n_1925), .B(n_1933), .C(n_1934), .Y(n_1924) );
NAND2xp5_ASAP7_75t_L g1925 ( .A(n_1926), .B(n_1930), .Y(n_1925) );
INVx2_ASAP7_75t_L g1940 ( .A(n_1941), .Y(n_1940) );
INVx2_ASAP7_75t_L g1941 ( .A(n_1942), .Y(n_1941) );
CKINVDCx5p33_ASAP7_75t_R g1948 ( .A(n_1949), .Y(n_1948) );
BUFx2_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
INVx1_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
INVx1_ASAP7_75t_L g1951 ( .A(n_1952), .Y(n_1951) );
INVx1_ASAP7_75t_L g1954 ( .A(n_1955), .Y(n_1954) );
CKINVDCx5p33_ASAP7_75t_R g1955 ( .A(n_1956), .Y(n_1955) );
A2O1A1Ixp33_ASAP7_75t_L g2001 ( .A1(n_1957), .A2(n_2002), .B(n_2004), .C(n_2005), .Y(n_2001) );
INVxp33_ASAP7_75t_L g1958 ( .A(n_1959), .Y(n_1958) );
INVx1_ASAP7_75t_L g1999 ( .A(n_1960), .Y(n_1999) );
BUFx2_ASAP7_75t_SL g1960 ( .A(n_1961), .Y(n_1960) );
AND4x1_ASAP7_75t_L g1961 ( .A(n_1962), .B(n_1964), .C(n_1977), .D(n_1995), .Y(n_1961) );
INVx2_ASAP7_75t_L g1975 ( .A(n_1976), .Y(n_1975) );
OAI31xp33_ASAP7_75t_L g1977 ( .A1(n_1978), .A2(n_1988), .A3(n_1993), .B(n_1994), .Y(n_1977) );
NOR2xp33_ASAP7_75t_L g1995 ( .A(n_1996), .B(n_1997), .Y(n_1995) );
HB1xp67_ASAP7_75t_L g2000 ( .A(n_2001), .Y(n_2000) );
INVx1_ASAP7_75t_L g2002 ( .A(n_2003), .Y(n_2002) );
endmodule