module fake_netlist_1_5514_n_50 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_50);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_50;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_47;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_48;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_49;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
AND2x4_ASAP7_75t_L g16 ( .A(n_4), .B(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
NOR2xp33_ASAP7_75t_SL g18 ( .A(n_10), .B(n_6), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_9), .Y(n_20) );
OAI22x1_ASAP7_75t_R g21 ( .A1(n_11), .A2(n_1), .B1(n_5), .B2(n_8), .Y(n_21) );
BUFx12f_ASAP7_75t_L g22 ( .A(n_0), .Y(n_22) );
HB1xp67_ASAP7_75t_L g23 ( .A(n_15), .Y(n_23) );
AOI22xp5_ASAP7_75t_L g24 ( .A1(n_16), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_23), .B(n_2), .Y(n_25) );
OAI221xp5_ASAP7_75t_L g26 ( .A1(n_17), .A2(n_3), .B1(n_4), .B2(n_5), .C(n_7), .Y(n_26) );
NOR2xp33_ASAP7_75t_L g27 ( .A(n_19), .B(n_7), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_24), .B(n_16), .Y(n_28) );
OAI21x1_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_20), .B(n_19), .Y(n_29) );
O2A1O1Ixp33_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_17), .B(n_16), .C(n_18), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_16), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OR2x2_ASAP7_75t_SL g33 ( .A(n_32), .B(n_21), .Y(n_33) );
AND2x4_ASAP7_75t_L g34 ( .A(n_31), .B(n_28), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AND2x2_ASAP7_75t_L g37 ( .A(n_34), .B(n_28), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_35), .Y(n_38) );
OAI322xp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_30), .A3(n_27), .B1(n_31), .B2(n_33), .C1(n_20), .C2(n_21), .Y(n_39) );
AOI21xp33_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_30), .B(n_28), .Y(n_40) );
NAND4xp75_ASAP7_75t_L g41 ( .A(n_40), .B(n_33), .C(n_31), .D(n_20), .Y(n_41) );
AND2x2_ASAP7_75t_L g42 ( .A(n_38), .B(n_28), .Y(n_42) );
NAND3xp33_ASAP7_75t_L g43 ( .A(n_38), .B(n_32), .C(n_29), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
AOI22xp5_ASAP7_75t_L g45 ( .A1(n_41), .A2(n_22), .B1(n_39), .B2(n_29), .Y(n_45) );
OR2x2_ASAP7_75t_L g46 ( .A(n_43), .B(n_8), .Y(n_46) );
OAI22x1_ASAP7_75t_L g47 ( .A1(n_45), .A2(n_22), .B1(n_12), .B2(n_13), .Y(n_47) );
INVx2_ASAP7_75t_SL g48 ( .A(n_46), .Y(n_48) );
OAI21xp5_ASAP7_75t_SL g49 ( .A1(n_48), .A2(n_44), .B(n_22), .Y(n_49) );
AO21x2_ASAP7_75t_L g50 ( .A1(n_49), .A2(n_47), .B(n_48), .Y(n_50) );
endmodule