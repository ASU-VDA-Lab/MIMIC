module fake_jpeg_24605_n_67 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_66;

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_7),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_18),
.B(n_20),
.Y(n_29)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_1),
.C(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_11),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_8),
.B1(n_12),
.B2(n_21),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_40),
.B(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_19),
.B1(n_12),
.B2(n_8),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_23),
.C(n_18),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_29),
.A2(n_11),
.B1(n_15),
.B2(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_46),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_15),
.B(n_13),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_13),
.Y(n_46)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_16),
.CI(n_27),
.CON(n_47),
.SN(n_47)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_53),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_33),
.B1(n_36),
.B2(n_40),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.C(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_56),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_31),
.C(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_51),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_32),
.B2(n_6),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_55),
.B(n_49),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_4),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_63),
.B(n_4),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_4),
.Y(n_67)
);


endmodule