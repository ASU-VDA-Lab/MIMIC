module fake_jpeg_11599_n_557 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_557);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_557;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_54),
.B(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_56),
.Y(n_122)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_65),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_23),
.B(n_16),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_67),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_26),
.B(n_9),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_22),
.A2(n_32),
.B1(n_40),
.B2(n_30),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_76),
.A2(n_78),
.B1(n_25),
.B2(n_42),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_42),
.A2(n_25),
.B1(n_22),
.B2(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_80),
.B(n_101),
.Y(n_138)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_81),
.Y(n_163)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_82),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx12f_ASAP7_75t_SL g120 ( 
.A(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_24),
.Y(n_93)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_30),
.Y(n_98)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_98),
.Y(n_154)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_99),
.Y(n_171)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_15),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_107),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_31),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_38),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_49),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_108),
.B(n_119),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_64),
.A2(n_49),
.B1(n_47),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_112),
.A2(n_148),
.B1(n_19),
.B2(n_52),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_53),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_161),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_134),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_89),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_135),
.B(n_39),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_47),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_140),
.B(n_159),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_141),
.A2(n_146),
.B1(n_153),
.B2(n_21),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_58),
.A2(n_38),
.B(n_46),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_142),
.B(n_175),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_78),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_55),
.A2(n_31),
.B1(n_46),
.B2(n_35),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_84),
.B(n_18),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_107),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_63),
.A2(n_46),
.B1(n_51),
.B2(n_43),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_71),
.A2(n_46),
.B1(n_51),
.B2(n_34),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_156),
.B(n_169),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_83),
.A2(n_46),
.B1(n_51),
.B2(n_34),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_39),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_105),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_56),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_88),
.A2(n_33),
.B1(n_43),
.B2(n_35),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_94),
.B(n_25),
.Y(n_175)
);

AOI22x1_ASAP7_75t_SL g176 ( 
.A1(n_111),
.A2(n_97),
.B1(n_104),
.B2(n_77),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_176),
.A2(n_187),
.B1(n_192),
.B2(n_109),
.Y(n_250)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_60),
.B1(n_62),
.B2(n_98),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_179),
.Y(n_273)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_131),
.Y(n_180)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_181),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_183),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_184),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_175),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_185),
.B(n_191),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_136),
.A2(n_65),
.B1(n_102),
.B2(n_86),
.Y(n_187)
);

INVx13_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx4_ASAP7_75t_SL g261 ( 
.A(n_188),
.Y(n_261)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_189),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_190),
.B(n_226),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_115),
.Y(n_195)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_124),
.Y(n_197)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_68),
.A3(n_74),
.B1(n_73),
.B2(n_27),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_198),
.B(n_227),
.Y(n_283)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_199),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_156),
.A2(n_35),
.B1(n_27),
.B2(n_28),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_202),
.A2(n_212),
.B1(n_213),
.B2(n_216),
.Y(n_281)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_203),
.Y(n_245)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

BUFx8_ASAP7_75t_L g205 ( 
.A(n_120),
.Y(n_205)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_134),
.A2(n_107),
.B1(n_103),
.B2(n_43),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_206),
.Y(n_268)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_207),
.Y(n_290)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_34),
.B1(n_27),
.B2(n_28),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_209),
.A2(n_132),
.B1(n_167),
.B2(n_117),
.Y(n_255)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_138),
.A2(n_28),
.B1(n_33),
.B2(n_50),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_214),
.Y(n_262)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_215),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_121),
.A2(n_19),
.B1(n_52),
.B2(n_50),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_217),
.Y(n_272)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_218),
.Y(n_276)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_219),
.Y(n_278)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_125),
.B(n_103),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_222),
.A2(n_236),
.B(n_238),
.Y(n_277)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_154),
.Y(n_223)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_155),
.A2(n_33),
.B1(n_52),
.B2(n_50),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_224),
.A2(n_228),
.B1(n_109),
.B2(n_123),
.Y(n_285)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_160),
.Y(n_225)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_225),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_128),
.B(n_19),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_120),
.B(n_36),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_169),
.A2(n_21),
.B1(n_36),
.B2(n_39),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_145),
.Y(n_229)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_229),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_172),
.B(n_21),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_231),
.B(n_235),
.Y(n_296)
);

AO22x2_ASAP7_75t_L g232 ( 
.A1(n_149),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_145),
.B(n_130),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_110),
.Y(n_234)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_110),
.B(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_133),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_237),
.B(n_122),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_133),
.B(n_8),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_118),
.B(n_8),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_10),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_240),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_186),
.A2(n_216),
.B1(n_193),
.B2(n_192),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_244),
.A2(n_259),
.B1(n_187),
.B2(n_196),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_254),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_250),
.A2(n_255),
.B1(n_202),
.B2(n_177),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_252),
.B(n_182),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_186),
.A2(n_118),
.B1(n_117),
.B2(n_132),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_263),
.B(n_11),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_191),
.A2(n_174),
.B1(n_114),
.B2(n_158),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_193),
.B(n_167),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_286),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_209),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_L g323 ( 
.A1(n_270),
.A2(n_293),
.B(n_282),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_230),
.B(n_123),
.CI(n_174),
.CON(n_275),
.SN(n_275)
);

OAI32xp33_ASAP7_75t_L g341 ( 
.A1(n_275),
.A2(n_10),
.A3(n_13),
.B1(n_12),
.B2(n_5),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_285),
.A2(n_297),
.B(n_39),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_198),
.B(n_158),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_157),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_295),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_188),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_232),
.B(n_157),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_228),
.A2(n_163),
.B1(n_123),
.B2(n_162),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_298),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_196),
.C(n_206),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_300),
.B(n_303),
.C(n_339),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g365 ( 
.A1(n_301),
.A2(n_349),
.B1(n_279),
.B2(n_290),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_284),
.C(n_274),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_305),
.Y(n_386)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_307),
.B(n_312),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_309),
.A2(n_328),
.B1(n_331),
.B2(n_340),
.Y(n_359)
);

BUFx12f_ASAP7_75t_L g310 ( 
.A(n_293),
.Y(n_310)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_310),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_256),
.A2(n_176),
.B1(n_177),
.B2(n_205),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_311),
.A2(n_348),
.B1(n_255),
.B2(n_290),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_261),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_272),
.Y(n_313)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_313),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_232),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_315),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_267),
.B(n_232),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_317),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_298),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_320),
.B(n_332),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_296),
.A2(n_205),
.B(n_180),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_249),
.B(n_276),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_252),
.B(n_241),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_322),
.B(n_325),
.Y(n_373)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_323),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_218),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_342),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_261),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_256),
.A2(n_183),
.B1(n_220),
.B2(n_194),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_286),
.A2(n_207),
.B1(n_122),
.B2(n_189),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_210),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_330),
.B(n_341),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_204),
.B1(n_201),
.B2(n_181),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_242),
.Y(n_333)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_333),
.Y(n_375)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_334),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_241),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_335),
.B(n_337),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_281),
.A2(n_162),
.B1(n_219),
.B2(n_184),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_336),
.A2(n_246),
.B1(n_276),
.B2(n_253),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_248),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_338),
.A2(n_280),
.B(n_258),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_281),
.B(n_7),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_268),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_275),
.B(n_0),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_266),
.B(n_289),
.Y(n_343)
);

OAI21xp33_ASAP7_75t_L g369 ( 
.A1(n_343),
.A2(n_345),
.B(n_14),
.Y(n_369)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_243),
.Y(n_344)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_344),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_275),
.A2(n_5),
.B1(n_6),
.B2(n_11),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_242),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_243),
.B(n_0),
.C(n_1),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_245),
.C(n_251),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_270),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_297),
.Y(n_349)
);

NOR2x1_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_277),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_364),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_354),
.A2(n_358),
.B1(n_360),
.B2(n_365),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_330),
.Y(n_356)
);

XNOR2x1_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_368),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_314),
.A2(n_285),
.B1(n_266),
.B2(n_246),
.Y(n_360)
);

NAND2xp33_ASAP7_75t_SL g397 ( 
.A(n_361),
.B(n_321),
.Y(n_397)
);

O2A1O1Ixp33_ASAP7_75t_L g367 ( 
.A1(n_315),
.A2(n_280),
.B(n_253),
.C(n_278),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_367),
.A2(n_371),
.B(n_389),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_303),
.B(n_260),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_L g416 ( 
.A1(n_369),
.A2(n_14),
.B(n_1),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_302),
.A2(n_330),
.B(n_308),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_339),
.A2(n_291),
.B1(n_260),
.B2(n_289),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_372),
.A2(n_382),
.B1(n_388),
.B2(n_390),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_300),
.A2(n_326),
.B1(n_301),
.B2(n_336),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_376),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_308),
.B(n_262),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_313),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_324),
.A2(n_291),
.B1(n_278),
.B2(n_287),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_309),
.A2(n_262),
.B1(n_251),
.B2(n_245),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_331),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_318),
.Y(n_409)
);

OAI22x1_ASAP7_75t_SL g388 ( 
.A1(n_328),
.A2(n_287),
.B1(n_271),
.B2(n_288),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_316),
.A2(n_288),
.B1(n_271),
.B2(n_273),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_378),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_392),
.Y(n_434)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_357),
.A2(n_304),
.A3(n_341),
.B1(n_319),
.B2(n_345),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_393),
.Y(n_445)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_353),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_395),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_370),
.A2(n_326),
.B(n_338),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_396),
.A2(n_397),
.B(n_381),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_376),
.A2(n_317),
.B1(n_319),
.B2(n_335),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_398),
.A2(n_412),
.B1(n_420),
.B2(n_424),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_310),
.Y(n_399)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_399),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_332),
.C(n_344),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_405),
.C(n_409),
.Y(n_427)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_415),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_382),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_403),
.B(n_423),
.Y(n_435)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_404),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_355),
.B(n_305),
.C(n_334),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_352),
.B(n_310),
.Y(n_408)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_408),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_310),
.Y(n_410)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_410),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_361),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_357),
.B(n_320),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_414),
.Y(n_448)
);

AOI222xp33_ASAP7_75t_L g415 ( 
.A1(n_371),
.A2(n_340),
.B1(n_347),
.B2(n_333),
.C1(n_273),
.C2(n_248),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_416),
.A2(n_370),
.B1(n_381),
.B2(n_372),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_418),
.Y(n_444)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_354),
.A2(n_306),
.B1(n_329),
.B2(n_299),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_356),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_426),
.C(n_405),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_390),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_422),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_364),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_360),
.A2(n_299),
.B1(n_258),
.B2(n_2),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_350),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_425),
.B(n_386),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_363),
.B(n_351),
.Y(n_426)
);

MAJx2_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_427),
.C(n_433),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_401),
.A2(n_422),
.B1(n_407),
.B2(n_414),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_417),
.B1(n_420),
.B2(n_424),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_411),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_431),
.B(n_440),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_385),
.C(n_363),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_433),
.B(n_441),
.C(n_447),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_391),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_391),
.C(n_387),
.Y(n_441)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_384),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_402),
.B(n_389),
.C(n_383),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_450),
.C(n_452),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_383),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_451),
.A2(n_396),
.B(n_401),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_398),
.B(n_379),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_399),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_439),
.Y(n_457)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_457),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_395),
.Y(n_459)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_459),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_440),
.B(n_413),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_460),
.B(n_467),
.Y(n_500)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_439),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_464),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_435),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_463),
.B(n_445),
.Y(n_489)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_443),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_471),
.C(n_473),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_407),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_447),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_469),
.A2(n_453),
.B(n_437),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_445),
.A2(n_394),
.B1(n_406),
.B2(n_415),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_470),
.A2(n_472),
.B1(n_477),
.B2(n_480),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_427),
.B(n_408),
.C(n_392),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_431),
.B(n_362),
.C(n_419),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_443),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_476),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_434),
.A2(n_425),
.B1(n_404),
.B2(n_358),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_430),
.A2(n_359),
.B1(n_388),
.B2(n_367),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_436),
.A2(n_393),
.B1(n_379),
.B2(n_418),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_481),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_430),
.A2(n_374),
.B1(n_375),
.B2(n_380),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_432),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_441),
.C(n_449),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_483),
.B(n_487),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_484),
.B(n_485),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_461),
.B(n_456),
.Y(n_485)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_458),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_456),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_488),
.B(n_500),
.Y(n_515)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_450),
.C(n_452),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_498),
.C(n_501),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_471),
.B(n_432),
.Y(n_491)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_491),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_459),
.B(n_446),
.Y(n_493)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_469),
.A2(n_451),
.B(n_454),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_496),
.A2(n_486),
.B(n_495),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_455),
.C(n_429),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_455),
.C(n_446),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_502),
.A2(n_475),
.B(n_479),
.Y(n_510)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_503),
.B(n_511),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_468),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_506),
.B(n_484),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_496),
.A2(n_475),
.B(n_479),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_509),
.A2(n_510),
.B(n_517),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_501),
.Y(n_511)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_492),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_514),
.B(n_444),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_497),
.A2(n_470),
.B1(n_472),
.B2(n_468),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_486),
.B1(n_502),
.B2(n_483),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_482),
.B(n_460),
.C(n_480),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_518),
.B(n_519),
.C(n_485),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_444),
.C(n_477),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_513),
.B(n_490),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_526),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_521),
.B(n_525),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_524),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_504),
.A2(n_494),
.B1(n_457),
.B2(n_497),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_503),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_500),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_527),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_532),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_488),
.C(n_375),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_519),
.C(n_513),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_508),
.A2(n_374),
.B1(n_380),
.B2(n_0),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_509),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_1),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g536 ( 
.A1(n_531),
.A2(n_512),
.B(n_507),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_536),
.A2(n_537),
.B(n_528),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_SL g539 ( 
.A(n_531),
.B(n_517),
.C(n_510),
.Y(n_539)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_539),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_540),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_539),
.A2(n_523),
.B(n_526),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_544),
.A2(n_547),
.B(n_535),
.Y(n_548)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_534),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_545),
.B(n_546),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_541),
.A2(n_516),
.B1(n_523),
.B2(n_505),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_548),
.B(n_550),
.Y(n_551)
);

A2O1A1Ixp33_ASAP7_75t_SL g550 ( 
.A1(n_542),
.A2(n_538),
.B(n_529),
.C(n_533),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_549),
.B(n_543),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_552),
.A2(n_544),
.B(n_537),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_553),
.A2(n_551),
.B(n_521),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_520),
.C(n_532),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_555),
.B(n_515),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_556),
.B(n_515),
.Y(n_557)
);


endmodule