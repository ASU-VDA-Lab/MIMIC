module fake_jpeg_31842_n_153 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_7),
.B(n_27),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

BUFx4f_ASAP7_75t_SL g61 ( 
.A(n_22),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_10),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_33),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_20),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_71),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_54),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_84),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_70),
.B1(n_75),
.B2(n_65),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_82),
.A2(n_60),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_69),
.B(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_49),
.Y(n_92)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_88),
.Y(n_91)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_96),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_61),
.B(n_53),
.C(n_58),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_64),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_98),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_63),
.B(n_59),
.C(n_50),
.D(n_65),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_79),
.A2(n_60),
.B1(n_23),
.B2(n_24),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_100),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_3),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_60),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_6),
.Y(n_120)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_6),
.Y(n_118)
);

NOR3xp33_ASAP7_75t_SL g112 ( 
.A(n_95),
.B(n_81),
.C(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_120),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_47),
.B(n_26),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_91),
.B(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_122),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_46),
.B(n_28),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_7),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_8),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_34),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_128),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_29),
.C(n_11),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_9),
.B1(n_14),
.B2(n_15),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_133),
.B1(n_35),
.B2(n_36),
.Y(n_142)
);

NAND2xp33_ASAP7_75t_SL g132 ( 
.A(n_119),
.B(n_108),
.Y(n_132)
);

AOI221xp5_ASAP7_75t_L g141 ( 
.A1(n_132),
.A2(n_114),
.B1(n_111),
.B2(n_109),
.C(n_108),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_115),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_25),
.C(n_30),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_134),
.A2(n_107),
.B1(n_114),
.B2(n_113),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_141),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_143),
.B1(n_45),
.B2(n_126),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_145),
.B(n_146),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_139),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_130),
.B(n_137),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_149),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

AOI31xp33_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_143),
.A3(n_135),
.B(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_140),
.Y(n_153)
);


endmodule