module fake_jpeg_2950_n_722 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_722);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_722;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_717;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_718;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_720;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_719;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_553;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_721;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_0),
.C(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_65),
.B(n_68),
.Y(n_153)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_66),
.Y(n_171)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_67),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_37),
.B(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_70),
.B(n_84),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_74),
.Y(n_149)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_78),
.B(n_111),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_81),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_83),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_8),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_85),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_86),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_87),
.B(n_100),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_89),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_91),
.Y(n_202)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_92),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_93),
.Y(n_187)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_94),
.Y(n_205)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_96),
.Y(n_220)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_97),
.Y(n_164)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx11_ASAP7_75t_L g211 ( 
.A(n_98),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_99),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_21),
.B(n_8),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_107),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_28),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_108),
.B(n_19),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_109),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_23),
.Y(n_110)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_36),
.B(n_10),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_33),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_114),
.Y(n_212)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_33),
.Y(n_116)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_116),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_117),
.Y(n_216)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_45),
.Y(n_118)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_118),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_43),
.Y(n_120)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_121),
.Y(n_208)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_48),
.Y(n_122)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_45),
.Y(n_123)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_20),
.Y(n_124)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_125),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g126 ( 
.A(n_30),
.Y(n_126)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_45),
.Y(n_128)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_23),
.Y(n_129)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_129),
.Y(n_186)
);

BUFx12_ASAP7_75t_L g130 ( 
.A(n_30),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g197 ( 
.A(n_130),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g132 ( 
.A(n_27),
.Y(n_132)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_40),
.Y(n_133)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_134),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_61),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_135),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_84),
.A2(n_40),
.B1(n_60),
.B2(n_59),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_136),
.A2(n_155),
.B1(n_6),
.B2(n_11),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_143),
.B(n_192),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_68),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_145),
.B(n_213),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_109),
.A2(n_40),
.B1(n_30),
.B2(n_46),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_32),
.B1(n_61),
.B2(n_57),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g242 ( 
.A1(n_157),
.A2(n_225),
.B1(n_126),
.B2(n_41),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_74),
.A2(n_40),
.B1(n_32),
.B2(n_53),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_162),
.A2(n_166),
.B1(n_218),
.B2(n_42),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_87),
.A2(n_31),
.B1(n_59),
.B2(n_58),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_100),
.B(n_57),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_168),
.B(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_108),
.B(n_56),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_180),
.B(n_196),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_107),
.B(n_105),
.C(n_119),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_183),
.B(n_10),
.C(n_2),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_118),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_65),
.B(n_56),
.Y(n_196)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_76),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_204),
.Y(n_283)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_123),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_117),
.A2(n_32),
.B1(n_53),
.B2(n_46),
.Y(n_218)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_69),
.Y(n_222)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_128),
.B(n_60),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_224),
.B(n_226),
.Y(n_268)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_72),
.A2(n_41),
.B1(n_27),
.B2(n_50),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_97),
.B(n_58),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_102),
.Y(n_227)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_82),
.B(n_31),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_228),
.B(n_17),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_167),
.A2(n_38),
.B1(n_28),
.B2(n_42),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_231),
.A2(n_247),
.B1(n_273),
.B2(n_284),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_135),
.B(n_89),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_232),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_167),
.B(n_86),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_233),
.B(n_240),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_153),
.A2(n_83),
.B1(n_90),
.B2(n_99),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_234),
.A2(n_217),
.B1(n_191),
.B2(n_144),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_93),
.B1(n_44),
.B2(n_55),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_235),
.A2(n_238),
.B1(n_278),
.B2(n_309),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_149),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_236),
.Y(n_360)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_237),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_153),
.A2(n_44),
.B1(n_55),
.B2(n_50),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_142),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_239),
.B(n_250),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_193),
.B(n_38),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_241),
.B(n_242),
.Y(n_323)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_243),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_244),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_137),
.B(n_130),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_245),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_41),
.B1(n_27),
.B2(n_126),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_249),
.B(n_269),
.Y(n_338)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_160),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_251),
.B(n_253),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_197),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_254),
.Y(n_357)
);

NAND2x2_ASAP7_75t_SL g256 ( 
.A(n_225),
.B(n_0),
.Y(n_256)
);

NAND2x1_ASAP7_75t_SL g355 ( 
.A(n_256),
.B(n_141),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_258),
.B(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_177),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_260),
.B(n_275),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_150),
.Y(n_261)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_194),
.B(n_7),
.C(n_2),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_205),
.C(n_202),
.Y(n_315)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_139),
.Y(n_264)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_264),
.Y(n_364)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_159),
.Y(n_265)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_155),
.A2(n_0),
.B1(n_3),
.B2(n_5),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_267),
.A2(n_274),
.B1(n_279),
.B2(n_217),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_158),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

NAND2x1_ASAP7_75t_L g272 ( 
.A(n_168),
.B(n_3),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_272),
.B(n_157),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_225),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_169),
.A2(n_6),
.B(n_11),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_276),
.A2(n_162),
.B(n_218),
.Y(n_334)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_173),
.Y(n_277)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_277),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g278 ( 
.A1(n_181),
.A2(n_6),
.B1(n_11),
.B2(n_15),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_169),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_178),
.Y(n_280)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_280),
.Y(n_343)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_281),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g363 ( 
.A(n_282),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_199),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_207),
.Y(n_285)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_285),
.Y(n_372)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_198),
.Y(n_286)
);

CKINVDCx6p67_ASAP7_75t_R g326 ( 
.A(n_286),
.Y(n_326)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_201),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_287),
.B(n_289),
.Y(n_331)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_178),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_288),
.Y(n_368)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_164),
.Y(n_289)
);

BUFx16f_ASAP7_75t_L g290 ( 
.A(n_141),
.Y(n_290)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_290),
.Y(n_361)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_188),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_293),
.Y(n_337)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_147),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_184),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_295),
.B(n_298),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_179),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_297),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_220),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_199),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_300),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_174),
.B(n_19),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_179),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_301),
.B(n_302),
.Y(n_365)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_191),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_176),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_303),
.B(n_304),
.Y(n_366)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_189),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_305),
.B(n_306),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_180),
.B(n_17),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_202),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_308),
.B(n_310),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_216),
.A2(n_18),
.B1(n_19),
.B2(n_152),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_138),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_313),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_315),
.B(n_245),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_146),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_340),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_200),
.C(n_175),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_318),
.B(n_362),
.C(n_243),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_230),
.B(n_157),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_329),
.B(n_342),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_256),
.A2(n_205),
.B1(n_189),
.B2(n_170),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_334),
.A2(n_355),
.B(n_373),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_256),
.A2(n_161),
.B1(n_172),
.B2(n_140),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_335),
.A2(n_346),
.B1(n_350),
.B2(n_359),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_339),
.A2(n_354),
.B1(n_371),
.B2(n_247),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_300),
.B(n_165),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_266),
.B(n_186),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_257),
.A2(n_203),
.B1(n_156),
.B2(n_185),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_232),
.A2(n_182),
.B1(n_215),
.B2(n_154),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_272),
.B(n_144),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_367),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_240),
.B(n_165),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_353),
.B(n_283),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_245),
.B(n_248),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g419 ( 
.A(n_358),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_242),
.A2(n_211),
.B1(n_212),
.B2(n_223),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_276),
.B(n_229),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_151),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_242),
.A2(n_151),
.B1(n_187),
.B2(n_229),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_370),
.A2(n_252),
.B1(n_290),
.B2(n_305),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_273),
.A2(n_235),
.B1(n_241),
.B2(n_238),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_241),
.A2(n_187),
.B(n_231),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_263),
.A2(n_267),
.B1(n_294),
.B2(n_264),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_375),
.A2(n_290),
.B1(n_303),
.B2(n_255),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_376),
.A2(n_413),
.B1(n_416),
.B2(n_422),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_338),
.B(n_236),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_379),
.B(n_395),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_380),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_345),
.B(n_258),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_381),
.B(n_391),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_316),
.B(n_262),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_323),
.A2(n_371),
.B1(n_329),
.B2(n_348),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_384),
.A2(n_397),
.B1(n_421),
.B2(n_339),
.Y(n_453)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_386),
.Y(n_429)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_333),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

INVx6_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_390),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_345),
.B(n_265),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g392 ( 
.A(n_338),
.B(n_317),
.C(n_342),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_356),
.Y(n_394)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_321),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_246),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_323),
.A2(n_309),
.B1(n_291),
.B2(n_283),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_400),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_321),
.Y(n_401)
);

BUFx24_ASAP7_75t_SL g469 ( 
.A(n_401),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_320),
.B(n_297),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_402),
.Y(n_427)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_347),
.Y(n_403)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_403),
.Y(n_455)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_347),
.Y(n_404)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_404),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_407),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_336),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_337),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_410),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_330),
.B(n_282),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_409),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_330),
.B(n_293),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_417),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_373),
.A2(n_284),
.B1(n_280),
.B2(n_302),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_414),
.B(n_415),
.Y(n_466)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_255),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_331),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_418),
.B(n_420),
.Y(n_437)
);

OAI32xp33_ASAP7_75t_L g420 ( 
.A1(n_323),
.A2(n_259),
.A3(n_286),
.B1(n_288),
.B2(n_237),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_323),
.A2(n_259),
.B1(n_244),
.B2(n_261),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_313),
.A2(n_301),
.B1(n_296),
.B2(n_281),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_349),
.B(n_317),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_424),
.Y(n_438)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_336),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_313),
.A2(n_354),
.B1(n_334),
.B2(n_375),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_425),
.A2(n_411),
.B1(n_384),
.B2(n_417),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_325),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_365),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_382),
.A2(n_319),
.B(n_358),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_425),
.A2(n_348),
.B1(n_349),
.B2(n_351),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_434),
.A2(n_464),
.B1(n_389),
.B2(n_383),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_440),
.A2(n_434),
.B1(n_463),
.B2(n_464),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_382),
.A2(n_399),
.B(n_419),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_447),
.Y(n_478)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_448),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_385),
.B(n_367),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_453),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_399),
.A2(n_355),
.B(n_358),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_452),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_385),
.B(n_349),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_463),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_397),
.A2(n_355),
.B(n_358),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_458),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_377),
.A2(n_326),
.B(n_344),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_460),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_349),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_387),
.A2(n_322),
.B1(n_353),
.B2(n_315),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_418),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_467),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_387),
.A2(n_326),
.B(n_322),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_405),
.A2(n_326),
.B(n_344),
.Y(n_468)
);

OAI21xp33_ASAP7_75t_L g487 ( 
.A1(n_468),
.A2(n_381),
.B(n_379),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_470),
.B(n_501),
.Y(n_519)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_471),
.Y(n_513)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_461),
.Y(n_472)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_472),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_427),
.B(n_395),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_474),
.B(n_493),
.Y(n_512)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_461),
.Y(n_476)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_476),
.Y(n_518)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_477),
.Y(n_525)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_466),
.Y(n_480)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_480),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_434),
.A2(n_421),
.B1(n_403),
.B2(n_404),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_481),
.A2(n_484),
.B1(n_502),
.B2(n_432),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_482),
.A2(n_499),
.B1(n_507),
.B2(n_459),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_423),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_483),
.B(n_495),
.C(n_452),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_440),
.A2(n_420),
.B1(n_392),
.B2(n_386),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_442),
.B(n_410),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_496),
.Y(n_523)
);

OAI21xp33_ASAP7_75t_L g511 ( 
.A1(n_487),
.A2(n_468),
.B(n_444),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_449),
.B(n_324),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_488),
.B(n_491),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_449),
.B(n_324),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_442),
.B(n_318),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_492),
.B(n_464),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_427),
.B(n_391),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_466),
.Y(n_494)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_494),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_442),
.B(n_393),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_398),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_465),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_498),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_428),
.A2(n_394),
.B1(n_340),
.B2(n_390),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_433),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g502 ( 
.A1(n_437),
.A2(n_368),
.B1(n_365),
.B2(n_341),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_433),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_503),
.B(n_505),
.Y(n_527)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_429),
.Y(n_504)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_504),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_433),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_446),
.Y(n_506)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_506),
.Y(n_530)
);

CKINVDCx14_ASAP7_75t_R g507 ( 
.A(n_446),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_511),
.B(n_540),
.Y(n_553)
);

AOI21xp33_ASAP7_75t_L g514 ( 
.A1(n_508),
.A2(n_460),
.B(n_431),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_514),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_492),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_524),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_472),
.Y(n_516)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_516),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_475),
.A2(n_437),
.B1(n_428),
.B2(n_447),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_543),
.B1(n_504),
.B2(n_429),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_481),
.A2(n_453),
.B1(n_447),
.B2(n_450),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_521),
.A2(n_522),
.B1(n_526),
.B2(n_536),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_475),
.A2(n_467),
.B1(n_457),
.B2(n_458),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_470),
.B(n_457),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_502),
.A2(n_484),
.B1(n_498),
.B2(n_486),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_500),
.A2(n_456),
.B1(n_473),
.B2(n_486),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_529),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_490),
.B(n_455),
.Y(n_532)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_532),
.Y(n_549)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_490),
.Y(n_533)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_535),
.B(n_537),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_486),
.A2(n_467),
.B1(n_458),
.B2(n_455),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_430),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_538),
.B(n_432),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_430),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_539),
.B(n_495),
.C(n_462),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_497),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_473),
.A2(n_452),
.B(n_456),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_541),
.B(n_542),
.Y(n_560)
);

OAI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_478),
.A2(n_458),
.B(n_435),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_471),
.A2(n_454),
.B1(n_459),
.B2(n_438),
.Y(n_543)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_544),
.Y(n_565)
);

OAI21xp33_ASAP7_75t_L g545 ( 
.A1(n_497),
.A2(n_508),
.B(n_478),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_545),
.B(n_439),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_547),
.B(n_489),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_550),
.B(n_554),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g590 ( 
.A(n_552),
.B(n_557),
.Y(n_590)
);

AOI32xp33_ASAP7_75t_L g554 ( 
.A1(n_530),
.A2(n_479),
.A3(n_477),
.B1(n_480),
.B2(n_494),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_510),
.B(n_532),
.Y(n_555)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_515),
.B(n_523),
.C(n_535),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_556),
.B(n_558),
.C(n_561),
.Y(n_600)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_438),
.C(n_489),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_516),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_559),
.B(n_569),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_537),
.B(n_445),
.C(n_441),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_562),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_527),
.B(n_441),
.Y(n_564)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_527),
.B(n_436),
.Y(n_566)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_566),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_436),
.C(n_445),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_567),
.B(n_581),
.C(n_366),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_533),
.B(n_476),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g607 ( 
.A1(n_570),
.A2(n_326),
.B(n_451),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_512),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g584 ( 
.A(n_571),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_546),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_573),
.B(n_575),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_534),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_574),
.Y(n_588)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_530),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_576),
.B(n_577),
.Y(n_612)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_509),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_525),
.B(n_505),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_524),
.B(n_469),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_509),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_539),
.B(n_369),
.C(n_414),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_SL g585 ( 
.A(n_583),
.B(n_522),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_585),
.B(n_589),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_560),
.A2(n_542),
.B(n_536),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g617 ( 
.A1(n_586),
.A2(n_592),
.B1(n_593),
.B2(n_594),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_583),
.B(n_519),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_576),
.A2(n_547),
.B1(n_526),
.B2(n_521),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_591),
.A2(n_608),
.B1(n_563),
.B2(n_578),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_572),
.A2(n_519),
.B1(n_531),
.B2(n_528),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_572),
.A2(n_513),
.B1(n_541),
.B2(n_517),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_565),
.A2(n_573),
.B1(n_562),
.B2(n_549),
.Y(n_594)
);

FAx1_ASAP7_75t_SL g596 ( 
.A(n_551),
.B(n_558),
.CI(n_556),
.CON(n_596),
.SN(n_596)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_596),
.B(n_600),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_565),
.A2(n_518),
.B1(n_503),
.B2(n_501),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g630 ( 
.A1(n_598),
.A2(n_603),
.B1(n_613),
.B2(n_580),
.Y(n_630)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_552),
.B(n_341),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_599),
.B(n_604),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_549),
.A2(n_439),
.B1(n_451),
.B2(n_368),
.Y(n_603)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_561),
.B(n_369),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_548),
.B(n_366),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g623 ( 
.A(n_605),
.B(n_557),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_607),
.B(n_568),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_SL g608 ( 
.A1(n_582),
.A2(n_451),
.B1(n_426),
.B2(n_388),
.Y(n_608)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_610),
.B(n_567),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_548),
.B(n_451),
.C(n_407),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_611),
.B(n_568),
.C(n_581),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_582),
.A2(n_426),
.B1(n_424),
.B2(n_343),
.Y(n_613)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_615),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_609),
.Y(n_616)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_616),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g618 ( 
.A(n_601),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_618),
.B(n_620),
.Y(n_640)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_606),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_621),
.B(n_622),
.Y(n_653)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_SL g652 ( 
.A(n_623),
.B(n_620),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_624),
.B(n_631),
.Y(n_658)
);

MAJx2_ASAP7_75t_L g659 ( 
.A(n_625),
.B(n_629),
.C(n_631),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_584),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_626),
.B(n_634),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_627),
.A2(n_628),
.B1(n_635),
.B2(n_400),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_591),
.A2(n_597),
.B1(n_602),
.B2(n_612),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_600),
.B(n_553),
.C(n_564),
.Y(n_629)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_629),
.B(n_632),
.C(n_633),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_630),
.A2(n_593),
.B1(n_586),
.B2(n_608),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g631 ( 
.A(n_589),
.B(n_566),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_604),
.B(n_555),
.C(n_563),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_611),
.B(n_569),
.C(n_577),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_590),
.B(n_314),
.C(n_364),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_612),
.A2(n_343),
.B1(n_312),
.B2(n_400),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_595),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_636),
.Y(n_656)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_594),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_637),
.Y(n_651)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_592),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_638),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_588),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_639),
.A2(n_331),
.B(n_328),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_641),
.A2(n_400),
.B1(n_312),
.B2(n_372),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_628),
.A2(n_587),
.B(n_598),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_642),
.A2(n_647),
.B(n_325),
.Y(n_679)
);

XOR2xp5_ASAP7_75t_L g643 ( 
.A(n_614),
.B(n_585),
.Y(n_643)
);

XOR2xp5_ASAP7_75t_L g667 ( 
.A(n_643),
.B(n_644),
.Y(n_667)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_614),
.B(n_590),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_617),
.A2(n_607),
.B(n_603),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_630),
.A2(n_599),
.B1(n_610),
.B2(n_613),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_SL g666 ( 
.A1(n_648),
.A2(n_625),
.B1(n_627),
.B2(n_596),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_652),
.B(n_654),
.Y(n_664)
);

CKINVDCx14_ASAP7_75t_R g654 ( 
.A(n_632),
.Y(n_654)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_655),
.Y(n_663)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_659),
.Y(n_670)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_624),
.B(n_605),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_660),
.B(n_634),
.Y(n_662)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_661),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_662),
.B(n_665),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_649),
.B(n_658),
.C(n_659),
.Y(n_665)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_666),
.A2(n_671),
.B1(n_676),
.B2(n_677),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_650),
.B(n_633),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g687 ( 
.A(n_668),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_649),
.B(n_619),
.C(n_623),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g685 ( 
.A(n_669),
.B(n_672),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_640),
.B(n_596),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_658),
.B(n_619),
.C(n_635),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_660),
.B(n_314),
.C(n_333),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g686 ( 
.A(n_673),
.B(n_675),
.C(n_678),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_652),
.B(n_364),
.C(n_328),
.Y(n_675)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_656),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_644),
.B(n_372),
.C(n_357),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_679),
.A2(n_680),
.B1(n_656),
.B2(n_651),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_646),
.A2(n_357),
.B1(n_325),
.B2(n_360),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_665),
.B(n_657),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_681),
.B(n_683),
.Y(n_695)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_664),
.A2(n_653),
.B(n_645),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_682),
.A2(n_691),
.B(n_675),
.Y(n_698)
);

XNOR2xp5_ASAP7_75t_L g683 ( 
.A(n_672),
.B(n_642),
.Y(n_683)
);

XNOR2xp5_ASAP7_75t_L g688 ( 
.A(n_669),
.B(n_648),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_688),
.B(n_689),
.Y(n_700)
);

MAJIxp5_ASAP7_75t_L g689 ( 
.A(n_663),
.B(n_655),
.C(n_641),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_670),
.A2(n_666),
.B(n_679),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_674),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_692),
.B(n_693),
.Y(n_702)
);

XNOR2xp5_ASAP7_75t_L g693 ( 
.A(n_673),
.B(n_647),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_694),
.B(n_651),
.Y(n_696)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_696),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_685),
.B(n_684),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_697),
.Y(n_706)
);

AOI21xp33_ASAP7_75t_L g709 ( 
.A1(n_698),
.A2(n_703),
.B(n_686),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_687),
.B(n_680),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_699),
.B(n_704),
.Y(n_708)
);

OAI21xp5_ASAP7_75t_L g701 ( 
.A1(n_690),
.A2(n_667),
.B(n_678),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_701),
.A2(n_695),
.B(n_702),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_692),
.B(n_676),
.Y(n_703)
);

MAJIxp5_ASAP7_75t_L g704 ( 
.A(n_688),
.B(n_667),
.C(n_643),
.Y(n_704)
);

O2A1O1Ixp33_ASAP7_75t_SL g705 ( 
.A1(n_696),
.A2(n_689),
.B(n_693),
.C(n_683),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_705),
.A2(n_709),
.B(n_711),
.Y(n_715)
);

OAI21xp33_ASAP7_75t_SL g713 ( 
.A1(n_707),
.A2(n_361),
.B(n_363),
.Y(n_713)
);

MAJIxp5_ASAP7_75t_L g711 ( 
.A(n_700),
.B(n_686),
.C(n_352),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_SL g712 ( 
.A(n_706),
.B(n_703),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_712),
.Y(n_717)
);

OAI311xp33_ASAP7_75t_L g716 ( 
.A1(n_713),
.A2(n_714),
.A3(n_708),
.B1(n_361),
.C1(n_360),
.Y(n_716)
);

MAJIxp5_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_710),
.C(n_327),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_716),
.B(n_360),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_718),
.Y(n_719)
);

MAJIxp5_ASAP7_75t_L g720 ( 
.A(n_719),
.B(n_715),
.C(n_717),
.Y(n_720)
);

BUFx24_ASAP7_75t_SL g721 ( 
.A(n_720),
.Y(n_721)
);

XOR2xp5_ASAP7_75t_L g722 ( 
.A(n_721),
.B(n_361),
.Y(n_722)
);


endmodule