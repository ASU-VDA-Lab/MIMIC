module fake_jpeg_31429_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_36),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_47),
.B(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_53),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_15),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_72),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_28),
.B(n_13),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_64),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_61),
.B(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_26),
.Y(n_71)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_71),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_33),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_33),
.B(n_13),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_76),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_74),
.Y(n_120)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_20),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_27),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_79),
.Y(n_124)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_34),
.Y(n_78)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_35),
.B(n_2),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_85),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_34),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_87),
.B(n_88),
.Y(n_127)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_91),
.Y(n_128)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_90),
.B(n_41),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_31),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_87),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_99),
.A2(n_92),
.B(n_48),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_17),
.B1(n_46),
.B2(n_43),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g143 ( 
.A1(n_100),
.A2(n_138),
.B1(n_140),
.B2(n_66),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_102),
.A2(n_119),
.B1(n_132),
.B2(n_62),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_52),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_118),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_58),
.A2(n_42),
.B1(n_46),
.B2(n_43),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_30),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_1),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_78),
.A2(n_41),
.B1(n_29),
.B2(n_24),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_63),
.B1(n_49),
.B2(n_82),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_29),
.B1(n_24),
.B2(n_23),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_23),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_55),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_70),
.A2(n_1),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_142),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_143),
.A2(n_157),
.B1(n_113),
.B2(n_97),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_67),
.B(n_77),
.C(n_85),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_67),
.B(n_10),
.C(n_11),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_151),
.B(n_167),
.Y(n_188)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_147),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_159),
.Y(n_191)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_96),
.A2(n_74),
.B1(n_91),
.B2(n_85),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_100),
.A2(n_91),
.B(n_76),
.C(n_65),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_171),
.B(n_113),
.Y(n_199)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_99),
.B(n_84),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_168),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_166),
.Y(n_207)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_100),
.Y(n_168)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_169),
.B(n_170),
.Y(n_209)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

HAxp5_ASAP7_75t_SL g171 ( 
.A(n_138),
.B(n_124),
.CON(n_171),
.SN(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_94),
.B(n_115),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_173),
.Y(n_211)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

AO21x2_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_126),
.B(n_93),
.Y(n_210)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_175),
.A2(n_177),
.B1(n_179),
.B2(n_98),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_128),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_135),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_135),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_112),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_123),
.Y(n_185)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_174),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_140),
.B1(n_102),
.B2(n_111),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_196),
.B1(n_200),
.B2(n_202),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_148),
.A2(n_108),
.B1(n_120),
.B2(n_117),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_136),
.C(n_104),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_176),
.C(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_199),
.B(n_206),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_167),
.B1(n_143),
.B2(n_171),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_97),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_176),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_143),
.A2(n_117),
.B1(n_106),
.B2(n_110),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_163),
.A2(n_106),
.B1(n_110),
.B2(n_93),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_203),
.A2(n_205),
.B1(n_175),
.B2(n_154),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_155),
.A2(n_162),
.B1(n_144),
.B2(n_145),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_213),
.B(n_223),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_202),
.C(n_203),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_182),
.B(n_147),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_191),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_185),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_158),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_211),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_204),
.B(n_146),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_225),
.B(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_227),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_161),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_160),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_169),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_150),
.B(n_173),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_208),
.B(n_184),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_234),
.Y(n_254)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_196),
.B(n_149),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_184),
.B(n_188),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_239),
.A2(n_240),
.B(n_246),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_236),
.A2(n_188),
.B(n_210),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_208),
.B(n_210),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_228),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_234),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_214),
.B(n_231),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_257),
.Y(n_262)
);

NAND2x1_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_210),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_258),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_221),
.B1(n_237),
.B2(n_219),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_268),
.B1(n_247),
.B2(n_244),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_218),
.B1(n_231),
.B2(n_232),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_260),
.A2(n_270),
.B1(n_272),
.B2(n_240),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_254),
.B(n_214),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_266),
.C(n_269),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_225),
.Y(n_267)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_267),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_221),
.B1(n_226),
.B2(n_231),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_227),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_239),
.A2(n_231),
.B1(n_215),
.B2(n_220),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_250),
.A2(n_230),
.B1(n_223),
.B2(n_212),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_250),
.B1(n_245),
.B2(n_241),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_245),
.A2(n_217),
.B1(n_189),
.B2(n_213),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_216),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_243),
.B(n_189),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_243),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_244),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_252),
.C(n_253),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_279),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_252),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_285),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_257),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_282),
.C(n_288),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_253),
.B1(n_255),
.B2(n_241),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_260),
.B1(n_264),
.B2(n_270),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_262),
.B(n_255),
.C(n_240),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_289),
.A2(n_258),
.B1(n_279),
.B2(n_278),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_246),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_261),
.C(n_247),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_294),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_290),
.A2(n_275),
.B(n_263),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_248),
.B(n_183),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_288),
.CI(n_282),
.CON(n_296),
.SN(n_296)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

NOR3xp33_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_264),
.C(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_291),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_194),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_258),
.B1(n_248),
.B2(n_242),
.Y(n_300)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_242),
.C(n_180),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_277),
.C(n_192),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_258),
.B1(n_248),
.B2(n_210),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_310),
.C(n_311),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_293),
.B1(n_297),
.B2(n_299),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_309),
.A2(n_296),
.B1(n_190),
.B2(n_183),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_235),
.C(n_181),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_181),
.C(n_190),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_312),
.B(n_298),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_302),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_315),
.A2(n_318),
.B1(n_319),
.B2(n_302),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_305),
.B(n_295),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_296),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_307),
.A2(n_313),
.B1(n_303),
.B2(n_309),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_312),
.B(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_311),
.B(n_310),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_325),
.B(n_198),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_323),
.B(n_324),
.C(n_320),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_328),
.B(n_166),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_324),
.A2(n_320),
.B(n_319),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_198),
.B(n_142),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_330),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.C(n_327),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_170),
.Y(n_334)
);


endmodule