module real_aes_6626_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_503;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_0), .Y(n_122) );
INVx1_ASAP7_75t_L g262 ( .A(n_1), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_2), .A2(n_31), .B1(n_215), .B2(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_3), .B(n_206), .Y(n_231) );
INVx1_ASAP7_75t_L g197 ( .A(n_4), .Y(n_197) );
AND2x6_ASAP7_75t_L g230 ( .A(n_4), .B(n_195), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_4), .B(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_5), .Y(n_117) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_6), .A2(n_26), .B1(n_89), .B2(n_94), .Y(n_97) );
INVx1_ASAP7_75t_L g211 ( .A(n_7), .Y(n_211) );
INVx1_ASAP7_75t_L g255 ( .A(n_8), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_9), .B(n_219), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_10), .B(n_207), .Y(n_267) );
AO32x2_ASAP7_75t_L g289 ( .A1(n_11), .A2(n_206), .A3(n_235), .B1(n_246), .B2(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_12), .B(n_215), .Y(n_302) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_13), .A2(n_28), .B1(n_89), .B2(n_90), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_14), .B(n_207), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_15), .A2(n_41), .B1(n_215), .B2(n_292), .Y(n_293) );
INVx1_ASAP7_75t_L g523 ( .A(n_15), .Y(n_523) );
AOI22xp33_ASAP7_75t_SL g314 ( .A1(n_16), .A2(n_62), .B1(n_215), .B2(n_219), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_17), .B(n_215), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_18), .A2(n_80), .B1(n_174), .B2(n_175), .Y(n_79) );
INVx1_ASAP7_75t_L g174 ( .A(n_18), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_19), .Y(n_154) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_20), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_21), .B(n_248), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_22), .A2(n_60), .B1(n_106), .B2(n_112), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_23), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_24), .B(n_248), .Y(n_286) );
INVx2_ASAP7_75t_L g217 ( .A(n_25), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_27), .B(n_215), .Y(n_238) );
OAI221xp5_ASAP7_75t_L g188 ( .A1(n_28), .A2(n_46), .B1(n_57), .B2(n_189), .C(n_190), .Y(n_188) );
INVxp67_ASAP7_75t_L g191 ( .A(n_28), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_29), .B(n_248), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g83 ( .A1(n_30), .A2(n_33), .B1(n_84), .B2(n_100), .Y(n_83) );
AOI22xp5_ASAP7_75t_SL g512 ( .A1(n_31), .A2(n_80), .B1(n_175), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_31), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_32), .Y(n_139) );
XNOR2xp5_ASAP7_75t_L g524 ( .A(n_34), .B(n_175), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_35), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_36), .B(n_215), .Y(n_214) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_37), .A2(n_71), .B1(n_292), .B2(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_38), .B(n_215), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_39), .B(n_215), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_40), .B(n_227), .Y(n_226) );
AOI22xp33_ASAP7_75t_SL g271 ( .A1(n_42), .A2(n_47), .B1(n_215), .B2(n_219), .Y(n_271) );
OAI22xp5_ASAP7_75t_SL g179 ( .A1(n_43), .A2(n_64), .B1(n_180), .B2(n_181), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_43), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_44), .B(n_215), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_45), .B(n_215), .Y(n_297) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_46), .A2(n_68), .B1(n_89), .B2(n_90), .Y(n_88) );
INVxp67_ASAP7_75t_L g192 ( .A(n_46), .Y(n_192) );
INVx1_ASAP7_75t_L g195 ( .A(n_48), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_49), .A2(n_177), .B1(n_183), .B2(n_184), .Y(n_176) );
INVx1_ASAP7_75t_L g183 ( .A(n_49), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_50), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_51), .B(n_215), .Y(n_263) );
INVx1_ASAP7_75t_L g210 ( .A(n_52), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_53), .Y(n_189) );
AO32x2_ASAP7_75t_L g310 ( .A1(n_54), .A2(n_206), .A3(n_246), .B1(n_311), .B2(n_315), .Y(n_310) );
INVx1_ASAP7_75t_L g241 ( .A(n_55), .Y(n_241) );
INVx1_ASAP7_75t_L g281 ( .A(n_56), .Y(n_281) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_57), .A2(n_73), .B1(n_89), .B2(n_94), .Y(n_93) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_58), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_59), .B(n_219), .Y(n_282) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_61), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_63), .Y(n_127) );
INVx1_ASAP7_75t_L g181 ( .A(n_64), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_65), .B(n_292), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_66), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_67), .B(n_219), .Y(n_285) );
INVx2_ASAP7_75t_L g208 ( .A(n_69), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_70), .B(n_219), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_72), .A2(n_76), .B1(n_219), .B2(n_220), .Y(n_270) );
INVx1_ASAP7_75t_L g89 ( .A(n_74), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_74), .Y(n_91) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_75), .A2(n_178), .B1(n_179), .B2(n_182), .Y(n_177) );
INVx1_ASAP7_75t_L g182 ( .A(n_75), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_75), .B(n_219), .Y(n_239) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_185), .B1(n_198), .B2(n_507), .C(n_511), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_176), .Y(n_78) );
INVx1_ASAP7_75t_L g175 ( .A(n_80), .Y(n_175) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_137), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_116), .C(n_126), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_105), .Y(n_82) );
BUFx2_ASAP7_75t_SL g84 ( .A(n_85), .Y(n_84) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_95), .Y(n_85) );
AND2x6_ASAP7_75t_L g102 ( .A(n_86), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g121 ( .A(n_86), .B(n_111), .Y(n_121) );
AND2x6_ASAP7_75t_L g153 ( .A(n_86), .B(n_148), .Y(n_153) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g131 ( .A(n_87), .B(n_93), .Y(n_131) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g109 ( .A(n_88), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_88), .B(n_93), .Y(n_115) );
AND2x2_ASAP7_75t_L g143 ( .A(n_88), .B(n_97), .Y(n_143) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g94 ( .A(n_91), .Y(n_94) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx1_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
INVx1_ASAP7_75t_L g159 ( .A(n_93), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_95), .B(n_109), .Y(n_125) );
AND2x4_ASAP7_75t_L g130 ( .A(n_95), .B(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g135 ( .A(n_95), .B(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
OR2x2_ASAP7_75t_L g104 ( .A(n_96), .B(n_99), .Y(n_104) );
AND2x2_ASAP7_75t_L g111 ( .A(n_96), .B(n_99), .Y(n_111) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g148 ( .A(n_97), .B(n_99), .Y(n_148) );
INVx1_ASAP7_75t_L g144 ( .A(n_98), .Y(n_144) );
AND2x2_ASAP7_75t_L g164 ( .A(n_98), .B(n_159), .Y(n_164) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g114 ( .A(n_99), .Y(n_114) );
INVx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx11_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OR2x2_ASAP7_75t_L g168 ( .A(n_104), .B(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx8_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_L g150 ( .A(n_110), .Y(n_150) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_111), .B(n_131), .Y(n_173) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g136 ( .A(n_115), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_118), .B1(n_122), .B2(n_123), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx6_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_132), .B2(n_133), .Y(n_126) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g169 ( .A(n_131), .Y(n_169) );
INVx1_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
BUFx2_ASAP7_75t_SL g134 ( .A(n_135), .Y(n_134) );
NOR3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_151), .C(n_165), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B1(n_145), .B2(n_146), .Y(n_138) );
INVx3_ASAP7_75t_SL g140 ( .A(n_141), .Y(n_140) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x4_ASAP7_75t_L g157 ( .A(n_143), .B(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g163 ( .A(n_143), .B(n_164), .Y(n_163) );
OR2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
OAI221xp5_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B1(n_155), .B2(n_160), .C(n_161), .Y(n_151) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B1(n_170), .B2(n_171), .Y(n_165) );
BUFx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_177), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_187), .Y(n_186) );
AND3x1_ASAP7_75t_SL g187 ( .A(n_188), .B(n_193), .C(n_196), .Y(n_187) );
INVxp67_ASAP7_75t_L g517 ( .A(n_188), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_191), .B(n_192), .Y(n_190) );
INVx1_ASAP7_75t_SL g518 ( .A(n_193), .Y(n_518) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_193), .A2(n_510), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g528 ( .A(n_193), .Y(n_528) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_194), .B(n_197), .Y(n_522) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_SL g527 ( .A(n_196), .B(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_197), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g198 ( .A(n_199), .B(n_431), .Y(n_198) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_200), .B(n_389), .Y(n_199) );
NOR4xp25_ASAP7_75t_L g200 ( .A(n_201), .B(n_329), .C(n_365), .D(n_379), .Y(n_200) );
OAI221xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_273), .B1(n_305), .B2(n_316), .C(n_320), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_202), .B(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_249), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_232), .Y(n_204) );
AND2x2_ASAP7_75t_L g326 ( .A(n_205), .B(n_233), .Y(n_326) );
INVx3_ASAP7_75t_L g334 ( .A(n_205), .Y(n_334) );
AND2x2_ASAP7_75t_L g388 ( .A(n_205), .B(n_252), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_205), .B(n_251), .Y(n_424) );
AND2x2_ASAP7_75t_L g482 ( .A(n_205), .B(n_344), .Y(n_482) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_212), .B(n_231), .Y(n_205) );
INVx4_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g235 ( .A(n_207), .Y(n_235) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AND2x2_ASAP7_75t_SL g248 ( .A(n_208), .B(n_209), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_224), .B(n_230), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_218), .B(n_221), .Y(n_213) );
INVx3_ASAP7_75t_L g280 ( .A(n_215), .Y(n_280) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g292 ( .A(n_216), .Y(n_292) );
BUFx3_ASAP7_75t_L g313 ( .A(n_216), .Y(n_313) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g220 ( .A(n_217), .Y(n_220) );
INVx1_ASAP7_75t_L g228 ( .A(n_217), .Y(n_228) );
INVx2_ASAP7_75t_L g256 ( .A(n_219), .Y(n_256) );
INVx3_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g229 ( .A(n_221), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_238), .B(n_239), .Y(n_237) );
O2A1O1Ixp5_ASAP7_75t_SL g279 ( .A1(n_221), .A2(n_280), .B(n_281), .C(n_282), .Y(n_279) );
INVx5_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OAI22xp5_ASAP7_75t_SL g311 ( .A1(n_222), .A2(n_245), .B1(n_312), .B2(n_314), .Y(n_311) );
INVx3_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_223), .Y(n_245) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_223), .Y(n_260) );
INVx1_ASAP7_75t_L g300 ( .A(n_223), .Y(n_300) );
AND2x2_ASAP7_75t_L g510 ( .A(n_223), .B(n_228), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_229), .Y(n_224) );
INVx2_ASAP7_75t_L g242 ( .A(n_227), .Y(n_242) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_229), .A2(n_242), .B(n_262), .C(n_263), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_229), .A2(n_245), .B1(n_270), .B2(n_271), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g290 ( .A1(n_229), .A2(n_245), .B1(n_291), .B2(n_293), .Y(n_290) );
BUFx3_ASAP7_75t_L g246 ( .A(n_230), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_230), .A2(n_254), .B(n_261), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_230), .A2(n_279), .B(n_283), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g295 ( .A1(n_230), .A2(n_296), .B(n_301), .Y(n_295) );
AND2x4_ASAP7_75t_L g509 ( .A(n_230), .B(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g317 ( .A(n_232), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_232), .B(n_252), .Y(n_331) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_233), .B(n_252), .Y(n_346) );
AND2x2_ASAP7_75t_L g358 ( .A(n_233), .B(n_334), .Y(n_358) );
OR2x2_ASAP7_75t_L g360 ( .A(n_233), .B(n_318), .Y(n_360) );
AND2x2_ASAP7_75t_L g395 ( .A(n_233), .B(n_318), .Y(n_395) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_233), .Y(n_440) );
INVx1_ASAP7_75t_L g448 ( .A(n_233), .Y(n_448) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_236), .B(n_247), .Y(n_233) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_234), .A2(n_253), .B(n_264), .Y(n_252) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_240), .B(n_246), .Y(n_236) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_243), .C(n_244), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_244), .A2(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND3xp33_ASAP7_75t_L g268 ( .A(n_246), .B(n_269), .C(n_272), .Y(n_268) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_248), .A2(n_278), .B(n_286), .Y(n_277) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_248), .A2(n_295), .B(n_304), .Y(n_294) );
INVx2_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_249), .A2(n_366), .B1(n_370), .B2(n_374), .C(n_375), .Y(n_365) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g325 ( .A(n_250), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_265), .Y(n_250) );
INVx2_ASAP7_75t_L g324 ( .A(n_251), .Y(n_324) );
AND2x2_ASAP7_75t_L g377 ( .A(n_251), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g396 ( .A(n_251), .B(n_334), .Y(n_396) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g459 ( .A(n_252), .B(n_334), .Y(n_459) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_257), .C(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_259), .A2(n_284), .B(n_285), .Y(n_283) );
INVx4_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g381 ( .A(n_265), .B(n_326), .Y(n_381) );
OAI322xp33_ASAP7_75t_L g449 ( .A1(n_265), .A2(n_405), .A3(n_450), .B1(n_452), .B2(n_455), .C1(n_457), .C2(n_461), .Y(n_449) );
INVx3_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NOR2x1_ASAP7_75t_L g332 ( .A(n_266), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g345 ( .A(n_266), .Y(n_345) );
AND2x2_ASAP7_75t_L g454 ( .A(n_266), .B(n_334), .Y(n_454) );
AND2x2_ASAP7_75t_L g486 ( .A(n_266), .B(n_358), .Y(n_486) );
OR2x2_ASAP7_75t_L g489 ( .A(n_266), .B(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g319 ( .A(n_267), .Y(n_319) );
AO21x1_ASAP7_75t_L g318 ( .A1(n_269), .A2(n_272), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_287), .Y(n_274) );
INVx1_ASAP7_75t_L g502 ( .A(n_275), .Y(n_502) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g307 ( .A(n_276), .B(n_294), .Y(n_307) );
INVx2_ASAP7_75t_L g342 ( .A(n_276), .Y(n_342) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g364 ( .A(n_277), .Y(n_364) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_277), .Y(n_372) );
OR2x2_ASAP7_75t_L g496 ( .A(n_277), .B(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g321 ( .A(n_287), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g361 ( .A(n_287), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g413 ( .A(n_287), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_294), .Y(n_287) );
AND2x2_ASAP7_75t_L g308 ( .A(n_288), .B(n_309), .Y(n_308) );
NOR2xp67_ASAP7_75t_L g368 ( .A(n_288), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g422 ( .A(n_288), .B(n_310), .Y(n_422) );
OR2x2_ASAP7_75t_L g430 ( .A(n_288), .B(n_364), .Y(n_430) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
AND2x2_ASAP7_75t_L g349 ( .A(n_289), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g373 ( .A(n_289), .B(n_294), .Y(n_373) );
AND2x2_ASAP7_75t_L g437 ( .A(n_289), .B(n_310), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_294), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_294), .B(n_342), .Y(n_341) );
INVx2_ASAP7_75t_L g350 ( .A(n_294), .Y(n_350) );
INVx1_ASAP7_75t_L g355 ( .A(n_294), .Y(n_355) );
AND2x2_ASAP7_75t_L g367 ( .A(n_294), .B(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_294), .Y(n_445) );
INVx1_ASAP7_75t_L g497 ( .A(n_294), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
AND2x2_ASAP7_75t_L g474 ( .A(n_306), .B(n_383), .Y(n_474) );
INVx2_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g401 ( .A(n_308), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g500 ( .A(n_308), .B(n_435), .Y(n_500) );
INVx1_ASAP7_75t_L g322 ( .A(n_309), .Y(n_322) );
AND2x2_ASAP7_75t_L g348 ( .A(n_309), .B(n_342), .Y(n_348) );
BUFx2_ASAP7_75t_L g407 ( .A(n_309), .Y(n_407) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_310), .Y(n_328) );
INVx1_ASAP7_75t_L g338 ( .A(n_310), .Y(n_338) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_316), .B(n_323), .Y(n_476) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AOI32xp33_ASAP7_75t_L g320 ( .A1(n_317), .A2(n_321), .A3(n_323), .B1(n_325), .B2(n_327), .Y(n_320) );
AND2x2_ASAP7_75t_L g460 ( .A(n_317), .B(n_333), .Y(n_460) );
AND2x2_ASAP7_75t_L g498 ( .A(n_317), .B(n_396), .Y(n_498) );
INVx1_ASAP7_75t_L g378 ( .A(n_318), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_322), .B(n_384), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_323), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_323), .B(n_326), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_323), .B(n_395), .Y(n_477) );
OR2x2_ASAP7_75t_L g491 ( .A(n_323), .B(n_360), .Y(n_491) );
INVx3_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g418 ( .A(n_324), .B(n_326), .Y(n_418) );
OR2x2_ASAP7_75t_L g427 ( .A(n_324), .B(n_414), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_326), .B(n_377), .Y(n_399) );
INVx2_ASAP7_75t_L g414 ( .A(n_328), .Y(n_414) );
OR2x2_ASAP7_75t_L g429 ( .A(n_328), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g444 ( .A(n_328), .B(n_445), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_328), .A2(n_421), .B(n_502), .C(n_503), .Y(n_501) );
OAI321xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_335), .A3(n_340), .B1(n_343), .B2(n_347), .C(n_351), .Y(n_329) );
INVx1_ASAP7_75t_L g442 ( .A(n_330), .Y(n_442) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g453 ( .A(n_331), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g405 ( .A(n_333), .Y(n_405) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_334), .B(n_448), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g472 ( .A1(n_335), .A2(n_473), .B1(n_475), .B2(n_477), .C(n_478), .Y(n_472) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
AND2x2_ASAP7_75t_L g410 ( .A(n_337), .B(n_384), .Y(n_410) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_338), .B(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_340), .A2(n_381), .B(n_426), .C(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g392 ( .A(n_342), .B(n_349), .Y(n_392) );
BUFx2_ASAP7_75t_L g402 ( .A(n_342), .Y(n_402) );
INVx1_ASAP7_75t_L g417 ( .A(n_342), .Y(n_417) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OR2x2_ASAP7_75t_L g423 ( .A(n_345), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g506 ( .A(n_345), .Y(n_506) );
INVx1_ASAP7_75t_L g499 ( .A(n_346), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
AND2x2_ASAP7_75t_L g352 ( .A(n_348), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g456 ( .A(n_348), .B(n_373), .Y(n_456) );
INVx1_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .B1(n_359), .B2(n_361), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_353), .B(n_469), .Y(n_468) );
INVxp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g421 ( .A(n_354), .B(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_SL g384 ( .A(n_355), .B(n_364), .Y(n_384) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g376 ( .A(n_358), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g386 ( .A(n_360), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_363), .A2(n_481), .B1(n_483), .B2(n_484), .C(n_485), .Y(n_480) );
INVx1_ASAP7_75t_L g369 ( .A(n_364), .Y(n_369) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_364), .Y(n_435) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_367), .B(n_486), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_368), .A2(n_373), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_371), .B(n_381), .Y(n_478) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx1_ASAP7_75t_L g447 ( .A(n_372), .Y(n_447) );
AND2x2_ASAP7_75t_L g406 ( .A(n_373), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g495 ( .A(n_373), .Y(n_495) );
INVx1_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx1_ASAP7_75t_L g466 ( .A(n_377), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_382), .B1(n_385), .B2(n_386), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_383), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g451 ( .A(n_384), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_384), .B(n_422), .Y(n_488) );
OR2x2_ASAP7_75t_L g461 ( .A(n_385), .B(n_414), .Y(n_461) );
INVx1_ASAP7_75t_L g400 ( .A(n_386), .Y(n_400) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_388), .B(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g389 ( .A(n_390), .B(n_408), .C(n_419), .Y(n_389) );
OAI211xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B(n_397), .C(n_403), .Y(n_390) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_392), .A2(n_463), .B1(n_467), .B2(n_470), .C(n_472), .Y(n_462) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
AND2x2_ASAP7_75t_L g404 ( .A(n_395), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g458 ( .A(n_395), .B(n_459), .Y(n_458) );
OAI211xp5_ASAP7_75t_L g443 ( .A1(n_396), .A2(n_444), .B(n_446), .C(n_448), .Y(n_443) );
INVx2_ASAP7_75t_L g490 ( .A(n_396), .Y(n_490) );
OAI21xp5_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_400), .B(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g469 ( .A(n_402), .B(n_422), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_411), .B(n_412), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
OAI21xp5_ASAP7_75t_SL g412 ( .A1(n_413), .A2(n_415), .B(n_418), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_413), .B(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_418), .B(n_505), .Y(n_504) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B(n_425), .Y(n_419) );
INVx1_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g446 ( .A(n_422), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND4x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_462), .C(n_479), .D(n_501), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_449), .Y(n_432) );
OAI211xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_438), .B(n_441), .C(n_443), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_SL g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_437), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_448), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx1_ASAP7_75t_L g483 ( .A(n_458), .Y(n_483) );
INVx2_ASAP7_75t_SL g471 ( .A(n_459), .Y(n_471) );
OR2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g484 ( .A(n_469), .Y(n_484) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_SL g479 ( .A(n_480), .B(n_487), .Y(n_479) );
INVx1_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OAI221xp5_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B1(n_491), .B2(n_492), .C(n_493), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_495), .B(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OAI322xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_514), .A3(n_518), .B1(n_519), .B2(n_523), .C1(n_524), .C2(n_525), .Y(n_511) );
INVx1_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
endmodule