module fake_netlist_1_5614_n_455 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_455);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_455;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g68 ( .A(n_22), .Y(n_68) );
INVx1_ASAP7_75t_L g69 ( .A(n_2), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_35), .Y(n_70) );
BUFx6f_ASAP7_75t_L g71 ( .A(n_1), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_30), .Y(n_72) );
INVx2_ASAP7_75t_L g73 ( .A(n_62), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_58), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_40), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_53), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_17), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_37), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_26), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_54), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_31), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_21), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_33), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_32), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_9), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_59), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_56), .Y(n_87) );
BUFx2_ASAP7_75t_L g88 ( .A(n_20), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_47), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_42), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_39), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_65), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_46), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_29), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_13), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_38), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_16), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_50), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_23), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_80), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_96), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_82), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_73), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_88), .B(n_0), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_88), .B(n_0), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_99), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_99), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_96), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_96), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_90), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_70), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_76), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_68), .B(n_1), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_72), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_81), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_72), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_79), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_93), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_68), .B(n_2), .Y(n_125) );
NAND2x1p5_ASAP7_75t_L g126 ( .A(n_119), .B(n_74), .Y(n_126) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_106), .Y(n_127) );
OR2x2_ASAP7_75t_L g128 ( .A(n_121), .B(n_69), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_121), .B(n_69), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_106), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_119), .B(n_77), .Y(n_132) );
AO22x2_ASAP7_75t_L g133 ( .A1(n_109), .A2(n_102), .B1(n_81), .B2(n_86), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_119), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_115), .B(n_99), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_107), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_118), .B(n_94), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_116), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g139 ( .A1(n_110), .A2(n_77), .B1(n_100), .B2(n_98), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_109), .B(n_85), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_116), .B(n_97), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_117), .B(n_74), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_107), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_107), .Y(n_145) );
NAND3x1_ASAP7_75t_L g146 ( .A(n_108), .B(n_100), .C(n_98), .Y(n_146) );
INVx8_ASAP7_75t_L g147 ( .A(n_111), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_114), .Y(n_148) );
AOI22x1_ASAP7_75t_L g149 ( .A1(n_117), .A2(n_93), .B1(n_86), .B2(n_91), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_120), .Y(n_150) );
INVx1_ASAP7_75t_SL g151 ( .A(n_103), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_151), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_134), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_127), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_126), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_126), .Y(n_157) );
INVx2_ASAP7_75t_SL g158 ( .A(n_138), .Y(n_158) );
NOR2x1_ASAP7_75t_L g159 ( .A(n_142), .B(n_108), .Y(n_159) );
NOR3xp33_ASAP7_75t_SL g160 ( .A(n_137), .B(n_125), .C(n_91), .Y(n_160) );
BUFx4f_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_150), .B(n_109), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_127), .Y(n_164) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_133), .A2(n_122), .B1(n_120), .B2(n_125), .Y(n_165) );
BUFx8_ASAP7_75t_L g166 ( .A(n_140), .Y(n_166) );
OR2x6_ASAP7_75t_L g167 ( .A(n_133), .B(n_122), .Y(n_167) );
NAND2xp33_ASAP7_75t_SL g168 ( .A(n_128), .B(n_85), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_136), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_135), .B(n_101), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_132), .B(n_104), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_136), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_140), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_127), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
AND2x4_ASAP7_75t_L g177 ( .A(n_130), .B(n_102), .Y(n_177) );
INVx3_ASAP7_75t_L g178 ( .A(n_127), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_144), .Y(n_179) );
NOR3xp33_ASAP7_75t_SL g180 ( .A(n_143), .B(n_75), .C(n_78), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_127), .Y(n_181) );
NOR2xp33_ASAP7_75t_R g182 ( .A(n_147), .B(n_105), .Y(n_182) );
INVx3_ASAP7_75t_SL g183 ( .A(n_147), .Y(n_183) );
AND2x4_ASAP7_75t_L g184 ( .A(n_130), .B(n_141), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_141), .B(n_124), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_169), .Y(n_186) );
NOR2x1_ASAP7_75t_SL g187 ( .A(n_167), .B(n_128), .Y(n_187) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
AND2x4_ASAP7_75t_L g189 ( .A(n_157), .B(n_130), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_169), .Y(n_190) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_185), .A2(n_129), .B(n_148), .C(n_93), .Y(n_191) );
OR2x6_ASAP7_75t_L g192 ( .A(n_155), .B(n_133), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_155), .Y(n_194) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_157), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_167), .A2(n_146), .B1(n_139), .B2(n_148), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_172), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_176), .A2(n_149), .B1(n_129), .B2(n_145), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_161), .Y(n_200) );
BUFx8_ASAP7_75t_SL g201 ( .A(n_152), .Y(n_201) );
CKINVDCx11_ASAP7_75t_R g202 ( .A(n_183), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_172), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_156), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_156), .B(n_104), .Y(n_205) );
AOI222xp33_ASAP7_75t_L g206 ( .A1(n_184), .A2(n_147), .B1(n_112), .B2(n_113), .C1(n_114), .C2(n_124), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_153), .B(n_147), .Y(n_207) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
BUFx12f_ASAP7_75t_L g209 ( .A(n_166), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_161), .B(n_149), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_175), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_158), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_174), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_175), .Y(n_214) );
INVx1_ASAP7_75t_SL g215 ( .A(n_183), .Y(n_215) );
AOI21x1_ASAP7_75t_L g216 ( .A1(n_154), .A2(n_114), .B(n_124), .Y(n_216) );
NAND2xp33_ASAP7_75t_L g217 ( .A(n_158), .B(n_146), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_179), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_200), .B(n_176), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_198), .B(n_184), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_192), .A2(n_176), .B1(n_167), .B2(n_161), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_186), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_186), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_186), .Y(n_224) );
OAI22xp33_ASAP7_75t_L g225 ( .A1(n_192), .A2(n_167), .B1(n_176), .B2(n_183), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_192), .A2(n_167), .B1(n_184), .B2(n_177), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_192), .A2(n_184), .B1(n_177), .B2(n_165), .Y(n_227) );
OAI221xp5_ASAP7_75t_L g228 ( .A1(n_192), .A2(n_168), .B1(n_180), .B2(n_185), .C(n_162), .Y(n_228) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_216), .A2(n_180), .B(n_75), .Y(n_229) );
BUFx4f_ASAP7_75t_SL g230 ( .A(n_209), .Y(n_230) );
NOR3xp33_ASAP7_75t_SL g231 ( .A(n_207), .B(n_182), .C(n_163), .Y(n_231) );
NAND3xp33_ASAP7_75t_SL g232 ( .A(n_206), .B(n_160), .C(n_173), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_197), .A2(n_158), .B1(n_179), .B2(n_177), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_198), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_186), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_191), .A2(n_159), .B(n_163), .Y(n_236) );
AOI221xp5_ASAP7_75t_L g237 ( .A1(n_203), .A2(n_171), .B1(n_162), .B2(n_177), .C(n_113), .Y(n_237) );
AND2x6_ASAP7_75t_L g238 ( .A(n_195), .B(n_171), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_189), .A2(n_166), .B1(n_159), .B2(n_170), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_186), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_186), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_189), .B(n_160), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_197), .A2(n_112), .B1(n_78), .B2(n_83), .Y(n_243) );
NOR2x1_ASAP7_75t_SL g244 ( .A(n_188), .B(n_181), .Y(n_244) );
BUFx12f_ASAP7_75t_L g245 ( .A(n_230), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_224), .A2(n_216), .B(n_212), .Y(n_246) );
OAI221xp5_ASAP7_75t_L g247 ( .A1(n_228), .A2(n_217), .B1(n_204), .B2(n_208), .C(n_200), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_233), .A2(n_214), .B1(n_203), .B2(n_211), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_234), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_235), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_237), .B(n_189), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_228), .A2(n_210), .B(n_189), .C(n_215), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_233), .B(n_194), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_225), .A2(n_209), .B1(n_194), .B2(n_218), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_243), .A2(n_218), .B1(n_214), .B2(n_211), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_SL g256 ( .A1(n_236), .A2(n_199), .B(n_178), .C(n_164), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_234), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_226), .A2(n_205), .B1(n_218), .B2(n_193), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_220), .B(n_205), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_237), .B(n_205), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g261 ( .A1(n_243), .A2(n_166), .B1(n_187), .B2(n_205), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_232), .A2(n_166), .B1(n_202), .B2(n_201), .Y(n_262) );
INVx4_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_220), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_218), .B1(n_193), .B2(n_190), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_249), .B(n_229), .Y(n_266) );
OR2x2_ASAP7_75t_L g267 ( .A(n_253), .B(n_227), .Y(n_267) );
NOR4xp25_ASAP7_75t_SL g268 ( .A(n_247), .B(n_235), .C(n_84), .D(n_87), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_249), .B(n_229), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_250), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_249), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_257), .Y(n_272) );
BUFx10_ASAP7_75t_L g273 ( .A(n_250), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_263), .B(n_250), .Y(n_274) );
AND2x2_ASAP7_75t_L g275 ( .A(n_257), .B(n_229), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_248), .Y(n_276) );
HB1xp67_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
NOR3xp33_ASAP7_75t_SL g278 ( .A(n_254), .B(n_236), .C(n_84), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_250), .Y(n_279) );
OAI221xp5_ASAP7_75t_L g280 ( .A1(n_261), .A2(n_231), .B1(n_239), .B2(n_221), .C(n_242), .Y(n_280) );
OAI221xp5_ASAP7_75t_L g281 ( .A1(n_262), .A2(n_242), .B1(n_190), .B2(n_212), .C(n_87), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_248), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_253), .B(n_219), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_263), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_263), .Y(n_286) );
NOR4xp25_ASAP7_75t_SL g287 ( .A(n_264), .B(n_83), .C(n_89), .D(n_92), .Y(n_287) );
AOI33xp33_ASAP7_75t_L g288 ( .A1(n_272), .A2(n_89), .A3(n_92), .B1(n_95), .B2(n_255), .B3(n_259), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_284), .B(n_229), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_271), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_275), .B(n_259), .Y(n_291) );
OAI221xp5_ASAP7_75t_SL g292 ( .A1(n_281), .A2(n_260), .B1(n_252), .B2(n_251), .C(n_265), .Y(n_292) );
OAI21xp5_ASAP7_75t_SL g293 ( .A1(n_281), .A2(n_258), .B(n_219), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_284), .B(n_258), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_267), .B(n_263), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_283), .B(n_193), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
OAI33xp33_ASAP7_75t_L g299 ( .A1(n_276), .A2(n_95), .A3(n_282), .B1(n_267), .B2(n_271), .B3(n_7), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_276), .B(n_246), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_282), .B(n_187), .Y(n_301) );
AOI33xp33_ASAP7_75t_L g302 ( .A1(n_287), .A2(n_219), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_266), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_283), .B(n_246), .Y(n_304) );
AND2x2_ASAP7_75t_SL g305 ( .A(n_274), .B(n_219), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_266), .B(n_244), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_266), .Y(n_307) );
OAI33xp33_ASAP7_75t_L g308 ( .A1(n_287), .A2(n_3), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_8), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_269), .B(n_244), .Y(n_309) );
BUFx2_ASAP7_75t_L g310 ( .A(n_270), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_274), .B(n_222), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_269), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_280), .A2(n_71), .B1(n_131), .B2(n_145), .C(n_256), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_283), .B(n_238), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_299), .B(n_280), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_306), .B(n_283), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_306), .B(n_283), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_291), .B(n_270), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_283), .Y(n_319) );
NAND4xp25_ASAP7_75t_L g320 ( .A(n_302), .B(n_285), .C(n_286), .D(n_274), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_296), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_309), .B(n_277), .Y(n_322) );
NOR2xp33_ASAP7_75t_R g323 ( .A(n_305), .B(n_245), .Y(n_323) );
NAND5xp2_ASAP7_75t_SL g324 ( .A(n_305), .B(n_245), .C(n_8), .D(n_9), .E(n_10), .Y(n_324) );
NOR3xp33_ASAP7_75t_SL g325 ( .A(n_308), .B(n_278), .C(n_10), .Y(n_325) );
INVxp33_ASAP7_75t_L g326 ( .A(n_310), .Y(n_326) );
AND2x2_ASAP7_75t_SL g327 ( .A(n_305), .B(n_274), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_310), .B(n_277), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_298), .B(n_279), .Y(n_329) );
OAI31xp33_ASAP7_75t_L g330 ( .A1(n_293), .A2(n_285), .A3(n_286), .B(n_268), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
NAND2xp33_ASAP7_75t_SL g332 ( .A(n_288), .B(n_286), .Y(n_332) );
AOI33xp33_ASAP7_75t_L g333 ( .A1(n_303), .A2(n_268), .A3(n_11), .B1(n_12), .B2(n_13), .B3(n_14), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_292), .B(n_71), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_307), .Y(n_335) );
NOR2xp67_ASAP7_75t_SL g336 ( .A(n_293), .B(n_193), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_307), .B(n_273), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_307), .B(n_71), .Y(n_338) );
NAND2x1_ASAP7_75t_SL g339 ( .A(n_296), .B(n_223), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_312), .B(n_273), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_312), .Y(n_341) );
INVx2_ASAP7_75t_SL g342 ( .A(n_296), .Y(n_342) );
NAND2xp33_ASAP7_75t_R g343 ( .A(n_296), .B(n_240), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_290), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_289), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_294), .B(n_71), .Y(n_346) );
INVxp67_ASAP7_75t_L g347 ( .A(n_304), .Y(n_347) );
OAI31xp33_ASAP7_75t_L g348 ( .A1(n_332), .A2(n_314), .A3(n_304), .B(n_295), .Y(n_348) );
AOI322xp5_ASAP7_75t_L g349 ( .A1(n_315), .A2(n_314), .A3(n_301), .B1(n_289), .B2(n_313), .C1(n_311), .C2(n_71), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_345), .B(n_300), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_SL g351 ( .A1(n_334), .A2(n_240), .B(n_224), .C(n_164), .Y(n_351) );
OAI21xp33_ASAP7_75t_L g352 ( .A1(n_334), .A2(n_71), .B(n_300), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_331), .B(n_335), .Y(n_354) );
AOI21xp5_ASAP7_75t_L g355 ( .A1(n_330), .A2(n_297), .B(n_311), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_341), .B(n_311), .Y(n_356) );
AOI222xp33_ASAP7_75t_L g357 ( .A1(n_315), .A2(n_311), .B1(n_238), .B2(n_145), .C1(n_131), .C2(n_15), .Y(n_357) );
NAND3x2_ASAP7_75t_L g358 ( .A(n_319), .B(n_3), .C(n_11), .Y(n_358) );
AOI22xp33_ASAP7_75t_SL g359 ( .A1(n_327), .A2(n_297), .B1(n_238), .B2(n_193), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g360 ( .A1(n_320), .A2(n_297), .B(n_241), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_322), .B(n_297), .Y(n_361) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_343), .A2(n_326), .B1(n_338), .B2(n_321), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_329), .B(n_12), .Y(n_363) );
OAI322xp33_ASAP7_75t_L g364 ( .A1(n_347), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_17), .C1(n_18), .C2(n_19), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_346), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_344), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_316), .B(n_19), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_324), .A2(n_241), .B(n_240), .C(n_224), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_340), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_317), .B(n_20), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_347), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_342), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_327), .B(n_238), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_326), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_325), .A2(n_241), .B(n_240), .C(n_154), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_328), .B(n_238), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_328), .B(n_145), .Y(n_378) );
AOI32xp33_ASAP7_75t_L g379 ( .A1(n_337), .A2(n_223), .A3(n_222), .B1(n_238), .B2(n_174), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_325), .B(n_145), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_323), .B(n_24), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_336), .Y(n_383) );
AOI21xp33_ASAP7_75t_SL g384 ( .A1(n_333), .A2(n_25), .B(n_27), .Y(n_384) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_380), .B(n_333), .Y(n_385) );
NAND3x1_ASAP7_75t_L g386 ( .A(n_348), .B(n_28), .C(n_34), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_358), .A2(n_131), .B1(n_196), .B2(n_195), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_353), .B(n_36), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_375), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_366), .B(n_131), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_372), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_361), .B(n_41), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_373), .Y(n_393) );
INVxp67_ASAP7_75t_L g394 ( .A(n_378), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
XNOR2xp5_ASAP7_75t_L g396 ( .A(n_368), .B(n_43), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_371), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_382), .Y(n_398) );
CKINVDCx14_ASAP7_75t_R g399 ( .A(n_374), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_370), .Y(n_400) );
NOR4xp25_ASAP7_75t_SL g401 ( .A(n_384), .B(n_44), .C(n_45), .D(n_49), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_362), .B(n_196), .Y(n_402) );
OAI22xp33_ASAP7_75t_L g403 ( .A1(n_355), .A2(n_196), .B1(n_195), .B2(n_213), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_356), .B(n_51), .Y(n_404) );
NAND3xp33_ASAP7_75t_SL g405 ( .A(n_376), .B(n_52), .C(n_55), .Y(n_405) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_383), .B(n_196), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_350), .B(n_57), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_363), .Y(n_408) );
AOI21xp5_ASAP7_75t_SL g409 ( .A1(n_376), .A2(n_195), .B(n_188), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_365), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_L g412 ( .A1(n_355), .A2(n_188), .B(n_213), .C(n_64), .Y(n_412) );
AOI21xp33_ASAP7_75t_L g413 ( .A1(n_385), .A2(n_357), .B(n_381), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_395), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_412), .A2(n_359), .B1(n_352), .B2(n_360), .C(n_379), .Y(n_415) );
AOI211x1_ASAP7_75t_L g416 ( .A1(n_402), .A2(n_362), .B(n_360), .C(n_377), .Y(n_416) );
NOR2x1_ASAP7_75t_L g417 ( .A(n_409), .B(n_364), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_411), .Y(n_418) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_412), .A2(n_351), .B(n_369), .C(n_349), .Y(n_419) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_408), .A2(n_351), .B1(n_359), .B2(n_369), .C1(n_174), .C2(n_213), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_402), .A2(n_188), .B(n_213), .Y(n_421) );
AOI322xp5_ASAP7_75t_L g422 ( .A1(n_397), .A2(n_60), .A3(n_63), .B1(n_66), .B2(n_67), .C1(n_154), .C2(n_213), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_386), .A2(n_181), .B(n_178), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_403), .A2(n_213), .B1(n_181), .B2(n_178), .Y(n_424) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_387), .A2(n_188), .B(n_181), .C(n_178), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_391), .Y(n_426) );
XNOR2x1_ASAP7_75t_L g427 ( .A(n_398), .B(n_164), .Y(n_427) );
NOR3xp33_ASAP7_75t_L g428 ( .A(n_405), .B(n_164), .C(n_181), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_410), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_394), .A2(n_181), .B1(n_398), .B2(n_393), .Y(n_430) );
INVx2_ASAP7_75t_SL g431 ( .A(n_389), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_386), .A2(n_400), .B1(n_399), .B2(n_404), .Y(n_432) );
AND3x4_ASAP7_75t_L g433 ( .A(n_417), .B(n_399), .C(n_396), .Y(n_433) );
NAND4xp75_ASAP7_75t_L g434 ( .A(n_416), .B(n_392), .C(n_406), .D(n_404), .Y(n_434) );
XNOR2xp5_ASAP7_75t_L g435 ( .A(n_427), .B(n_388), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g436 ( .A1(n_415), .A2(n_423), .B1(n_431), .B2(n_421), .Y(n_436) );
XNOR2xp5_ASAP7_75t_L g437 ( .A(n_430), .B(n_407), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_415), .A2(n_390), .B1(n_401), .B2(n_423), .Y(n_438) );
AOI311xp33_ASAP7_75t_L g439 ( .A1(n_418), .A2(n_429), .A3(n_421), .B(n_428), .C(n_425), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_420), .B(n_419), .C(n_422), .D(n_424), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_432), .A2(n_417), .B1(n_385), .B2(n_413), .Y(n_441) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_413), .A2(n_419), .B(n_412), .C(n_417), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_414), .B(n_426), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_442), .B(n_436), .Y(n_444) );
NAND2xp33_ASAP7_75t_SL g445 ( .A(n_433), .B(n_435), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_441), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_437), .Y(n_447) );
AO22x2_ASAP7_75t_L g448 ( .A1(n_444), .A2(n_434), .B1(n_443), .B2(n_439), .Y(n_448) );
INVx1_ASAP7_75t_SL g449 ( .A(n_447), .Y(n_449) );
XNOR2xp5_ASAP7_75t_L g450 ( .A(n_446), .B(n_440), .Y(n_450) );
NOR2xp67_ASAP7_75t_L g451 ( .A(n_450), .B(n_438), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_449), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_452), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g454 ( .A1(n_453), .A2(n_451), .B1(n_448), .B2(n_445), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_454), .Y(n_455) );
endmodule