module fake_netlist_6_4797_n_1234 (n_52, n_1, n_91, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_53, n_44, n_232, n_16, n_163, n_46, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1234);

input n_52;
input n_1;
input n_91;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1234;

wire n_992;
wire n_801;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_530;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_694;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_615;
wire n_1127;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_738;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_958;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1223;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_335;
wire n_463;
wire n_848;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_380;
wire n_1190;
wire n_397;
wire n_1213;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_548;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_652;
wire n_560;
wire n_569;
wire n_737;
wire n_1229;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_649;

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_50),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_102),
.Y(n_328)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_140),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_312),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_321),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_220),
.Y(n_333)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_154),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_57),
.Y(n_335)
);

BUFx8_ASAP7_75t_SL g336 ( 
.A(n_170),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_134),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_77),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_145),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_308),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_63),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_309),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_88),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_248),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_3),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_71),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_272),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_164),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_131),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_310),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_48),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_204),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_171),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_156),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_153),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_290),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_5),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_281),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_189),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_216),
.Y(n_363)
);

BUFx10_ASAP7_75t_L g364 ( 
.A(n_166),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_206),
.Y(n_365)
);

BUFx8_ASAP7_75t_SL g366 ( 
.A(n_15),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_266),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_110),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_37),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_69),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_205),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_279),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_62),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_128),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_187),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_46),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_146),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_265),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_306),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_56),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_254),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_0),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_277),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_313),
.Y(n_384)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_219),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_24),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_61),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_104),
.Y(n_388)
);

BUFx10_ASAP7_75t_L g389 ( 
.A(n_252),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_68),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_4),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_72),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_105),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_80),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_286),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_66),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_178),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_151),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_182),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_307),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_17),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_180),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_107),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_260),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_169),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_188),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_33),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_84),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_155),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_317),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_21),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_133),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_249),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_160),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_143),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_179),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_120),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_304),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_82),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_200),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_67),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_163),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_148),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_269),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_194),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_274),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_172),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_259),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_158),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_223),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_239),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_199),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_15),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_99),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_1),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_49),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_242),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_60),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_203),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_294),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_92),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_213),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_109),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_59),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_135),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_132),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_319),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_100),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_318),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_235),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_302),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_251),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_157),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_83),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_73),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_280),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_278),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_250),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_76),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_245),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_268),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_126),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_258),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_305),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_10),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_91),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_55),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_25),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_70),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_65),
.Y(n_471)
);

BUFx5_ASAP7_75t_L g472 ( 
.A(n_196),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_320),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_47),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_288),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_149),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_101),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_96),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_241),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_38),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_270),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_324),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_21),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_209),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_19),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_225),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_174),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_94),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_210),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_264),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_276),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_195),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_16),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_176),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_41),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_244),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_296),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_198),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_285),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_22),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_256),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_64),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_97),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_53),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_301),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_162),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_159),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_89),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_118),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_7),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_217),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_41),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_24),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_52),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_267),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_299),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_212),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_227),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_10),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_5),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_314),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_273),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_38),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_315),
.Y(n_524)
);

BUFx5_ASAP7_75t_L g525 ( 
.A(n_98),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_289),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_40),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_192),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_138),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_262),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_17),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_3),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_27),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_191),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_141),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_31),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_18),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_411),
.B(n_0),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_391),
.Y(n_539)
);

BUFx12f_ASAP7_75t_L g540 ( 
.A(n_355),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_344),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_429),
.B(n_1),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_429),
.B(n_515),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_344),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_344),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_329),
.B(n_2),
.Y(n_546)
);

BUFx8_ASAP7_75t_SL g547 ( 
.A(n_366),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_344),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_424),
.B(n_2),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_515),
.B(n_4),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_391),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_382),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_534),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_535),
.B(n_43),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_326),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_6),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_385),
.B(n_6),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_409),
.B(n_7),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_391),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_425),
.B(n_8),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_328),
.B(n_8),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_472),
.Y(n_563)
);

BUFx3_ASAP7_75t_L g564 ( 
.A(n_355),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_330),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_328),
.B(n_9),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_495),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_495),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_334),
.B(n_9),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_428),
.B(n_11),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_472),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_348),
.Y(n_572)
);

BUFx12f_ASAP7_75t_L g573 ( 
.A(n_364),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_509),
.B(n_11),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_534),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_334),
.B(n_12),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_369),
.Y(n_577)
);

INVx5_ASAP7_75t_L g578 ( 
.A(n_534),
.Y(n_578)
);

BUFx8_ASAP7_75t_L g579 ( 
.A(n_500),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_534),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_374),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

BUFx8_ASAP7_75t_L g583 ( 
.A(n_523),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_386),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_374),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_364),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_518),
.B(n_12),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_427),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_521),
.B(n_327),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_389),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_389),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_340),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_350),
.B(n_13),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_408),
.B(n_13),
.Y(n_595)
);

AND2x6_ASAP7_75t_L g596 ( 
.A(n_352),
.B(n_44),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_472),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_367),
.B(n_14),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_450),
.B(n_14),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_408),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_421),
.B(n_16),
.Y(n_601)
);

CKINVDCx6p67_ASAP7_75t_R g602 ( 
.A(n_421),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_434),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_480),
.B(n_18),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_336),
.Y(n_606)
);

BUFx8_ASAP7_75t_SL g607 ( 
.A(n_336),
.Y(n_607)
);

CKINVDCx11_ASAP7_75t_R g608 ( 
.A(n_360),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_485),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

BUFx12f_ASAP7_75t_L g611 ( 
.A(n_407),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_496),
.B(n_19),
.Y(n_612)
);

NOR2x1_ASAP7_75t_L g613 ( 
.A(n_338),
.B(n_45),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_342),
.B(n_388),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_476),
.B(n_20),
.Y(n_615)
);

INVx5_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_331),
.Y(n_617)
);

BUFx12f_ASAP7_75t_L g618 ( 
.A(n_436),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_472),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_466),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_332),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_476),
.B(n_20),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_525),
.B(n_22),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_513),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_525),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_347),
.Y(n_626)
);

NOR2x1_ASAP7_75t_L g627 ( 
.A(n_349),
.B(n_51),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_525),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_525),
.B(n_23),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_469),
.B(n_23),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_356),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_525),
.B(n_25),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_412),
.B(n_26),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_358),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_525),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_467),
.B(n_26),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_362),
.B(n_54),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_483),
.B(n_27),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_531),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

AND2x6_ASAP7_75t_L g642 ( 
.A(n_470),
.B(n_58),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_487),
.B(n_28),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_363),
.B(n_28),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_493),
.Y(n_645)
);

CKINVDCx6p67_ASAP7_75t_R g646 ( 
.A(n_346),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_510),
.B(n_29),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_533),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_365),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_368),
.B(n_29),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_536),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_512),
.B(n_30),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_520),
.B(n_527),
.Y(n_653)
);

BUFx12f_ASAP7_75t_L g654 ( 
.A(n_333),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_543),
.A2(n_537),
.B1(n_371),
.B2(n_378),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_572),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_548),
.Y(n_657)
);

AO22x2_ASAP7_75t_L g658 ( 
.A1(n_562),
.A2(n_380),
.B1(n_381),
.B2(n_370),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_552),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_542),
.A2(n_401),
.B1(n_403),
.B2(n_398),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_614),
.A2(n_418),
.B1(n_420),
.B2(n_417),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_539),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_556),
.B(n_383),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_617),
.B(n_501),
.Y(n_664)
);

AO22x2_ASAP7_75t_L g665 ( 
.A1(n_562),
.A2(n_392),
.B1(n_393),
.B2(n_387),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_R g666 ( 
.A1(n_577),
.A2(n_397),
.B1(n_402),
.B2(n_395),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_L g667 ( 
.A1(n_558),
.A2(n_497),
.B1(n_514),
.B2(n_494),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_550),
.A2(n_517),
.B1(n_529),
.B2(n_522),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_621),
.B(n_410),
.Y(n_669)
);

AO22x2_ASAP7_75t_L g670 ( 
.A1(n_566),
.A2(n_416),
.B1(n_426),
.B2(n_414),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_606),
.B(n_443),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_SL g672 ( 
.A1(n_601),
.A2(n_445),
.B1(n_455),
.B2(n_444),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_653),
.B(n_335),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_546),
.A2(n_339),
.B1(n_341),
.B2(n_337),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_539),
.Y(n_675)
);

XNOR2xp5_ASAP7_75t_L g676 ( 
.A(n_595),
.B(n_30),
.Y(n_676)
);

AO22x2_ASAP7_75t_L g677 ( 
.A1(n_566),
.A2(n_458),
.B1(n_460),
.B2(n_456),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_560),
.Y(n_678)
);

AO22x2_ASAP7_75t_L g679 ( 
.A1(n_576),
.A2(n_468),
.B1(n_474),
.B2(n_465),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_560),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_559),
.A2(n_345),
.B1(n_351),
.B2(n_343),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_565),
.B(n_484),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_633),
.A2(n_354),
.B1(n_357),
.B2(n_353),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_636),
.A2(n_361),
.B1(n_372),
.B2(n_359),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_545),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_581),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_586),
.B(n_486),
.Y(n_687)
);

AO22x2_ASAP7_75t_L g688 ( 
.A1(n_576),
.A2(n_489),
.B1(n_490),
.B2(n_491),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_586),
.B(n_373),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_586),
.B(n_592),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_607),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_551),
.A2(n_498),
.B1(n_503),
.B2(n_504),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_545),
.Y(n_693)
);

AO22x2_ASAP7_75t_L g694 ( 
.A1(n_538),
.A2(n_511),
.B1(n_32),
.B2(n_33),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_545),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_547),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_615),
.A2(n_530),
.B1(n_528),
.B2(n_526),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_554),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_569),
.B(n_375),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_554),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_592),
.B(n_376),
.Y(n_701)
);

AND2x2_ASAP7_75t_SL g702 ( 
.A(n_643),
.B(n_31),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_598),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_581),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_377),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_557),
.B(n_379),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_564),
.B(n_384),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_622),
.A2(n_620),
.B1(n_602),
.B2(n_570),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_600),
.A2(n_524),
.B1(n_516),
.B2(n_508),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_585),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_600),
.B(n_390),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_600),
.B(n_620),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_611),
.B(n_34),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_585),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_585),
.Y(n_716)
);

OA22x2_ASAP7_75t_L g717 ( 
.A1(n_567),
.A2(n_507),
.B1(n_506),
.B2(n_505),
.Y(n_717)
);

OA22x2_ASAP7_75t_L g718 ( 
.A1(n_568),
.A2(n_502),
.B1(n_499),
.B2(n_492),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_645),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_R g720 ( 
.A1(n_584),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_587),
.B(n_589),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_587),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_645),
.B(n_394),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_554),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_575),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_575),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_618),
.A2(n_442),
.B1(n_481),
.B2(n_479),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_630),
.A2(n_482),
.B1(n_477),
.B2(n_475),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_645),
.B(n_396),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_587),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_574),
.A2(n_473),
.B1(n_471),
.B2(n_464),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_575),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_589),
.B(n_399),
.Y(n_733)
);

XNOR2xp5_ASAP7_75t_L g734 ( 
.A(n_639),
.B(n_36),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_647),
.A2(n_652),
.B1(n_561),
.B2(n_573),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_589),
.B(n_400),
.Y(n_736)
);

BUFx10_ASAP7_75t_L g737 ( 
.A(n_603),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_540),
.A2(n_463),
.B1(n_462),
.B2(n_461),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_590),
.B(n_404),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_593),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_591),
.A2(n_459),
.B1(n_457),
.B2(n_454),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_580),
.Y(n_743)
);

OA22x2_ASAP7_75t_L g744 ( 
.A1(n_553),
.A2(n_453),
.B1(n_452),
.B2(n_451),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_685),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_661),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_721),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_722),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_696),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_663),
.B(n_682),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_693),
.Y(n_751)
);

AND2x2_ASAP7_75t_SL g752 ( 
.A(n_702),
.B(n_598),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_722),
.Y(n_753)
);

XOR2xp5_ASAP7_75t_L g754 ( 
.A(n_691),
.B(n_405),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_656),
.B(n_646),
.Y(n_755)
);

OAI21xp5_ASAP7_75t_L g756 ( 
.A1(n_717),
.A2(n_638),
.B(n_555),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_713),
.B(n_654),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_741),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_695),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_698),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_733),
.Y(n_761)
);

XOR2xp5_ASAP7_75t_L g762 ( 
.A(n_691),
.B(n_406),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_739),
.B(n_588),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_700),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_736),
.B(n_640),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_657),
.B(n_563),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_686),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_724),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_725),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_726),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_732),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_740),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_743),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_668),
.B(n_579),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_659),
.B(n_571),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_704),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_710),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_669),
.B(n_637),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_711),
.Y(n_779)
);

XOR2x2_ASAP7_75t_L g780 ( 
.A(n_676),
.B(n_608),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_664),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_SL g782 ( 
.A(n_667),
.B(n_642),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_715),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_662),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_718),
.A2(n_744),
.B(n_681),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_R g786 ( 
.A(n_707),
.B(n_413),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_683),
.B(n_579),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_684),
.B(n_583),
.Y(n_788)
);

XOR2xp5_ASAP7_75t_L g789 ( 
.A(n_727),
.B(n_415),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_690),
.B(n_609),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_716),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_673),
.B(n_609),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_730),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_675),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_678),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_674),
.A2(n_638),
.B(n_555),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_701),
.B(n_624),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_680),
.Y(n_798)
);

NOR2xp67_ASAP7_75t_L g799 ( 
.A(n_738),
.B(n_544),
.Y(n_799)
);

INVxp33_ASAP7_75t_L g800 ( 
.A(n_676),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_669),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_737),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_687),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_692),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_705),
.B(n_712),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_699),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_697),
.B(n_593),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_658),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_671),
.B(n_648),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_658),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_665),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_665),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_707),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_670),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_670),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_SL g816 ( 
.A(n_660),
.B(n_642),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_677),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_699),
.B(n_582),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_677),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_679),
.Y(n_820)
);

INVxp33_ASAP7_75t_L g821 ( 
.A(n_734),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_679),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_723),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_728),
.B(n_583),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_688),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_688),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_742),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_655),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_792),
.B(n_655),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_797),
.B(n_694),
.Y(n_830)
);

INVxp67_ASAP7_75t_SL g831 ( 
.A(n_801),
.Y(n_831)
);

AND2x4_ASAP7_75t_SL g832 ( 
.A(n_801),
.B(n_671),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_763),
.B(n_694),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_763),
.B(n_703),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_748),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_805),
.B(n_703),
.Y(n_837)
);

AND2x2_ASAP7_75t_SL g838 ( 
.A(n_752),
.B(n_623),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_781),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_766),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_753),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_766),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_750),
.B(n_729),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_784),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_775),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_775),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_794),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_749),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_780),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_818),
.B(n_734),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_828),
.B(n_708),
.Y(n_851)
);

BUFx6f_ASAP7_75t_L g852 ( 
.A(n_801),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_818),
.B(n_778),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_778),
.B(n_735),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_795),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_798),
.Y(n_856)
);

NOR2xp67_ASAP7_75t_L g857 ( 
.A(n_802),
.B(n_719),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_786),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_823),
.B(n_604),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_827),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_790),
.B(n_624),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_745),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_751),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_764),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_765),
.B(n_641),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_765),
.B(n_641),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_759),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_755),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_767),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_760),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_816),
.B(n_731),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_803),
.B(n_555),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_807),
.B(n_761),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_809),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_806),
.B(n_651),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_806),
.B(n_804),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_804),
.B(n_597),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_813),
.B(n_625),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_768),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_785),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_769),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_770),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_771),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_758),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_808),
.B(n_638),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_776),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_785),
.B(n_628),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_774),
.B(n_746),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_807),
.B(n_635),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_810),
.Y(n_890)
);

NAND2xp33_ASAP7_75t_L g891 ( 
.A(n_796),
.B(n_638),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_811),
.B(n_626),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_812),
.B(n_626),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_814),
.B(n_626),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_772),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_777),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_809),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_816),
.B(n_672),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_773),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_782),
.B(n_642),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_779),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_R g902 ( 
.A(n_782),
.B(n_706),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_815),
.B(n_817),
.Y(n_903)
);

INVx1_ASAP7_75t_SL g904 ( 
.A(n_757),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_783),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_791),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_756),
.B(n_593),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_793),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_756),
.B(n_605),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_819),
.B(n_631),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_831),
.B(n_826),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_903),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_843),
.B(n_842),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_832),
.Y(n_914)
);

NAND2x1p5_ASAP7_75t_L g915 ( 
.A(n_852),
.B(n_820),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_888),
.B(n_821),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_850),
.B(n_800),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_869),
.B(n_825),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_903),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_873),
.B(n_789),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_850),
.B(n_880),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_863),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_885),
.B(n_822),
.Y(n_923)
);

BUFx4f_ASAP7_75t_L g924 ( 
.A(n_832),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_863),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_876),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_864),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_864),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_876),
.Y(n_929)
);

OR2x2_ASAP7_75t_L g930 ( 
.A(n_880),
.B(n_754),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_842),
.B(n_796),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_840),
.Y(n_932)
);

CKINVDCx8_ASAP7_75t_R g933 ( 
.A(n_848),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_858),
.B(n_787),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_840),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_848),
.B(n_824),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_868),
.B(n_762),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_852),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_869),
.B(n_799),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_847),
.Y(n_940)
);

INVx4_ASAP7_75t_L g941 ( 
.A(n_852),
.Y(n_941)
);

BUFx12f_ASAP7_75t_L g942 ( 
.A(n_874),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_891),
.A2(n_549),
.B(n_544),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_889),
.B(n_788),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_845),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_889),
.B(n_709),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_903),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_869),
.B(n_714),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_845),
.B(n_605),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_874),
.Y(n_950)
);

OR2x6_ASAP7_75t_L g951 ( 
.A(n_837),
.B(n_714),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_852),
.Y(n_952)
);

AND2x2_ASAP7_75t_SL g953 ( 
.A(n_834),
.B(n_720),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_853),
.B(n_689),
.Y(n_954)
);

AND2x4_ASAP7_75t_L g955 ( 
.A(n_853),
.B(n_613),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_906),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_847),
.Y(n_957)
);

INVx2_ASAP7_75t_SL g958 ( 
.A(n_865),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_906),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_865),
.B(n_627),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_846),
.B(n_605),
.Y(n_961)
);

NOR2x1_ASAP7_75t_L g962 ( 
.A(n_900),
.B(n_644),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_846),
.B(n_650),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_858),
.B(n_419),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_852),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_877),
.B(n_594),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_875),
.B(n_631),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_892),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_877),
.B(n_599),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_908),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_965),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_942),
.Y(n_972)
);

BUFx5_ASAP7_75t_L g973 ( 
.A(n_970),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_914),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_965),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_917),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_921),
.B(n_860),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_933),
.Y(n_978)
);

BUFx12f_ASAP7_75t_L g979 ( 
.A(n_948),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_912),
.Y(n_980)
);

INVx5_ASAP7_75t_L g981 ( 
.A(n_923),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_916),
.B(n_860),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_924),
.Y(n_983)
);

CKINVDCx14_ASAP7_75t_R g984 ( 
.A(n_937),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_923),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_922),
.Y(n_986)
);

INVx3_ASAP7_75t_SL g987 ( 
.A(n_951),
.Y(n_987)
);

INVx4_ASAP7_75t_L g988 ( 
.A(n_941),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_925),
.Y(n_989)
);

INVx8_ASAP7_75t_L g990 ( 
.A(n_923),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_927),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_930),
.Y(n_992)
);

INVx1_ASAP7_75t_SL g993 ( 
.A(n_926),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_913),
.A2(n_834),
.B1(n_835),
.B2(n_871),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_926),
.Y(n_995)
);

INVx6_ASAP7_75t_L g996 ( 
.A(n_912),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_928),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_932),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_948),
.Y(n_999)
);

INVx1_ASAP7_75t_SL g1000 ( 
.A(n_929),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_932),
.B(n_887),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_920),
.B(n_875),
.Y(n_1002)
);

AND2x4_ASAP7_75t_L g1003 ( 
.A(n_958),
.B(n_968),
.Y(n_1003)
);

AO21x2_ASAP7_75t_L g1004 ( 
.A1(n_931),
.A2(n_891),
.B(n_872),
.Y(n_1004)
);

BUFx2_ASAP7_75t_SL g1005 ( 
.A(n_919),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_919),
.Y(n_1006)
);

BUFx10_ASAP7_75t_L g1007 ( 
.A(n_964),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_935),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_950),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_947),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_941),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_935),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_947),
.Y(n_1013)
);

CKINVDCx12_ASAP7_75t_R g1014 ( 
.A(n_951),
.Y(n_1014)
);

INVxp67_ASAP7_75t_L g1015 ( 
.A(n_968),
.Y(n_1015)
);

INVx5_ASAP7_75t_L g1016 ( 
.A(n_938),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_1002),
.A2(n_838),
.B1(n_934),
.B2(n_835),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_980),
.Y(n_1018)
);

CKINVDCx11_ASAP7_75t_R g1019 ( 
.A(n_972),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_994),
.A2(n_944),
.B1(n_929),
.B2(n_966),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_994),
.A2(n_969),
.B1(n_945),
.B2(n_946),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_998),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_976),
.A2(n_838),
.B1(n_953),
.B2(n_902),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_982),
.B(n_967),
.Y(n_1024)
);

OAI22xp33_ASAP7_75t_R g1025 ( 
.A1(n_982),
.A2(n_666),
.B1(n_849),
.B2(n_851),
.Y(n_1025)
);

NAND2x1p5_ASAP7_75t_L g1026 ( 
.A(n_981),
.B(n_897),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_999),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_977),
.A2(n_945),
.B1(n_963),
.B2(n_1001),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1001),
.A2(n_959),
.B1(n_956),
.B2(n_952),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_981),
.B(n_839),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_992),
.A2(n_936),
.B1(n_904),
.B2(n_836),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1008),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_995),
.A2(n_854),
.B1(n_898),
.B2(n_954),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_SL g1034 ( 
.A1(n_984),
.A2(n_854),
.B(n_837),
.Y(n_1034)
);

CKINVDCx20_ASAP7_75t_R g1035 ( 
.A(n_992),
.Y(n_1035)
);

CKINVDCx11_ASAP7_75t_R g1036 ( 
.A(n_987),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_993),
.A2(n_1000),
.B1(n_1012),
.B2(n_939),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_978),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_993),
.B(n_1000),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_995),
.A2(n_954),
.B1(n_955),
.B2(n_829),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_986),
.Y(n_1041)
);

BUFx10_ASAP7_75t_L g1042 ( 
.A(n_1003),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1003),
.B(n_861),
.Y(n_1043)
);

BUFx8_ASAP7_75t_L g1044 ( 
.A(n_979),
.Y(n_1044)
);

INVx6_ASAP7_75t_L g1045 ( 
.A(n_983),
.Y(n_1045)
);

OAI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_987),
.A2(n_841),
.B1(n_851),
.B2(n_833),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1015),
.B(n_829),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_989),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1007),
.A2(n_955),
.B1(n_962),
.B2(n_960),
.Y(n_1049)
);

INVx8_ASAP7_75t_L g1050 ( 
.A(n_990),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1007),
.A2(n_960),
.B1(n_830),
.B2(n_911),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_984),
.A2(n_830),
.B1(n_911),
.B2(n_918),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_1014),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_991),
.A2(n_918),
.B1(n_887),
.B2(n_878),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_980),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_974),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_1023),
.A2(n_1015),
.B1(n_939),
.B2(n_1009),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1022),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1021),
.A2(n_1004),
.B(n_961),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_1019),
.Y(n_1060)
);

OAI22xp33_ASAP7_75t_SL g1061 ( 
.A1(n_1024),
.A2(n_629),
.B1(n_632),
.B2(n_612),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1017),
.A2(n_1049),
.B1(n_1033),
.B2(n_1051),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1040),
.A2(n_915),
.B1(n_1006),
.B2(n_996),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_1039),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1032),
.Y(n_1065)
);

OAI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1034),
.A2(n_849),
.B1(n_1013),
.B2(n_1010),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1041),
.Y(n_1067)
);

OAI222xp33_ASAP7_75t_L g1068 ( 
.A1(n_1020),
.A2(n_970),
.B1(n_907),
.B2(n_909),
.C1(n_957),
.C2(n_940),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1052),
.A2(n_996),
.B1(n_1006),
.B2(n_1005),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1025),
.A2(n_886),
.B1(n_884),
.B2(n_901),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_SL g1071 ( 
.A1(n_1035),
.A2(n_1037),
.B1(n_1028),
.B2(n_1053),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_1046),
.A2(n_859),
.B(n_861),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1031),
.A2(n_886),
.B1(n_884),
.B2(n_901),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_SL g1074 ( 
.A1(n_1043),
.A2(n_866),
.B(n_859),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_SL g1075 ( 
.A1(n_1044),
.A2(n_981),
.B1(n_990),
.B2(n_985),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1027),
.A2(n_1036),
.B1(n_886),
.B2(n_884),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1056),
.A2(n_857),
.B1(n_866),
.B2(n_878),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_1045),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_1018),
.Y(n_1079)
);

OAI222xp33_ASAP7_75t_L g1080 ( 
.A1(n_1029),
.A2(n_949),
.B1(n_997),
.B2(n_981),
.C1(n_893),
.C2(n_910),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_1054),
.A2(n_884),
.B1(n_886),
.B2(n_905),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_SL g1082 ( 
.A1(n_1044),
.A2(n_990),
.B1(n_985),
.B2(n_973),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1048),
.A2(n_886),
.B1(n_884),
.B2(n_905),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1047),
.A2(n_856),
.B1(n_855),
.B2(n_908),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_SL g1085 ( 
.A1(n_1050),
.A2(n_973),
.B1(n_894),
.B2(n_910),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1026),
.A2(n_896),
.B(n_870),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1042),
.B(n_892),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1030),
.A2(n_996),
.B1(n_1006),
.B2(n_1013),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_1045),
.A2(n_1010),
.B1(n_980),
.B2(n_908),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1038),
.B(n_1010),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_1018),
.Y(n_1091)
);

OAI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1050),
.A2(n_882),
.B1(n_883),
.B2(n_988),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1042),
.A2(n_867),
.B1(n_879),
.B2(n_899),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1018),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1055),
.A2(n_894),
.B1(n_893),
.B2(n_844),
.Y(n_1095)
);

OAI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1055),
.A2(n_1011),
.B1(n_988),
.B2(n_883),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1071),
.A2(n_596),
.B1(n_881),
.B2(n_895),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1064),
.B(n_1055),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1070),
.A2(n_1066),
.B1(n_1077),
.B2(n_1073),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_SL g1100 ( 
.A1(n_1062),
.A2(n_973),
.B1(n_1011),
.B2(n_596),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1072),
.A2(n_596),
.B1(n_895),
.B2(n_881),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1061),
.A2(n_596),
.B1(n_899),
.B2(n_882),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1065),
.B(n_1004),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1076),
.A2(n_1016),
.B1(n_975),
.B2(n_971),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1057),
.A2(n_1063),
.B1(n_1086),
.B2(n_1085),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_SL g1106 ( 
.A1(n_1069),
.A2(n_973),
.B1(n_885),
.B2(n_432),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1085),
.A2(n_862),
.B1(n_885),
.B2(n_431),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1058),
.B(n_973),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1093),
.A2(n_862),
.B1(n_433),
.B2(n_435),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1087),
.A2(n_422),
.B1(n_448),
.B2(n_449),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1084),
.A2(n_423),
.B1(n_446),
.B2(n_441),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1081),
.A2(n_430),
.B1(n_440),
.B2(n_439),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_SL g1113 ( 
.A1(n_1090),
.A2(n_973),
.B1(n_438),
.B2(n_437),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1067),
.B(n_890),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1082),
.A2(n_1075),
.B1(n_1092),
.B2(n_1095),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1074),
.A2(n_447),
.B1(n_975),
.B2(n_971),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1075),
.A2(n_1016),
.B1(n_943),
.B2(n_649),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_1082),
.A2(n_649),
.B1(n_634),
.B2(n_631),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1059),
.Y(n_1119)
);

AOI22xp33_ASAP7_75t_L g1120 ( 
.A1(n_1088),
.A2(n_1083),
.B1(n_1089),
.B2(n_1091),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1079),
.A2(n_649),
.B1(n_634),
.B2(n_1016),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1078),
.A2(n_1016),
.B1(n_634),
.B2(n_610),
.Y(n_1122)
);

NAND3xp33_ASAP7_75t_L g1123 ( 
.A(n_1096),
.B(n_610),
.C(n_619),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1094),
.A2(n_619),
.B1(n_616),
.B2(n_541),
.Y(n_1124)
);

AOI221xp5_ASAP7_75t_SL g1125 ( 
.A1(n_1080),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.C(n_580),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1060),
.A2(n_619),
.B1(n_616),
.B2(n_541),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1080),
.A2(n_616),
.B1(n_610),
.B2(n_578),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1068),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1068),
.A2(n_578),
.B1(n_549),
.B2(n_544),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1064),
.B(n_39),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1071),
.A2(n_578),
.B1(n_549),
.B2(n_42),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1071),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1071),
.A2(n_79),
.B1(n_81),
.B2(n_85),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1098),
.B(n_1108),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1132),
.B(n_86),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1131),
.A2(n_87),
.B1(n_90),
.B2(n_93),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1108),
.B(n_95),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1099),
.A2(n_103),
.B1(n_106),
.B2(n_108),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1103),
.B(n_111),
.Y(n_1139)
);

OA21x2_ASAP7_75t_L g1140 ( 
.A1(n_1119),
.A2(n_112),
.B(n_113),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1103),
.B(n_114),
.Y(n_1141)
);

NOR3xp33_ASAP7_75t_L g1142 ( 
.A(n_1125),
.B(n_1113),
.C(n_1106),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1130),
.B(n_115),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1133),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1105),
.B(n_121),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1128),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1128),
.B(n_1114),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1120),
.B(n_323),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1119),
.B(n_122),
.Y(n_1149)
);

NAND4xp25_ASAP7_75t_L g1150 ( 
.A(n_1110),
.B(n_123),
.C(n_124),
.D(n_125),
.Y(n_1150)
);

NAND3xp33_ASAP7_75t_L g1151 ( 
.A(n_1102),
.B(n_127),
.C(n_129),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1115),
.B(n_1116),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1127),
.A2(n_130),
.B1(n_136),
.B2(n_137),
.C(n_139),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_L g1154 ( 
.A(n_1100),
.B(n_142),
.C(n_144),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_L g1155 ( 
.A(n_1126),
.B(n_1111),
.C(n_1097),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1107),
.B(n_147),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1104),
.B(n_150),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1112),
.B(n_152),
.C(n_161),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1147),
.B(n_1134),
.Y(n_1159)
);

AO21x2_ASAP7_75t_L g1160 ( 
.A1(n_1146),
.A2(n_1123),
.B(n_1117),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1139),
.B(n_1129),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1141),
.B(n_1118),
.Y(n_1162)
);

NAND3xp33_ASAP7_75t_L g1163 ( 
.A(n_1142),
.B(n_1101),
.C(n_1109),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_SL g1164 ( 
.A(n_1150),
.B(n_1122),
.Y(n_1164)
);

NOR3xp33_ASAP7_75t_L g1165 ( 
.A(n_1152),
.B(n_1121),
.C(n_1124),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1149),
.A2(n_165),
.B(n_167),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1140),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_1137),
.B(n_168),
.Y(n_1168)
);

NOR3xp33_ASAP7_75t_L g1169 ( 
.A(n_1142),
.B(n_173),
.C(n_175),
.Y(n_1169)
);

AO21x2_ASAP7_75t_L g1170 ( 
.A1(n_1154),
.A2(n_177),
.B(n_181),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1159),
.B(n_1167),
.Y(n_1171)
);

NAND4xp75_ASAP7_75t_L g1172 ( 
.A(n_1162),
.B(n_1145),
.C(n_1148),
.D(n_1153),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1168),
.B(n_1140),
.Y(n_1173)
);

NAND4xp75_ASAP7_75t_L g1174 ( 
.A(n_1169),
.B(n_1143),
.C(n_1157),
.D(n_1156),
.Y(n_1174)
);

AND4x1_ASAP7_75t_L g1175 ( 
.A(n_1164),
.B(n_1135),
.C(n_1138),
.D(n_1155),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1160),
.Y(n_1176)
);

NAND4xp75_ASAP7_75t_SL g1177 ( 
.A(n_1170),
.B(n_1154),
.C(n_1151),
.D(n_1158),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1161),
.B(n_1136),
.Y(n_1178)
);

XOR2x2_ASAP7_75t_L g1179 ( 
.A(n_1163),
.B(n_1144),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1160),
.B(n_183),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1176),
.Y(n_1181)
);

XNOR2xp5_ASAP7_75t_L g1182 ( 
.A(n_1179),
.B(n_1163),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1171),
.Y(n_1183)
);

OA22x2_ASAP7_75t_L g1184 ( 
.A1(n_1173),
.A2(n_1168),
.B1(n_1170),
.B2(n_1165),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1178),
.B(n_1166),
.Y(n_1185)
);

INVx1_ASAP7_75t_SL g1186 ( 
.A(n_1180),
.Y(n_1186)
);

XNOR2xp5_ASAP7_75t_L g1187 ( 
.A(n_1175),
.B(n_1166),
.Y(n_1187)
);

AOI22x1_ASAP7_75t_L g1188 ( 
.A1(n_1187),
.A2(n_1177),
.B1(n_1175),
.B2(n_1174),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1183),
.Y(n_1189)
);

OA22x2_ASAP7_75t_L g1190 ( 
.A1(n_1182),
.A2(n_1172),
.B1(n_185),
.B2(n_186),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1187),
.Y(n_1191)
);

AOI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1185),
.A2(n_184),
.B1(n_190),
.B2(n_193),
.Y(n_1192)
);

AOI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1184),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_1193)
);

OA22x2_ASAP7_75t_L g1194 ( 
.A1(n_1186),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_1181),
.Y(n_1195)
);

OAI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1187),
.A2(n_214),
.B1(n_215),
.B2(n_218),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1183),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1189),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1197),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1188),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1195),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1191),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1194),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1200),
.A2(n_1193),
.B1(n_1190),
.B2(n_1196),
.Y(n_1204)
);

OA22x2_ASAP7_75t_L g1205 ( 
.A1(n_1202),
.A2(n_1188),
.B1(n_1192),
.B2(n_224),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1203),
.A2(n_1201),
.B1(n_1198),
.B2(n_1199),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1199),
.A2(n_221),
.B1(n_222),
.B2(n_226),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1200),
.A2(n_228),
.B(n_229),
.C(n_230),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1199),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1209),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1204),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1205),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1206),
.Y(n_1213)
);

AO22x2_ASAP7_75t_L g1214 ( 
.A1(n_1213),
.A2(n_1207),
.B1(n_1208),
.B2(n_237),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1212),
.B(n_234),
.Y(n_1215)
);

OA22x2_ASAP7_75t_L g1216 ( 
.A1(n_1211),
.A2(n_236),
.B1(n_238),
.B2(n_240),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1215),
.Y(n_1217)
);

XOR2xp5_ASAP7_75t_L g1218 ( 
.A(n_1214),
.B(n_1210),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1216),
.Y(n_1219)
);

AOI21xp33_ASAP7_75t_L g1220 ( 
.A1(n_1217),
.A2(n_322),
.B(n_246),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_1219),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1221),
.Y(n_1222)
);

AO22x2_ASAP7_75t_L g1223 ( 
.A1(n_1222),
.A2(n_1218),
.B1(n_1220),
.B2(n_253),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1222),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1224),
.Y(n_1225)
);

INVx2_ASAP7_75t_SL g1226 ( 
.A(n_1223),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1226),
.A2(n_243),
.B1(n_247),
.B2(n_255),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1225),
.A2(n_257),
.B1(n_261),
.B2(n_263),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1226),
.A2(n_271),
.B1(n_275),
.B2(n_283),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1229),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1230),
.A2(n_1227),
.B1(n_1228),
.B2(n_293),
.Y(n_1231)
);

INVxp67_ASAP7_75t_L g1232 ( 
.A(n_1231),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1232),
.A2(n_284),
.B1(n_292),
.B2(n_295),
.C(n_297),
.Y(n_1233)
);

AOI211xp5_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_298),
.B(n_300),
.C(n_303),
.Y(n_1234)
);


endmodule