module fake_jpeg_14286_n_644 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_644);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_644;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_2),
.B(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_9),
.B(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_28),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_62),
.B(n_65),
.Y(n_132)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_67),
.Y(n_187)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_68),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_69),
.B(n_72),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_70),
.Y(n_189)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_71),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_18),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_74),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_78),
.B(n_84),
.Y(n_175)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_79),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_80),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_81),
.Y(n_193)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_83),
.Y(n_216)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_50),
.Y(n_86)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_89),
.B(n_90),
.Y(n_177)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

CKINVDCx11_ASAP7_75t_R g91 ( 
.A(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_91),
.B(n_99),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_94),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_95),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_38),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_96),
.Y(n_166)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_29),
.Y(n_97)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_98),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_57),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_101),
.B(n_103),
.Y(n_213)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_38),
.Y(n_102)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_36),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_44),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_104),
.B(n_106),
.Y(n_215)
);

BUFx4f_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_32),
.Y(n_108)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_109),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_110),
.Y(n_180)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_44),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_112),
.B(n_115),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_24),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_114),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_40),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_116),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_33),
.Y(n_117)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_40),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_129),
.Y(n_147)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_123),
.Y(n_212)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_124),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_34),
.Y(n_125)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_61),
.B(n_14),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_127),
.B(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_49),
.Y(n_128)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_128),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_49),
.Y(n_130)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_130),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_141),
.B(n_110),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_71),
.B(n_55),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_149),
.B(n_172),
.Y(n_219)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_73),
.A2(n_34),
.B1(n_46),
.B2(n_19),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_151),
.A2(n_195),
.B1(n_86),
.B2(n_126),
.Y(n_226)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_60),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_155),
.B(n_96),
.C(n_118),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_74),
.A2(n_55),
.B1(n_60),
.B2(n_46),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_156),
.A2(n_168),
.B1(n_111),
.B2(n_110),
.Y(n_253)
);

BUFx8_ASAP7_75t_L g162 ( 
.A(n_102),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g249 ( 
.A(n_162),
.Y(n_249)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_58),
.B(n_51),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_163),
.B(n_87),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_63),
.A2(n_46),
.B1(n_24),
.B2(n_53),
.Y(n_168)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_170),
.Y(n_271)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_20),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_77),
.B(n_21),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_173),
.B(n_194),
.Y(n_241)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_80),
.Y(n_178)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_178),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_179),
.B(n_14),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_82),
.B(n_20),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_214),
.Y(n_228)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_76),
.Y(n_182)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_67),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_183),
.Y(n_218)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_88),
.B(n_21),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_97),
.A2(n_19),
.B1(n_53),
.B2(n_58),
.Y(n_195)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_105),
.Y(n_205)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_205),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_122),
.A2(n_19),
.B1(n_53),
.B2(n_39),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_207),
.A2(n_81),
.B1(n_98),
.B2(n_95),
.Y(n_263)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_105),
.Y(n_210)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_210),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_94),
.B(n_39),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_217),
.B(n_280),
.Y(n_322)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_220),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_221),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_155),
.A2(n_116),
.B(n_85),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_223),
.A2(n_188),
.B(n_135),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_100),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_225),
.B(n_230),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_226),
.A2(n_254),
.B1(n_267),
.B2(n_208),
.Y(n_293)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

CKINVDCx12_ASAP7_75t_R g229 ( 
.A(n_176),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_229),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_120),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_231),
.B(n_243),
.Y(n_320)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_232),
.Y(n_341)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_140),
.Y(n_233)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_233),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_237),
.B(n_270),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_238),
.Y(n_351)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_240),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_132),
.B(n_22),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_244),
.B(n_259),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_56),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_245),
.B(n_247),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_56),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_153),
.Y(n_248)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_248),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_147),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_250),
.B(n_252),
.Y(n_326)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_144),
.Y(n_251)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_251),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_132),
.B(n_51),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_253),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_151),
.A2(n_125),
.B1(n_123),
.B2(n_83),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_145),
.Y(n_256)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_143),
.A2(n_109),
.B1(n_54),
.B2(n_113),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_263),
.B1(n_143),
.B2(n_159),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_137),
.B(n_37),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_177),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_260),
.B(n_266),
.Y(n_343)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_169),
.Y(n_262)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_168),
.A2(n_93),
.B1(n_92),
.B2(n_70),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_264),
.A2(n_279),
.B1(n_281),
.B2(n_161),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_137),
.B(n_45),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_173),
.A2(n_45),
.B1(n_37),
.B2(n_27),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_193),
.Y(n_268)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_268),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_269),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_211),
.B(n_54),
.Y(n_270)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_160),
.Y(n_272)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_272),
.Y(n_329)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_164),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_193),
.Y(n_274)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_274),
.Y(n_337)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_162),
.Y(n_275)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_275),
.Y(n_316)
);

CKINVDCx12_ASAP7_75t_R g276 ( 
.A(n_135),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_276),
.B(n_277),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_194),
.B(n_27),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_175),
.B(n_179),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_282),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_156),
.A2(n_117),
.B1(n_22),
.B2(n_85),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_157),
.B(n_117),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_163),
.A2(n_197),
.B1(n_203),
.B2(n_191),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_175),
.B(n_0),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_174),
.B(n_0),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_285),
.Y(n_328)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_204),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_166),
.B(n_2),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_166),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_286),
.B(n_289),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_148),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_136),
.B(n_3),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_167),
.A2(n_87),
.B(n_4),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_185),
.C(n_200),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_192),
.Y(n_292)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_292),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_293),
.A2(n_315),
.B1(n_269),
.B2(n_265),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_294),
.A2(n_321),
.B1(n_336),
.B2(n_242),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g301 ( 
.A(n_217),
.B(n_158),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_301),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_228),
.A2(n_165),
.B1(n_199),
.B2(n_131),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_303),
.A2(n_317),
.B1(n_318),
.B2(n_334),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_306),
.A2(n_325),
.B(n_330),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_263),
.A2(n_191),
.B1(n_212),
.B2(n_206),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_241),
.A2(n_146),
.B1(n_202),
.B2(n_196),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_253),
.A2(n_154),
.B1(n_216),
.B2(n_138),
.Y(n_321)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_288),
.A2(n_200),
.B(n_136),
.C(n_161),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_L g389 ( 
.A1(n_323),
.A2(n_269),
.B(n_249),
.C(n_238),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_219),
.B(n_188),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_331),
.B(n_272),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_258),
.A2(n_139),
.B1(n_180),
.B2(n_152),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_288),
.A2(n_201),
.B1(n_133),
.B2(n_6),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_3),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_339),
.B(n_342),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_5),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_254),
.A2(n_201),
.B1(n_8),
.B2(n_11),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_347),
.A2(n_349),
.B1(n_224),
.B2(n_271),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_271),
.B(n_7),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_348),
.B(n_249),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_223),
.A2(n_7),
.B1(n_11),
.B2(n_12),
.Y(n_349)
);

OA22x2_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_11),
.B1(n_12),
.B2(n_284),
.Y(n_350)
);

AND2x2_ASAP7_75t_SL g360 ( 
.A(n_350),
.B(n_12),
.Y(n_360)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_227),
.Y(n_352)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_352),
.Y(n_356)
);

INVx13_ASAP7_75t_L g353 ( 
.A(n_351),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_346),
.A2(n_246),
.B(n_224),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_354),
.A2(n_376),
.B(n_335),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_293),
.A2(n_232),
.B1(n_240),
.B2(n_233),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_355),
.A2(n_379),
.B1(n_381),
.B2(n_387),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_357),
.B(n_361),
.Y(n_419)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_344),
.Y(n_359)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_383),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_320),
.B(n_222),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_273),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_368),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_364),
.B(n_349),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_298),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_365),
.A2(n_296),
.B(n_302),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_301),
.B(n_251),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_369),
.B(n_377),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_317),
.A2(n_220),
.B1(n_218),
.B2(n_239),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_370),
.A2(n_391),
.B1(n_392),
.B2(n_335),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_340),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_384),
.Y(n_412)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_373),
.Y(n_428)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_374),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_307),
.B(n_292),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_380),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_346),
.A2(n_246),
.B(n_275),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_301),
.B(n_239),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_300),
.Y(n_378)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_378),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_315),
.A2(n_291),
.B1(n_274),
.B2(n_234),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_222),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_306),
.A2(n_268),
.B1(n_218),
.B2(n_255),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_255),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_350),
.Y(n_415)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_313),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_314),
.B(n_236),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_385),
.B(n_398),
.Y(n_405)
);

INVx4_ASAP7_75t_SL g386 ( 
.A(n_323),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_386),
.Y(n_425)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_390),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g399 ( 
.A1(n_389),
.A2(n_395),
.B(n_325),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_324),
.B(n_287),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_305),
.Y(n_391)
);

BUFx12f_ASAP7_75t_L g392 ( 
.A(n_304),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_295),
.B(n_287),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_319),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_265),
.B1(n_256),
.B2(n_236),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_394),
.A2(n_347),
.B1(n_325),
.B2(n_333),
.Y(n_409)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_396),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_322),
.A2(n_12),
.B1(n_261),
.B2(n_318),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_397),
.A2(n_342),
.B1(n_316),
.B2(n_327),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_343),
.B(n_261),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_371),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_322),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_400),
.B(n_420),
.C(n_362),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_401),
.A2(n_404),
.B1(n_430),
.B2(n_394),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_367),
.A2(n_322),
.B1(n_350),
.B2(n_330),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_409),
.A2(n_431),
.B1(n_359),
.B2(n_358),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_411),
.A2(n_429),
.B(n_386),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_422),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_415),
.B(n_424),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_371),
.A2(n_311),
.B(n_350),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_417),
.A2(n_381),
.B(n_362),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_418),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_364),
.B(n_326),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_366),
.B(n_297),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_365),
.Y(n_423)
);

INVx13_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_369),
.B(n_311),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_427),
.A2(n_386),
.B(n_389),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_377),
.A2(n_309),
.B(n_308),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_367),
.A2(n_341),
.B1(n_338),
.B2(n_337),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_355),
.A2(n_341),
.B1(n_305),
.B2(n_332),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_329),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_433),
.B(n_356),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_375),
.Y(n_434)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_434),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_363),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_436),
.B(n_373),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_437),
.B(n_384),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_415),
.A2(n_395),
.B1(n_397),
.B2(n_368),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_438),
.B(n_443),
.Y(n_482)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_407),
.Y(n_440)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_440),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_430),
.Y(n_491)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_407),
.Y(n_442)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_442),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_406),
.A2(n_354),
.B1(n_376),
.B2(n_372),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_412),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_444),
.B(n_446),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_445),
.A2(n_461),
.B(n_471),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_406),
.A2(n_360),
.B1(n_361),
.B2(n_379),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_447),
.B(n_465),
.Y(n_495)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_448),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_449),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_409),
.A2(n_385),
.B1(n_360),
.B2(n_357),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_450),
.A2(n_452),
.B1(n_405),
.B2(n_419),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_434),
.B(n_360),
.Y(n_451)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_453),
.B(n_422),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_454),
.A2(n_429),
.B(n_421),
.Y(n_480)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_426),
.Y(n_455)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_455),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_420),
.B(n_356),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_464),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_457),
.Y(n_486)
);

BUFx12_ASAP7_75t_L g458 ( 
.A(n_408),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_458),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_462),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g464 ( 
.A(n_419),
.B(n_383),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_403),
.A2(n_391),
.B1(n_337),
.B2(n_332),
.Y(n_465)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_426),
.Y(n_467)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_467),
.Y(n_505)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_416),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_468),
.Y(n_475)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_428),
.Y(n_469)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_469),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g471 ( 
.A1(n_425),
.A2(n_378),
.B(n_374),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_402),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_472),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_400),
.B(n_329),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_424),
.C(n_414),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_452),
.A2(n_403),
.B1(n_417),
.B2(n_425),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_477),
.A2(n_499),
.B1(n_438),
.B2(n_447),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g526 ( 
.A1(n_480),
.A2(n_470),
.B(n_463),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_483),
.B(n_485),
.C(n_501),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_458),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_484),
.B(n_498),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_491),
.B(n_465),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_448),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_460),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_413),
.C(n_405),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_458),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_410),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_413),
.C(n_404),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_503),
.B(n_416),
.C(n_391),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_461),
.A2(n_411),
.B(n_421),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_504),
.A2(n_506),
.B(n_445),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_457),
.A2(n_421),
.B(n_408),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_439),
.A2(n_435),
.B1(n_431),
.B2(n_410),
.Y(n_507)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_507),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_481),
.B(n_449),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g542 ( 
.A(n_509),
.B(n_511),
.Y(n_542)
);

XOR2x1_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_439),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_518),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_478),
.B(n_500),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_485),
.B(n_445),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_512),
.B(n_516),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_513),
.B(n_491),
.Y(n_550)
);

OA21x2_ASAP7_75t_SL g514 ( 
.A1(n_500),
.A2(n_459),
.B(n_451),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_514),
.B(n_525),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_483),
.B(n_459),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_517),
.A2(n_528),
.B1(n_495),
.B2(n_482),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_501),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g519 ( 
.A1(n_478),
.A2(n_463),
.B1(n_454),
.B2(n_467),
.Y(n_519)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_519),
.Y(n_547)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_520),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_521),
.A2(n_529),
.B(n_506),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_490),
.B(n_464),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_522),
.B(n_526),
.Y(n_562)
);

AOI211xp5_ASAP7_75t_SL g524 ( 
.A1(n_486),
.A2(n_443),
.B(n_470),
.C(n_460),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_524),
.B(n_505),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_474),
.B(n_455),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_476),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_531),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_495),
.A2(n_471),
.B1(n_401),
.B2(n_442),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_489),
.A2(n_471),
.B(n_440),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_488),
.Y(n_530)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_530),
.Y(n_554)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_476),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_493),
.B(n_427),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_535),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_432),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_536),
.C(n_537),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g535 ( 
.A(n_493),
.B(n_432),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_428),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_538),
.A2(n_544),
.B1(n_548),
.B2(n_561),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_484),
.C(n_502),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_541),
.B(n_543),
.C(n_557),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_474),
.C(n_486),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_517),
.A2(n_497),
.B1(n_487),
.B2(n_504),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_515),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_546),
.B(n_549),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_523),
.A2(n_497),
.B1(n_487),
.B2(n_496),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_522),
.B(n_488),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_550),
.B(n_468),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_513),
.A2(n_491),
.B1(n_489),
.B2(n_492),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_551),
.A2(n_556),
.B1(n_529),
.B2(n_524),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_553),
.A2(n_558),
.B(n_544),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_508),
.A2(n_492),
.B1(n_494),
.B2(n_505),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_475),
.C(n_479),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_528),
.A2(n_479),
.B1(n_494),
.B2(n_475),
.Y(n_561)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_545),
.Y(n_565)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_565),
.Y(n_597)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_552),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_566),
.B(n_568),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g601 ( 
.A(n_567),
.B(n_574),
.Y(n_601)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_554),
.Y(n_568)
);

BUFx12_ASAP7_75t_L g569 ( 
.A(n_541),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_569),
.Y(n_593)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_556),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_575),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_557),
.B(n_534),
.C(n_516),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_572),
.B(n_543),
.C(n_539),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_558),
.A2(n_521),
.B(n_536),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_573),
.A2(n_580),
.B(n_582),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_512),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_561),
.B(n_535),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_542),
.B(n_532),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_576),
.B(n_559),
.Y(n_590)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_554),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_578),
.Y(n_589)
);

INVx13_ASAP7_75t_L g578 ( 
.A(n_548),
.Y(n_578)
);

FAx1_ASAP7_75t_SL g579 ( 
.A(n_555),
.B(n_510),
.CI(n_533),
.CON(n_579),
.SN(n_579)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_579),
.B(n_581),
.Y(n_600)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_550),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_553),
.A2(n_388),
.B(n_396),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_583),
.A2(n_396),
.B(n_353),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_584),
.B(n_590),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_SL g586 ( 
.A(n_574),
.B(n_539),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_598),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_564),
.B(n_540),
.C(n_547),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_588),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_564),
.B(n_540),
.C(n_560),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g591 ( 
.A1(n_573),
.A2(n_551),
.B(n_562),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_592),
.Y(n_604)
);

XOR2x1_ASAP7_75t_SL g592 ( 
.A(n_575),
.B(n_538),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g594 ( 
.A(n_565),
.B(n_562),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_594),
.B(n_579),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_595),
.B(n_583),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_572),
.B(n_319),
.C(n_308),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_589),
.A2(n_566),
.B1(n_571),
.B2(n_581),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_603),
.A2(n_605),
.B1(n_611),
.B2(n_614),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_599),
.A2(n_571),
.B1(n_582),
.B2(n_580),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_597),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_606),
.B(n_609),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_610),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_597),
.Y(n_611)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_588),
.B(n_563),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_613),
.Y(n_623)
);

XOR2xp5_ASAP7_75t_L g613 ( 
.A(n_601),
.B(n_569),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_599),
.A2(n_578),
.B1(n_568),
.B2(n_569),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_579),
.C(n_312),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_615),
.B(n_598),
.Y(n_617)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_617),
.Y(n_631)
);

FAx1_ASAP7_75t_SL g618 ( 
.A(n_604),
.B(n_596),
.CI(n_587),
.CON(n_618),
.SN(n_618)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_618),
.B(n_619),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_608),
.B(n_584),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_600),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_620),
.B(n_621),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_585),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_SL g622 ( 
.A1(n_615),
.A2(n_592),
.B1(n_601),
.B2(n_591),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_622),
.B(n_596),
.C(n_609),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_602),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_626),
.B(n_586),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g627 ( 
.A1(n_623),
.A2(n_613),
.B(n_604),
.Y(n_627)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_627),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_628),
.B(n_629),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_616),
.A2(n_611),
.B(n_595),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_632),
.A2(n_621),
.B(n_617),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_SL g635 ( 
.A1(n_633),
.A2(n_624),
.B(n_625),
.C(n_618),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_635),
.A2(n_636),
.B(n_632),
.Y(n_638)
);

O2A1O1Ixp33_ASAP7_75t_SL g640 ( 
.A1(n_638),
.A2(n_639),
.B(n_634),
.C(n_353),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_637),
.B(n_630),
.C(n_631),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g641 ( 
.A(n_640),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_641),
.A2(n_392),
.B(n_304),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_392),
.B(n_351),
.Y(n_643)
);

FAx1_ASAP7_75t_SL g644 ( 
.A(n_643),
.B(n_392),
.CI(n_312),
.CON(n_644),
.SN(n_644)
);


endmodule