module fake_jpeg_22949_n_182 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_182);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_51),
.B(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_33),
.B1(n_22),
.B2(n_23),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_69),
.B(n_17),
.C(n_30),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_33),
.B1(n_35),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_61),
.A2(n_71),
.B1(n_34),
.B2(n_25),
.Y(n_96)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_29),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_44),
.A2(n_24),
.B1(n_30),
.B2(n_26),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_44),
.A2(n_35),
.B1(n_17),
.B2(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_77),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_42),
.B1(n_39),
.B2(n_37),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_113)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_78),
.B(n_83),
.Y(n_115)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_37),
.C(n_39),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_80),
.B(n_90),
.C(n_60),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_81),
.A2(n_84),
.B(n_31),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_54),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_89),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_43),
.C(n_40),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_48),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_27),
.B1(n_18),
.B2(n_26),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_95),
.B1(n_58),
.B2(n_52),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_43),
.B1(n_40),
.B2(n_29),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_20),
.B1(n_27),
.B2(n_25),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_20),
.B1(n_34),
.B2(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_102),
.B(n_117),
.Y(n_134)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_104),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_107),
.B1(n_119),
.B2(n_5),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_108),
.C(n_114),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_80),
.C(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_65),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_0),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_52),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_81),
.A2(n_66),
.B(n_48),
.C(n_49),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_118),
.A2(n_79),
.B1(n_99),
.B2(n_93),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_73),
.A2(n_63),
.B1(n_49),
.B2(n_4),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_84),
.B(n_13),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_31),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_118),
.B(n_109),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_127),
.B(n_130),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_75),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_136),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_88),
.C(n_85),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_133),
.C(n_138),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_135),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_1),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_12),
.C(n_11),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_1),
.Y(n_136)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_2),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_120),
.A3(n_114),
.B1(n_115),
.B2(n_118),
.C1(n_5),
.C2(n_10),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_11),
.C(n_6),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_139),
.A2(n_113),
.B1(n_116),
.B2(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_130),
.B(n_9),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_146),
.A2(n_147),
.B(n_137),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_115),
.B(n_118),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_149),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_111),
.B(n_9),
.C(n_10),
.D(n_7),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_138),
.C(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_7),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_7),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_158),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_160),
.Y(n_165)
);

OAI321xp33_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_143),
.A3(n_150),
.B1(n_151),
.B2(n_148),
.C(n_140),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_125),
.C(n_128),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_125),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_129),
.C(n_144),
.Y(n_168)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_163),
.Y(n_166)
);

OA21x2_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_143),
.B(n_159),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_160),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_168),
.C(n_156),
.Y(n_171)
);

OAI31xp33_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_173),
.A3(n_162),
.B(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_167),
.C(n_168),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_157),
.Y(n_172)
);

AOI31xp67_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_147),
.A3(n_159),
.B(n_127),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_174),
.A2(n_173),
.B(n_172),
.C(n_169),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_176),
.B(n_175),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_144),
.B(n_9),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_180),
.A2(n_179),
.B(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_181),
.Y(n_182)
);


endmodule