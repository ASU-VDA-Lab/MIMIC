module real_aes_7159_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g179 ( .A1(n_0), .A2(n_180), .B(n_183), .C(n_187), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_1), .B(n_171), .Y(n_190) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_3), .B(n_181), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_4), .A2(n_144), .B(n_147), .C(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_5), .A2(n_139), .B(n_550), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_6), .A2(n_139), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_7), .B(n_171), .Y(n_556) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_8), .A2(n_173), .B(n_245), .Y(n_244) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_9), .A2(n_460), .B1(n_747), .B2(n_748), .C1(n_751), .C2(n_754), .Y(n_459) );
AND2x6_ASAP7_75t_L g144 ( .A(n_10), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_11), .A2(n_144), .B(n_147), .C(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g516 ( .A(n_12), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_13), .B(n_41), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_13), .B(n_41), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_14), .B(n_186), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g101 ( .A1(n_15), .A2(n_102), .B1(n_115), .B2(n_758), .Y(n_101) );
INVx1_ASAP7_75t_L g165 ( .A(n_16), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_17), .B(n_181), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g455 ( .A(n_18), .B(n_456), .Y(n_455) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_19), .A2(n_182), .B(n_536), .C(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_20), .B(n_171), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_21), .B(n_159), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_22), .A2(n_147), .B(n_150), .C(n_158), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_23), .A2(n_185), .B(n_253), .C(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_24), .B(n_186), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_25), .B(n_186), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_26), .Y(n_497) );
INVx1_ASAP7_75t_L g477 ( .A(n_27), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_28), .A2(n_147), .B(n_158), .C(n_248), .Y(n_247) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_29), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_30), .Y(n_523) );
INVx1_ASAP7_75t_L g491 ( .A(n_31), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_32), .A2(n_139), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g142 ( .A(n_33), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_34), .A2(n_197), .B(n_198), .C(n_202), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_35), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_36), .A2(n_185), .B(n_553), .C(n_555), .Y(n_552) );
INVxp67_ASAP7_75t_L g492 ( .A(n_37), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_38), .B(n_250), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_39), .A2(n_147), .B(n_158), .C(n_476), .Y(n_475) );
CKINVDCx14_ASAP7_75t_R g551 ( .A(n_40), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_42), .A2(n_187), .B(n_514), .C(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_43), .B(n_138), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_44), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_45), .B(n_181), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_46), .B(n_139), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_47), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_48), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_49), .A2(n_197), .B(n_202), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g184 ( .A(n_50), .Y(n_184) );
INVx1_ASAP7_75t_L g228 ( .A(n_51), .Y(n_228) );
INVx1_ASAP7_75t_L g564 ( .A(n_52), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_53), .B(n_139), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_54), .Y(n_167) );
CKINVDCx14_ASAP7_75t_R g512 ( .A(n_55), .Y(n_512) );
INVx1_ASAP7_75t_L g145 ( .A(n_56), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_57), .B(n_139), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_58), .B(n_171), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_59), .A2(n_157), .B(n_213), .C(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g164 ( .A(n_60), .Y(n_164) );
INVx1_ASAP7_75t_SL g554 ( .A(n_61), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_62), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_63), .B(n_181), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_64), .B(n_171), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_65), .B(n_182), .Y(n_263) );
INVx1_ASAP7_75t_L g500 ( .A(n_66), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g177 ( .A(n_67), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_68), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g210 ( .A1(n_69), .A2(n_147), .B(n_202), .C(n_211), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_70), .Y(n_237) );
INVx1_ASAP7_75t_L g114 ( .A(n_71), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_72), .A2(n_139), .B(n_511), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g123 ( .A1(n_73), .A2(n_93), .B1(n_124), .B2(n_125), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_73), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_74), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_75), .A2(n_139), .B(n_533), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_76), .A2(n_100), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_76), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_77), .A2(n_138), .B(n_487), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g474 ( .A(n_78), .Y(n_474) );
INVx1_ASAP7_75t_L g534 ( .A(n_79), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_80), .B(n_155), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_81), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_82), .A2(n_139), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g537 ( .A(n_83), .Y(n_537) );
INVx2_ASAP7_75t_L g162 ( .A(n_84), .Y(n_162) );
INVx1_ASAP7_75t_L g526 ( .A(n_85), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_86), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_87), .B(n_186), .Y(n_264) );
INVx2_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
OR2x2_ASAP7_75t_L g451 ( .A(n_88), .B(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g463 ( .A(n_88), .B(n_453), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_89), .A2(n_147), .B(n_202), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_90), .B(n_139), .Y(n_195) );
INVx1_ASAP7_75t_L g199 ( .A(n_91), .Y(n_199) );
INVxp67_ASAP7_75t_L g240 ( .A(n_92), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_93), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_94), .B(n_173), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_95), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g212 ( .A(n_96), .Y(n_212) );
INVx1_ASAP7_75t_L g259 ( .A(n_97), .Y(n_259) );
INVx2_ASAP7_75t_L g567 ( .A(n_98), .Y(n_567) );
AND2x2_ASAP7_75t_L g230 ( .A(n_99), .B(n_161), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_100), .Y(n_749) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g758 ( .A(n_104), .Y(n_758) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g453 ( .A(n_110), .B(n_454), .Y(n_453) );
OR2x2_ASAP7_75t_L g466 ( .A(n_111), .B(n_453), .Y(n_466) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_111), .B(n_452), .Y(n_753) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B(n_458), .Y(n_115) );
HB1xp67_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx3_ASAP7_75t_L g757 ( .A(n_117), .Y(n_757) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_449), .B(n_455), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B1(n_126), .B2(n_127), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_126), .A2(n_461), .B1(n_464), .B2(n_467), .Y(n_460) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_127), .A2(n_461), .B1(n_755), .B2(n_756), .Y(n_754) );
AND2x2_ASAP7_75t_SL g127 ( .A(n_128), .B(n_404), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_339), .Y(n_128) );
NAND4xp25_ASAP7_75t_SL g129 ( .A(n_130), .B(n_284), .C(n_308), .D(n_331), .Y(n_129) );
AOI221xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_221), .B1(n_255), .B2(n_268), .C(n_271), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_191), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_133), .A2(n_169), .B1(n_222), .B2(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_133), .B(n_192), .Y(n_342) );
AND2x2_ASAP7_75t_L g361 ( .A(n_133), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_133), .B(n_345), .Y(n_431) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_169), .Y(n_133) );
AND2x2_ASAP7_75t_L g299 ( .A(n_134), .B(n_192), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_134), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g322 ( .A(n_134), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g327 ( .A(n_134), .B(n_170), .Y(n_327) );
INVx2_ASAP7_75t_L g359 ( .A(n_134), .Y(n_359) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_134), .Y(n_403) );
AND2x2_ASAP7_75t_L g420 ( .A(n_134), .B(n_297), .Y(n_420) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g338 ( .A(n_135), .B(n_297), .Y(n_338) );
AND2x4_ASAP7_75t_L g352 ( .A(n_135), .B(n_169), .Y(n_352) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_135), .Y(n_356) );
AND2x2_ASAP7_75t_L g376 ( .A(n_135), .B(n_291), .Y(n_376) );
AND2x2_ASAP7_75t_L g426 ( .A(n_135), .B(n_193), .Y(n_426) );
AND2x2_ASAP7_75t_L g436 ( .A(n_135), .B(n_170), .Y(n_436) );
OR2x6_ASAP7_75t_L g135 ( .A(n_136), .B(n_166), .Y(n_135) );
AOI21xp5_ASAP7_75t_SL g136 ( .A1(n_137), .A2(n_146), .B(n_159), .Y(n_136) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
NAND2x1p5_ASAP7_75t_L g260 ( .A(n_140), .B(n_144), .Y(n_260) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx1_ASAP7_75t_L g254 ( .A(n_142), .Y(n_254) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_143), .Y(n_153) );
INVx3_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_143), .Y(n_186) );
INVx1_ASAP7_75t_L g250 ( .A(n_143), .Y(n_250) );
BUFx3_ASAP7_75t_L g158 ( .A(n_144), .Y(n_158) );
INVx4_ASAP7_75t_SL g189 ( .A(n_144), .Y(n_189) );
INVx5_ASAP7_75t_L g178 ( .A(n_147), .Y(n_178) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_154), .B(n_156), .Y(n_150) );
INVx2_ASAP7_75t_L g155 ( .A(n_152), .Y(n_155) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g214 ( .A(n_153), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_155), .A2(n_199), .B(n_200), .C(n_201), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_155), .A2(n_201), .B(n_228), .C(n_229), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_155), .A2(n_500), .B(n_501), .C(n_502), .Y(n_499) );
O2A1O1Ixp5_ASAP7_75t_L g525 ( .A1(n_155), .A2(n_502), .B(n_526), .C(n_527), .Y(n_525) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_156), .A2(n_181), .B(n_477), .C(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_157), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_160), .B(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g168 ( .A(n_161), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_161), .A2(n_195), .B(n_196), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_161), .A2(n_225), .B(n_226), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_161), .A2(n_260), .B(n_474), .C(n_475), .Y(n_473) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_161), .A2(n_510), .B(n_517), .Y(n_509) );
AND2x2_ASAP7_75t_SL g161 ( .A(n_162), .B(n_163), .Y(n_161) );
AND2x2_ASAP7_75t_L g174 ( .A(n_162), .B(n_163), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_168), .A2(n_522), .B(n_528), .Y(n_521) );
AND2x2_ASAP7_75t_L g292 ( .A(n_169), .B(n_192), .Y(n_292) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_169), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_169), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g382 ( .A(n_169), .Y(n_382) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g270 ( .A(n_170), .B(n_207), .Y(n_270) );
AND2x2_ASAP7_75t_L g297 ( .A(n_170), .B(n_208), .Y(n_297) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_175), .B(n_190), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_172), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_172), .A2(n_209), .B(n_219), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_172), .B(n_220), .Y(n_219) );
AO21x2_ASAP7_75t_L g257 ( .A1(n_172), .A2(n_258), .B(n_265), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_172), .B(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_172), .A2(n_496), .B(n_503), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_172), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_173), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_173), .A2(n_246), .B(n_247), .Y(n_245) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g267 ( .A(n_174), .Y(n_267) );
O2A1O1Ixp33_ASAP7_75t_SL g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_189), .Y(n_176) );
INVx2_ASAP7_75t_L g197 ( .A(n_178), .Y(n_197) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_178), .A2(n_189), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g487 ( .A1(n_178), .A2(n_189), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g511 ( .A1(n_178), .A2(n_189), .B(n_512), .C(n_513), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_178), .A2(n_189), .B(n_534), .C(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_178), .A2(n_189), .B(n_551), .C(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_SL g563 ( .A1(n_178), .A2(n_189), .B(n_564), .C(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_181), .B(n_240), .Y(n_239) );
OAI22xp33_ASAP7_75t_L g490 ( .A1(n_181), .A2(n_214), .B1(n_491), .B2(n_492), .Y(n_490) );
INVx5_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_182), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_185), .B(n_554), .Y(n_553) );
INVx4_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g514 ( .A(n_186), .Y(n_514) );
INVx2_ASAP7_75t_L g502 ( .A(n_187), .Y(n_502) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_188), .Y(n_201) );
INVx1_ASAP7_75t_L g538 ( .A(n_188), .Y(n_538) );
INVx1_ASAP7_75t_L g202 ( .A(n_189), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_191), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g191 ( .A(n_192), .B(n_205), .Y(n_191) );
OR2x2_ASAP7_75t_L g323 ( .A(n_192), .B(n_206), .Y(n_323) );
AND2x2_ASAP7_75t_L g360 ( .A(n_192), .B(n_270), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_192), .B(n_291), .Y(n_371) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_192), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_192), .B(n_327), .Y(n_444) );
INVx5_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
BUFx2_ASAP7_75t_L g269 ( .A(n_193), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_193), .B(n_206), .Y(n_278) );
AND2x2_ASAP7_75t_L g394 ( .A(n_193), .B(n_289), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_193), .B(n_327), .Y(n_416) );
OR2x6_ASAP7_75t_L g193 ( .A(n_194), .B(n_203), .Y(n_193) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_206), .Y(n_362) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_207), .Y(n_314) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx2_ASAP7_75t_L g291 ( .A(n_208), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_218), .Y(n_209) );
O2A1O1Ixp33_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_215), .C(n_216), .Y(n_211) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_214), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_214), .B(n_567), .Y(n_566) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx3_ASAP7_75t_L g555 ( .A(n_217), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_231), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_222), .B(n_304), .Y(n_423) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_223), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g275 ( .A(n_223), .B(n_276), .Y(n_275) );
INVx5_ASAP7_75t_SL g283 ( .A(n_223), .Y(n_283) );
OR2x2_ASAP7_75t_L g306 ( .A(n_223), .B(n_276), .Y(n_306) );
OR2x2_ASAP7_75t_L g316 ( .A(n_223), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g379 ( .A(n_223), .B(n_233), .Y(n_379) );
AND2x2_ASAP7_75t_SL g417 ( .A(n_223), .B(n_232), .Y(n_417) );
NOR4xp25_ASAP7_75t_L g438 ( .A(n_223), .B(n_359), .C(n_439), .D(n_440), .Y(n_438) );
AND2x2_ASAP7_75t_L g448 ( .A(n_223), .B(n_280), .Y(n_448) );
OR2x6_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g273 ( .A(n_232), .B(n_269), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_232), .B(n_275), .Y(n_442) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_242), .Y(n_232) );
OR2x2_ASAP7_75t_L g282 ( .A(n_233), .B(n_283), .Y(n_282) );
INVx3_ASAP7_75t_L g289 ( .A(n_233), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_233), .B(n_257), .Y(n_301) );
INVxp67_ASAP7_75t_L g304 ( .A(n_233), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_233), .B(n_276), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_233), .B(n_243), .Y(n_370) );
AND2x2_ASAP7_75t_L g385 ( .A(n_233), .B(n_280), .Y(n_385) );
OR2x2_ASAP7_75t_L g414 ( .A(n_233), .B(n_243), .Y(n_414) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_234), .A2(n_532), .B(n_539), .Y(n_531) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_234), .A2(n_549), .B(n_556), .Y(n_548) );
OA21x2_ASAP7_75t_L g561 ( .A1(n_234), .A2(n_562), .B(n_568), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_242), .B(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_242), .B(n_283), .Y(n_422) );
OR2x2_ASAP7_75t_L g443 ( .A(n_242), .B(n_320), .Y(n_443) );
INVx1_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g256 ( .A(n_243), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g280 ( .A(n_243), .B(n_276), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_243), .B(n_257), .Y(n_295) );
AND2x2_ASAP7_75t_L g365 ( .A(n_243), .B(n_289), .Y(n_365) );
AND2x2_ASAP7_75t_L g399 ( .A(n_243), .B(n_283), .Y(n_399) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_244), .B(n_283), .Y(n_302) );
AND2x2_ASAP7_75t_L g330 ( .A(n_244), .B(n_257), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_251), .B(n_252), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_252), .A2(n_263), .B(n_264), .Y(n_262) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_255), .B(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_256), .A2(n_345), .B1(n_381), .B2(n_398), .C(n_400), .Y(n_397) );
INVx5_ASAP7_75t_SL g276 ( .A(n_257), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_261), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_260), .A2(n_497), .B(n_498), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_260), .A2(n_523), .B(n_524), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_L g485 ( .A(n_267), .Y(n_485) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OAI33xp33_ASAP7_75t_L g296 ( .A1(n_269), .A2(n_297), .A3(n_298), .B1(n_300), .B2(n_303), .B3(n_307), .Y(n_296) );
OR2x2_ASAP7_75t_L g312 ( .A(n_269), .B(n_313), .Y(n_312) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_269), .A2(n_338), .A3(n_345), .B1(n_422), .B2(n_423), .C1(n_424), .C2(n_427), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_269), .B(n_297), .Y(n_439) );
A2O1A1Ixp33_ASAP7_75t_SL g445 ( .A1(n_269), .A2(n_297), .B(n_446), .C(n_448), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_270), .A2(n_285), .B1(n_290), .B2(n_293), .C(n_296), .Y(n_284) );
INVx1_ASAP7_75t_L g377 ( .A(n_270), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_270), .B(n_426), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B1(n_277), .B2(n_279), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g354 ( .A(n_275), .B(n_289), .Y(n_354) );
AND2x2_ASAP7_75t_L g412 ( .A(n_275), .B(n_413), .Y(n_412) );
OR2x2_ASAP7_75t_L g320 ( .A(n_276), .B(n_283), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_276), .B(n_289), .Y(n_348) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_278), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_278), .B(n_356), .Y(n_410) );
OAI321xp33_ASAP7_75t_L g429 ( .A1(n_278), .A2(n_351), .A3(n_430), .B1(n_431), .B2(n_432), .C(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g396 ( .A(n_279), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_280), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g335 ( .A(n_280), .B(n_283), .Y(n_335) );
AOI321xp33_ASAP7_75t_L g393 ( .A1(n_280), .A2(n_297), .A3(n_394), .B1(n_395), .B2(n_396), .C(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g310 ( .A(n_282), .B(n_295), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_283), .B(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_283), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_283), .B(n_369), .Y(n_406) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g329 ( .A(n_287), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g294 ( .A(n_288), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g402 ( .A(n_289), .Y(n_402) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_292), .B(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g325 ( .A(n_297), .Y(n_325) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_299), .B(n_334), .Y(n_383) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
OR2x2_ASAP7_75t_L g347 ( .A(n_302), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g392 ( .A(n_302), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_303), .A2(n_350), .B1(n_353), .B2(n_355), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g447 ( .A(n_306), .B(n_370), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B1(n_315), .B2(n_321), .C(n_324), .Y(n_308) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_L g345 ( .A(n_314), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
INVx1_ASAP7_75t_SL g391 ( .A(n_317), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_319), .B(n_369), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_319), .A2(n_387), .B(n_389), .Y(n_386) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g432 ( .A(n_320), .B(n_414), .Y(n_432) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_SL g334 ( .A(n_323), .Y(n_334) );
AOI21xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g378 ( .A(n_330), .B(n_379), .Y(n_378) );
INVxp67_ASAP7_75t_L g440 ( .A(n_330), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_335), .B(n_336), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_334), .B(n_352), .Y(n_388) );
INVxp67_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g409 ( .A(n_338), .Y(n_409) );
NAND5xp2_ASAP7_75t_L g339 ( .A(n_340), .B(n_357), .C(n_366), .D(n_386), .E(n_393), .Y(n_339) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B(n_346), .C(n_349), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
CKINVDCx16_ASAP7_75t_R g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_353), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g395 ( .A(n_355), .Y(n_395) );
OAI21xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_361), .B(n_363), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_358), .A2(n_412), .B1(n_415), .B2(n_417), .C(n_418), .Y(n_411) );
AND2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AOI321xp33_ASAP7_75t_L g366 ( .A1(n_359), .A2(n_367), .A3(n_371), .B1(n_372), .B2(n_378), .C(n_380), .Y(n_366) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g437 ( .A(n_371), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g372 ( .A(n_373), .B(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g389 ( .A(n_374), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NOR2xp67_ASAP7_75t_SL g401 ( .A(n_375), .B(n_382), .Y(n_401) );
AOI321xp33_ASAP7_75t_SL g433 ( .A1(n_378), .A2(n_434), .A3(n_435), .B1(n_436), .B2(n_437), .C(n_438), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .C(n_384), .Y(n_380) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_391), .B(n_399), .Y(n_428) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .C(n_403), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_429), .C(n_441), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g405 ( .A1(n_406), .A2(n_407), .B(n_411), .C(n_421), .Y(n_405) );
INVxp67_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_409), .B(n_410), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g441 ( .A1(n_410), .A2(n_442), .B1(n_443), .B2(n_444), .C(n_445), .Y(n_441) );
INVx1_ASAP7_75t_L g430 ( .A(n_412), .Y(n_430) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g434 ( .A(n_432), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
CKINVDCx14_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g457 ( .A(n_451), .Y(n_457) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_455), .A2(n_459), .B(n_757), .Y(n_458) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g756 ( .A(n_465), .Y(n_756) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g755 ( .A(n_467), .Y(n_755) );
OR4x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_637), .C(n_684), .D(n_724), .Y(n_467) );
NAND3xp33_ASAP7_75t_SL g468 ( .A(n_469), .B(n_583), .C(n_612), .Y(n_468) );
AOI211xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_505), .B(n_540), .C(n_576), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_470), .A2(n_596), .B(n_613), .C(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_472), .B(n_481), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_472), .B(n_575), .Y(n_574) );
INVx3_ASAP7_75t_SL g579 ( .A(n_472), .Y(n_579) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_472), .Y(n_591) );
AND2x4_ASAP7_75t_L g595 ( .A(n_472), .B(n_547), .Y(n_595) );
AND2x2_ASAP7_75t_L g606 ( .A(n_472), .B(n_495), .Y(n_606) );
OR2x2_ASAP7_75t_L g630 ( .A(n_472), .B(n_543), .Y(n_630) );
AND2x2_ASAP7_75t_L g643 ( .A(n_472), .B(n_548), .Y(n_643) );
AND2x2_ASAP7_75t_L g683 ( .A(n_472), .B(n_669), .Y(n_683) );
AND2x2_ASAP7_75t_L g690 ( .A(n_472), .B(n_653), .Y(n_690) );
AND2x2_ASAP7_75t_L g720 ( .A(n_472), .B(n_482), .Y(n_720) );
OR2x6_ASAP7_75t_L g472 ( .A(n_473), .B(n_479), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_481), .B(n_647), .Y(n_659) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_494), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_482), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g597 ( .A(n_482), .B(n_494), .Y(n_597) );
BUFx3_ASAP7_75t_L g605 ( .A(n_482), .Y(n_605) );
OR2x2_ASAP7_75t_L g626 ( .A(n_482), .B(n_508), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_482), .B(n_647), .Y(n_737) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B(n_493), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AO21x2_ASAP7_75t_L g543 ( .A1(n_484), .A2(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g544 ( .A(n_486), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_493), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_494), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g590 ( .A(n_494), .Y(n_590) );
AND2x2_ASAP7_75t_L g653 ( .A(n_494), .B(n_548), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_494), .A2(n_656), .B1(n_658), .B2(n_660), .C(n_661), .Y(n_655) );
AND2x2_ASAP7_75t_L g669 ( .A(n_494), .B(n_543), .Y(n_669) );
AND2x2_ASAP7_75t_L g695 ( .A(n_494), .B(n_579), .Y(n_695) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g575 ( .A(n_495), .B(n_548), .Y(n_575) );
BUFx2_ASAP7_75t_L g709 ( .A(n_495), .Y(n_709) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
OAI32xp33_ASAP7_75t_L g675 ( .A1(n_506), .A2(n_636), .A3(n_650), .B1(n_676), .B2(n_677), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
AND2x2_ASAP7_75t_L g616 ( .A(n_507), .B(n_560), .Y(n_616) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g598 ( .A(n_508), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_508), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g670 ( .A(n_508), .B(n_560), .Y(n_670) );
AND2x2_ASAP7_75t_L g681 ( .A(n_508), .B(n_573), .Y(n_681) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g582 ( .A(n_509), .B(n_561), .Y(n_582) );
AND2x2_ASAP7_75t_L g586 ( .A(n_509), .B(n_561), .Y(n_586) );
AND2x2_ASAP7_75t_L g621 ( .A(n_509), .B(n_572), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_509), .B(n_530), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g633 ( .A1(n_509), .A2(n_579), .B(n_590), .C(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g687 ( .A(n_509), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_509), .B(n_520), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_518), .B(n_570), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_518), .B(n_586), .Y(n_676) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
OR2x2_ASAP7_75t_L g581 ( .A(n_519), .B(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_530), .Y(n_519) );
AND2x2_ASAP7_75t_L g573 ( .A(n_520), .B(n_531), .Y(n_573) );
OR2x2_ASAP7_75t_L g588 ( .A(n_520), .B(n_531), .Y(n_588) );
AND2x2_ASAP7_75t_L g611 ( .A(n_520), .B(n_572), .Y(n_611) );
INVx1_ASAP7_75t_L g615 ( .A(n_520), .Y(n_615) );
AND2x2_ASAP7_75t_L g634 ( .A(n_520), .B(n_571), .Y(n_634) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_520), .A2(n_599), .B1(n_645), .B2(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_520), .B(n_687), .Y(n_711) );
AND2x2_ASAP7_75t_L g726 ( .A(n_520), .B(n_586), .Y(n_726) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx3_ASAP7_75t_L g558 ( .A(n_521), .Y(n_558) );
AND2x2_ASAP7_75t_L g600 ( .A(n_521), .B(n_531), .Y(n_600) );
AND2x2_ASAP7_75t_L g602 ( .A(n_521), .B(n_560), .Y(n_602) );
AND3x2_ASAP7_75t_L g664 ( .A(n_521), .B(n_628), .C(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g699 ( .A(n_530), .B(n_571), .Y(n_699) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g560 ( .A(n_531), .B(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_531), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_531), .B(n_570), .Y(n_632) );
NAND3xp33_ASAP7_75t_L g739 ( .A(n_531), .B(n_611), .C(n_687), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_557), .B1(n_569), .B2(n_574), .Y(n_540) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_546), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_543), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g651 ( .A(n_543), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g667 ( .A1(n_546), .A2(n_668), .A3(n_669), .B(n_670), .Y(n_667) );
AND2x2_ASAP7_75t_L g692 ( .A(n_546), .B(n_579), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_546), .B(n_605), .Y(n_738) );
AND2x2_ASAP7_75t_L g647 ( .A(n_547), .B(n_579), .Y(n_647) );
AND2x2_ASAP7_75t_L g708 ( .A(n_547), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g578 ( .A(n_548), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g636 ( .A(n_548), .Y(n_636) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
CKINVDCx16_ASAP7_75t_R g657 ( .A(n_558), .Y(n_657) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_559), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
AOI221x1_ASAP7_75t_SL g624 ( .A1(n_560), .A2(n_625), .B1(n_627), .B2(n_629), .C(n_631), .Y(n_624) );
INVx2_ASAP7_75t_L g572 ( .A(n_561), .Y(n_572) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_561), .Y(n_666) );
INVx1_ASAP7_75t_L g654 ( .A(n_569), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_570), .B(n_587), .Y(n_679) );
INVx1_ASAP7_75t_SL g742 ( .A(n_570), .Y(n_742) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g660 ( .A(n_573), .B(n_586), .Y(n_660) );
INVx1_ASAP7_75t_L g728 ( .A(n_574), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_574), .B(n_657), .Y(n_741) );
INVx2_ASAP7_75t_SL g580 ( .A(n_575), .Y(n_580) );
AND2x2_ASAP7_75t_L g623 ( .A(n_575), .B(n_579), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_575), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_575), .B(n_650), .Y(n_677) );
AOI21xp33_ASAP7_75t_SL g576 ( .A1(n_577), .A2(n_580), .B(n_581), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_578), .B(n_650), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_578), .B(n_605), .Y(n_746) );
OR2x2_ASAP7_75t_L g618 ( .A(n_579), .B(n_597), .Y(n_618) );
AND2x2_ASAP7_75t_L g717 ( .A(n_579), .B(n_708), .Y(n_717) );
OAI22xp5_ASAP7_75t_SL g592 ( .A1(n_580), .A2(n_593), .B1(n_598), .B2(n_601), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_580), .B(n_626), .Y(n_625) );
OR2x2_ASAP7_75t_L g640 ( .A(n_582), .B(n_588), .Y(n_640) );
INVx1_ASAP7_75t_L g704 ( .A(n_582), .Y(n_704) );
AOI311xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_589), .A3(n_591), .B(n_592), .C(n_603), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g730 ( .A1(n_587), .A2(n_719), .B1(n_731), .B2(n_734), .C(n_736), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_587), .B(n_742), .Y(n_744) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g641 ( .A(n_589), .Y(n_641) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_590), .A2(n_632), .B(n_633), .C(n_635), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
O2A1O1Ixp33_ASAP7_75t_SL g700 ( .A1(n_594), .A2(n_596), .B(n_701), .C(n_702), .Y(n_700) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_595), .B(n_669), .Y(n_735) );
INVx1_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
OAI221xp5_ASAP7_75t_L g617 ( .A1(n_598), .A2(n_618), .B1(n_619), .B2(n_622), .C(n_624), .Y(n_617) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g620 ( .A(n_600), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g703 ( .A(n_600), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
A2O1A1Ixp33_ASAP7_75t_L g661 ( .A1(n_604), .A2(n_662), .B(n_663), .C(n_667), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_605), .B(n_606), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_605), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_605), .B(n_708), .Y(n_707) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g627 ( .A(n_611), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_615), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g729 ( .A(n_618), .Y(n_729) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_621), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g656 ( .A(n_621), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_SL g733 ( .A(n_621), .Y(n_733) );
INVx1_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g674 ( .A(n_623), .B(n_650), .Y(n_674) );
INVx1_ASAP7_75t_SL g668 ( .A(n_630), .Y(n_668) );
INVx1_ASAP7_75t_L g645 ( .A(n_636), .Y(n_645) );
NAND3xp33_ASAP7_75t_SL g637 ( .A(n_638), .B(n_655), .C(n_671), .Y(n_637) );
AOI322xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .A3(n_642), .B1(n_644), .B2(n_648), .C1(n_652), .C2(n_654), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_639), .A2(n_692), .B(n_693), .C(n_700), .Y(n_691) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_642), .A2(n_663), .B1(n_694), .B2(n_696), .Y(n_693) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g652 ( .A(n_650), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g689 ( .A(n_650), .B(n_690), .Y(n_689) );
AOI32xp33_ASAP7_75t_L g740 ( .A1(n_650), .A2(n_741), .A3(n_742), .B1(n_743), .B2(n_745), .Y(n_740) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g662 ( .A(n_653), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_653), .A2(n_706), .B1(n_710), .B2(n_712), .C(n_715), .Y(n_705) );
AND2x2_ASAP7_75t_L g719 ( .A(n_653), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g722 ( .A(n_657), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g732 ( .A(n_657), .B(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g723 ( .A(n_666), .B(n_687), .Y(n_723) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B(n_675), .C(n_678), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B(n_682), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g684 ( .A1(n_685), .A2(n_688), .B(n_691), .C(n_705), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_699), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g714 ( .A(n_711), .Y(n_714) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_718), .B(n_721), .Y(n_715) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OAI211xp5_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_727), .B(n_730), .C(n_740), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_726), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI21xp33_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B(n_739), .Y(n_736) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
endmodule