module real_aes_5224_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_666;
wire n_320;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_948;
wire n_677;
wire n_958;
wire n_1046;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_559;
wire n_466;
wire n_1049;
wire n_636;
wire n_872;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_931;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_755;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_488;
wire n_1041;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_1056;
wire n_358;
wire n_385;
wire n_397;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_1040;
wire n_652;
wire n_703;
wire n_393;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_0), .A2(n_267), .B1(n_558), .B2(n_559), .Y(n_591) );
AO22x2_ASAP7_75t_L g572 ( .A1(n_1), .A2(n_573), .B1(n_593), .B2(n_594), .Y(n_572) );
INVxp67_ASAP7_75t_SL g593 ( .A(n_1), .Y(n_593) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_2), .Y(n_779) );
AND2x4_ASAP7_75t_L g787 ( .A(n_2), .B(n_788), .Y(n_787) );
AND2x4_ASAP7_75t_L g796 ( .A(n_2), .B(n_287), .Y(n_796) );
AOI22xp33_ASAP7_75t_SL g792 ( .A1(n_3), .A2(n_63), .B1(n_793), .B2(n_797), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_4), .A2(n_35), .B1(n_332), .B2(n_527), .Y(n_726) );
INVx1_ASAP7_75t_L g428 ( .A(n_5), .Y(n_428) );
INVx1_ASAP7_75t_L g688 ( .A(n_6), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g1015 ( .A1(n_7), .A2(n_180), .B1(n_307), .B2(n_352), .Y(n_1015) );
AOI22xp33_ASAP7_75t_L g1017 ( .A1(n_8), .A2(n_165), .B1(n_332), .B2(n_534), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_9), .A2(n_120), .B1(n_413), .B2(n_489), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_10), .A2(n_145), .B1(n_532), .B2(n_729), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_11), .A2(n_231), .B1(n_307), .B2(n_332), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_12), .A2(n_124), .B1(n_811), .B2(n_812), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_13), .A2(n_259), .B1(n_342), .B2(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_14), .A2(n_108), .B1(n_558), .B2(n_559), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_15), .A2(n_207), .B1(n_332), .B2(n_484), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_16), .A2(n_21), .B1(n_555), .B2(n_556), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_17), .A2(n_59), .B1(n_347), .B2(n_529), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_18), .A2(n_27), .B1(n_451), .B2(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g1050 ( .A(n_19), .B(n_502), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_20), .A2(n_90), .B1(n_647), .B2(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_22), .A2(n_135), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_23), .A2(n_36), .B1(n_413), .B2(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g1029 ( .A(n_24), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_25), .A2(n_31), .B1(n_431), .B2(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_26), .A2(n_176), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_28), .A2(n_242), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_29), .A2(n_143), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_30), .A2(n_150), .B1(n_442), .B2(n_559), .Y(n_612) );
INVx1_ASAP7_75t_L g711 ( .A(n_32), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_33), .A2(n_136), .B1(n_384), .B2(n_387), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_34), .A2(n_137), .B1(n_370), .B2(n_516), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_37), .A2(n_43), .B1(n_423), .B2(n_536), .C(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g519 ( .A(n_38), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_39), .A2(n_171), .B1(n_364), .B2(n_451), .Y(n_699) );
AOI21x1_ASAP7_75t_L g707 ( .A1(n_40), .A2(n_708), .B(n_710), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_41), .A2(n_192), .B1(n_438), .B2(n_439), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_42), .A2(n_497), .B(n_498), .Y(n_496) );
XOR2x2_ASAP7_75t_L g740 ( .A(n_44), .B(n_741), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_45), .A2(n_291), .B1(n_529), .B2(n_731), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_46), .A2(n_244), .B1(n_713), .B2(n_737), .Y(n_736) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_47), .A2(n_118), .B1(n_786), .B2(n_790), .Y(n_785) );
XNOR2x1_ASAP7_75t_L g511 ( .A(n_48), .B(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_49), .A2(n_200), .B1(n_646), .B2(n_648), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g422 ( .A1(n_50), .A2(n_423), .B(n_426), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_51), .A2(n_89), .B1(n_342), .B2(n_654), .Y(n_746) );
INVx1_ASAP7_75t_L g329 ( .A(n_52), .Y(n_329) );
INVxp67_ASAP7_75t_L g382 ( .A(n_52), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_52), .B(n_226), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_53), .A2(n_144), .B1(n_497), .B2(n_555), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_54), .A2(n_182), .B1(n_489), .B2(n_529), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_55), .A2(n_96), .B1(n_396), .B2(n_505), .Y(n_683) );
INVx1_ASAP7_75t_L g1049 ( .A(n_56), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_57), .A2(n_116), .B1(n_456), .B2(n_457), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_58), .A2(n_146), .B1(n_493), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_60), .A2(n_175), .B1(n_471), .B2(n_536), .Y(n_735) );
XNOR2x1_ASAP7_75t_L g620 ( .A(n_61), .B(n_621), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_61), .A2(n_277), .B1(n_801), .B2(n_822), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_62), .A2(n_203), .B1(n_793), .B2(n_797), .Y(n_828) );
XNOR2x1_ASAP7_75t_L g480 ( .A(n_63), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_64), .B(n_313), .Y(n_325) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_65), .A2(n_132), .B1(n_396), .B2(n_421), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_66), .A2(n_100), .B1(n_351), .B2(n_354), .Y(n_350) );
AOI21xp33_ASAP7_75t_SL g575 ( .A1(n_67), .A2(n_431), .B(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_68), .A2(n_274), .B1(n_532), .B2(n_729), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_69), .A2(n_212), .B1(n_352), .B2(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g566 ( .A(n_70), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_71), .A2(n_278), .B1(n_432), .B2(n_435), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_72), .A2(n_193), .B1(n_392), .B2(n_396), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_73), .A2(n_248), .B1(n_352), .B2(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_74), .A2(n_245), .B1(n_432), .B2(n_434), .Y(n_603) );
BUFx2_ASAP7_75t_L g581 ( .A(n_75), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_76), .A2(n_114), .B1(n_555), .B2(n_556), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_77), .A2(n_131), .B1(n_811), .B2(n_812), .Y(n_872) );
INVx1_ASAP7_75t_L g687 ( .A(n_78), .Y(n_687) );
INVx2_ASAP7_75t_L g777 ( .A(n_79), .Y(n_777) );
INVx1_ASAP7_75t_L g749 ( .A(n_80), .Y(n_749) );
INVx1_ASAP7_75t_SL g789 ( .A(n_81), .Y(n_789) );
AND2x4_ASAP7_75t_L g791 ( .A(n_81), .B(n_777), .Y(n_791) );
INVx1_ASAP7_75t_L g795 ( .A(n_81), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_82), .A2(n_263), .B1(n_396), .B2(n_431), .Y(n_548) );
INVx1_ASAP7_75t_L g750 ( .A(n_83), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_84), .A2(n_264), .B1(n_757), .B2(n_759), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_85), .A2(n_190), .B1(n_370), .B2(n_373), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_86), .B(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g1054 ( .A1(n_87), .A2(n_189), .B1(n_491), .B2(n_647), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_88), .A2(n_255), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_91), .A2(n_257), .B1(n_354), .B2(n_456), .Y(n_700) );
AOI22xp33_ASAP7_75t_SL g460 ( .A1(n_92), .A2(n_270), .B1(n_307), .B2(n_332), .Y(n_460) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_93), .Y(n_313) );
AOI22xp5_ASAP7_75t_L g837 ( .A1(n_94), .A2(n_178), .B1(n_793), .B2(n_797), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_95), .A2(n_228), .B1(n_438), .B2(n_439), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_97), .A2(n_206), .B1(n_358), .B2(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g541 ( .A(n_98), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_99), .A2(n_215), .B1(n_352), .B2(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g561 ( .A(n_101), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_102), .A2(n_292), .B1(n_556), .B2(n_558), .Y(n_609) );
INVx1_ASAP7_75t_L g819 ( .A(n_103), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_104), .A2(n_105), .B1(n_435), .B2(n_441), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g827 ( .A1(n_106), .A2(n_289), .B1(n_786), .B2(n_790), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_107), .A2(n_239), .B1(n_470), .B2(n_471), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_109), .A2(n_296), .B1(n_370), .B2(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g314 ( .A(n_110), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_110), .B(n_225), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_111), .A2(n_117), .B1(n_786), .B2(n_790), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_112), .A2(n_169), .B1(n_332), .B2(n_484), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_113), .A2(n_196), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_115), .A2(n_191), .B1(n_504), .B2(n_516), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_119), .A2(n_237), .B1(n_434), .B2(n_497), .Y(n_663) );
XNOR2x1_ASAP7_75t_L g598 ( .A(n_121), .B(n_599), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_122), .A2(n_205), .B1(n_477), .B2(n_478), .Y(n_476) );
INVx1_ASAP7_75t_L g765 ( .A(n_123), .Y(n_765) );
INVx1_ASAP7_75t_L g447 ( .A(n_125), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_125), .A2(n_229), .B1(n_793), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g753 ( .A(n_126), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_127), .A2(n_1041), .B1(n_1042), .B2(n_1056), .Y(n_1040) );
CKINVDCx5p33_ASAP7_75t_R g1041 ( .A(n_127), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_128), .A2(n_174), .B1(n_342), .B2(n_459), .Y(n_697) );
INVxp33_ASAP7_75t_SL g825 ( .A(n_129), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_130), .A2(n_290), .B1(n_441), .B2(n_442), .Y(n_589) );
XNOR2x1_ASAP7_75t_L g409 ( .A(n_133), .B(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_134), .A2(n_153), .B1(n_624), .B2(n_625), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_138), .A2(n_252), .B1(n_358), .B2(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g637 ( .A(n_139), .Y(n_637) );
INVx1_ASAP7_75t_L g577 ( .A(n_140), .Y(n_577) );
INVx1_ASAP7_75t_L g419 ( .A(n_141), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_142), .A2(n_183), .B1(n_808), .B2(n_809), .Y(n_873) );
CKINVDCx16_ASAP7_75t_R g1032 ( .A(n_142), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1037 ( .A1(n_142), .A2(n_1038), .B1(n_1040), .B2(n_1057), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_147), .A2(n_271), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI21xp33_ASAP7_75t_L g604 ( .A1(n_148), .A2(n_605), .B(n_606), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_149), .A2(n_260), .B1(n_438), .B2(n_439), .Y(n_551) );
INVx1_ASAP7_75t_L g607 ( .A(n_151), .Y(n_607) );
INVx1_ASAP7_75t_L g521 ( .A(n_152), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_154), .A2(n_285), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_155), .A2(n_184), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g587 ( .A1(n_156), .A2(n_256), .B1(n_421), .B2(n_435), .Y(n_587) );
AOI21xp33_ASAP7_75t_L g1047 ( .A1(n_157), .A2(n_628), .B(n_1048), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_158), .A2(n_167), .B1(n_485), .B2(n_760), .Y(n_1055) );
AOI22xp5_ASAP7_75t_L g1053 ( .A1(n_159), .A2(n_230), .B1(n_493), .B2(n_532), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1025 ( .A1(n_160), .A2(n_240), .B1(n_516), .B2(n_1026), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_161), .A2(n_163), .B1(n_491), .B2(n_529), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g743 ( .A1(n_162), .A2(n_258), .B1(n_459), .B2(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g549 ( .A1(n_164), .A2(n_199), .B1(n_373), .B2(n_516), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_166), .A2(n_214), .B1(n_396), .B2(n_421), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_168), .B(n_389), .Y(n_601) );
INVx1_ASAP7_75t_L g499 ( .A(n_170), .Y(n_499) );
INVx1_ASAP7_75t_L g823 ( .A(n_172), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_173), .A2(n_272), .B1(n_536), .B2(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g752 ( .A(n_177), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_179), .A2(n_210), .B1(n_652), .B2(n_653), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_181), .A2(n_370), .B(n_1028), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_185), .B(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_186), .A2(n_276), .B1(n_493), .B2(n_494), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_187), .A2(n_236), .B1(n_352), .B2(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g658 ( .A(n_188), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_194), .A2(n_213), .B1(n_627), .B2(n_629), .Y(n_626) );
OA22x2_ASAP7_75t_L g319 ( .A1(n_195), .A2(n_226), .B1(n_313), .B2(n_317), .Y(n_319) );
INVx1_ASAP7_75t_L g338 ( .A(n_195), .Y(n_338) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_197), .A2(n_632), .B(n_635), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_198), .A2(n_294), .B1(n_332), .B2(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_201), .A2(n_250), .B1(n_493), .B2(n_532), .Y(n_680) );
XOR2x2_ASAP7_75t_L g303 ( .A(n_202), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g640 ( .A(n_204), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_208), .A2(n_282), .B1(n_808), .B2(n_809), .Y(n_807) );
INVx1_ASAP7_75t_SL g738 ( .A(n_209), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_211), .A2(n_251), .B1(n_524), .B2(n_628), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_216), .A2(n_284), .B1(n_536), .B2(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g552 ( .A1(n_217), .A2(n_224), .B1(n_441), .B2(n_442), .Y(n_552) );
XOR2x2_ASAP7_75t_L g693 ( .A(n_218), .B(n_694), .Y(n_693) );
NAND2xp33_ASAP7_75t_L g1020 ( .A(n_219), .B(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g567 ( .A(n_220), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_221), .B(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g585 ( .A(n_222), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_223), .A2(n_254), .B1(n_438), .B2(n_439), .Y(n_592) );
INVx1_ASAP7_75t_L g331 ( .A(n_225), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_225), .B(n_336), .Y(n_407) );
OAI21xp33_ASAP7_75t_L g339 ( .A1(n_226), .A2(n_241), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g866 ( .A(n_227), .Y(n_866) );
INVx1_ASAP7_75t_L g865 ( .A(n_232), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g836 ( .A1(n_233), .A2(n_253), .B1(n_786), .B2(n_790), .Y(n_836) );
INVx1_ASAP7_75t_L g517 ( .A(n_234), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_235), .A2(n_275), .B1(n_441), .B2(n_442), .Y(n_669) );
INVx1_ASAP7_75t_L g466 ( .A(n_238), .Y(n_466) );
INVx1_ASAP7_75t_L g316 ( .A(n_241), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_241), .B(n_279), .Y(n_405) );
AOI21xp33_ASAP7_75t_L g464 ( .A1(n_243), .A2(n_370), .B(n_465), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g769 ( .A1(n_246), .A2(n_261), .B1(n_524), .B2(n_543), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_247), .A2(n_281), .B1(n_536), .B2(n_537), .C(n_540), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_249), .A2(n_425), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g667 ( .A(n_262), .Y(n_667) );
AOI21xp33_ASAP7_75t_L g665 ( .A1(n_265), .A2(n_605), .B(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_266), .A2(n_269), .B1(n_342), .B2(n_347), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_268), .A2(n_389), .B(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_273), .B(n_634), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_279), .B(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_280), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_283), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g714 ( .A(n_286), .Y(n_714) );
INVx1_ASAP7_75t_L g788 ( .A(n_287), .Y(n_788) );
HB1xp67_ASAP7_75t_L g1059 ( .A(n_287), .Y(n_1059) );
INVxp33_ASAP7_75t_L g817 ( .A(n_288), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_293), .A2(n_295), .B1(n_451), .B2(n_532), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_616), .B(n_771), .C(n_780), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g771 ( .A1(n_298), .A2(n_616), .B(n_772), .Y(n_771) );
XOR2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_507), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_443), .B2(n_506), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
XNOR2x1_ASAP7_75t_L g302 ( .A(n_303), .B(n_408), .Y(n_302) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_305), .B(n_368), .Y(n_304) );
NAND4xp25_ASAP7_75t_SL g305 ( .A(n_306), .B(n_341), .C(n_350), .D(n_357), .Y(n_305) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_308), .Y(n_484) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_308), .Y(n_527) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_308), .Y(n_760) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_320), .Y(n_308) );
AND2x4_ASAP7_75t_L g353 ( .A(n_309), .B(n_345), .Y(n_353) );
AND2x4_ASAP7_75t_L g361 ( .A(n_309), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g365 ( .A(n_309), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g438 ( .A(n_309), .B(n_362), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_309), .B(n_366), .Y(n_439) );
AND2x4_ASAP7_75t_L g441 ( .A(n_309), .B(n_349), .Y(n_441) );
AND2x4_ASAP7_75t_L g558 ( .A(n_309), .B(n_345), .Y(n_558) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_318), .Y(n_309) );
AND2x2_ASAP7_75t_L g372 ( .A(n_310), .B(n_319), .Y(n_372) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g344 ( .A(n_311), .B(n_319), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_315), .Y(n_311) );
NAND2xp33_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx2_ASAP7_75t_L g317 ( .A(n_313), .Y(n_317) );
INVx3_ASAP7_75t_L g324 ( .A(n_313), .Y(n_324) );
NAND2xp33_ASAP7_75t_L g330 ( .A(n_313), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g340 ( .A(n_313), .Y(n_340) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_313), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_314), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_316), .A2(n_340), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g380 ( .A(n_319), .B(n_381), .Y(n_380) );
AND2x4_ASAP7_75t_L g333 ( .A(n_320), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g442 ( .A(n_320), .B(n_334), .Y(n_442) );
AND2x4_ASAP7_75t_L g556 ( .A(n_320), .B(n_344), .Y(n_556) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g349 ( .A(n_321), .Y(n_349) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
AND2x4_ASAP7_75t_L g345 ( .A(n_322), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g362 ( .A(n_322), .B(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g367 ( .A(n_322), .Y(n_367) );
AND2x2_ASAP7_75t_L g376 ( .A(n_322), .B(n_377), .Y(n_376) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_324), .B(n_329), .Y(n_328) );
INVxp67_ASAP7_75t_L g336 ( .A(n_324), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g406 ( .A(n_325), .B(n_335), .C(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g346 ( .A(n_326), .Y(n_346) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g363 ( .A(n_327), .Y(n_363) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
BUFx3_ASAP7_75t_L g644 ( .A(n_332), .Y(n_644) );
BUFx12f_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx6_ASAP7_75t_L g486 ( .A(n_333), .Y(n_486) );
AND2x4_ASAP7_75t_L g356 ( .A(n_334), .B(n_345), .Y(n_356) );
AND2x4_ASAP7_75t_L g397 ( .A(n_334), .B(n_366), .Y(n_397) );
AND2x4_ASAP7_75t_L g435 ( .A(n_334), .B(n_366), .Y(n_435) );
AND2x4_ASAP7_75t_L g559 ( .A(n_334), .B(n_345), .Y(n_559) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_339), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
BUFx8_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_343), .Y(n_529) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x4_ASAP7_75t_L g348 ( .A(n_344), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g390 ( .A(n_344), .B(n_366), .Y(n_390) );
AND2x2_ASAP7_75t_L g395 ( .A(n_344), .B(n_362), .Y(n_395) );
AND2x2_ASAP7_75t_L g414 ( .A(n_344), .B(n_345), .Y(n_414) );
AND2x2_ASAP7_75t_L g425 ( .A(n_344), .B(n_366), .Y(n_425) );
AND2x4_ASAP7_75t_L g434 ( .A(n_344), .B(n_362), .Y(n_434) );
AND2x4_ASAP7_75t_L g555 ( .A(n_344), .B(n_345), .Y(n_555) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_347), .Y(n_643) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_348), .Y(n_415) );
BUFx3_ASAP7_75t_L g459 ( .A(n_348), .Y(n_459) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_348), .Y(n_489) );
BUFx12f_ASAP7_75t_L g534 ( .A(n_348), .Y(n_534) );
BUFx12f_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g758 ( .A(n_352), .Y(n_758) );
BUFx12f_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_353), .Y(n_456) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_353), .Y(n_647) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g417 ( .A(n_355), .Y(n_417) );
INVx4_ASAP7_75t_L g457 ( .A(n_355), .Y(n_457) );
INVx2_ASAP7_75t_L g491 ( .A(n_355), .Y(n_491) );
INVx1_ASAP7_75t_L g654 ( .A(n_355), .Y(n_654) );
INVx4_ASAP7_75t_L g678 ( .A(n_355), .Y(n_678) );
INVx2_ASAP7_75t_L g731 ( .A(n_355), .Y(n_731) );
INVx8_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx4f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g729 ( .A(n_360), .Y(n_729) );
INVx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_361), .Y(n_451) );
BUFx12f_ASAP7_75t_L g493 ( .A(n_361), .Y(n_493) );
AND2x4_ASAP7_75t_L g371 ( .A(n_362), .B(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g497 ( .A(n_362), .B(n_372), .Y(n_497) );
AND2x4_ASAP7_75t_L g366 ( .A(n_363), .B(n_367), .Y(n_366) );
BUFx3_ASAP7_75t_L g650 ( .A(n_364), .Y(n_650) );
BUFx5_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g454 ( .A(n_365), .Y(n_454) );
BUFx3_ASAP7_75t_L g494 ( .A(n_365), .Y(n_494) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_365), .Y(n_532) );
AND2x4_ASAP7_75t_L g386 ( .A(n_366), .B(n_372), .Y(n_386) );
AND2x2_ASAP7_75t_L g605 ( .A(n_366), .B(n_372), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g368 ( .A(n_369), .B(n_383), .C(n_391), .D(n_398), .Y(n_368) );
INVx4_ASAP7_75t_L g522 ( .A(n_370), .Y(n_522) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g431 ( .A(n_371), .Y(n_431) );
BUFx3_ASAP7_75t_L g628 ( .A(n_371), .Y(n_628) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g477 ( .A(n_374), .Y(n_477) );
INVx4_ASAP7_75t_L g713 ( .A(n_374), .Y(n_713) );
INVx2_ASAP7_75t_L g1026 ( .A(n_374), .Y(n_1026) );
INVx5_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g504 ( .A(n_375), .Y(n_504) );
BUFx4f_ASAP7_75t_L g524 ( .A(n_375), .Y(n_524) );
AND2x4_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
AND2x2_ASAP7_75t_L g432 ( .A(n_376), .B(n_380), .Y(n_432) );
AND2x4_ASAP7_75t_L g583 ( .A(n_376), .B(n_380), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g470 ( .A(n_385), .Y(n_470) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_386), .Y(n_421) );
BUFx3_ASAP7_75t_L g536 ( .A(n_386), .Y(n_536) );
BUFx8_ASAP7_75t_SL g563 ( .A(n_386), .Y(n_563) );
INVx1_ASAP7_75t_L g709 ( .A(n_387), .Y(n_709) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g768 ( .A(n_389), .Y(n_768) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx3_ASAP7_75t_L g475 ( .A(n_390), .Y(n_475) );
INVx2_ASAP7_75t_L g539 ( .A(n_390), .Y(n_539) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g478 ( .A(n_393), .Y(n_478) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_393), .Y(n_754) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g703 ( .A(n_394), .Y(n_703) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx3_ASAP7_75t_L g505 ( .A(n_395), .Y(n_505) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_395), .Y(n_516) );
INVx3_ASAP7_75t_L g518 ( .A(n_396), .Y(n_518) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_397), .Y(n_471) );
INVx3_ASAP7_75t_L g706 ( .A(n_397), .Y(n_706) );
INVx2_ASAP7_75t_SL g715 ( .A(n_399), .Y(n_715) );
INVx2_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_400), .Y(n_427) );
INVx1_ASAP7_75t_L g737 ( .A(n_400), .Y(n_737) );
INVx2_ASAP7_75t_L g1031 ( .A(n_400), .Y(n_1031) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx3_ASAP7_75t_L g468 ( .A(n_401), .Y(n_468) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_406), .Y(n_401) );
HB1xp67_ASAP7_75t_L g778 ( .A(n_403), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND4xp75_ASAP7_75t_L g410 ( .A(n_411), .B(n_418), .C(n_429), .D(n_436), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx4f_ASAP7_75t_L g488 ( .A(n_414), .Y(n_488) );
OA21x2_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_422), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_420), .A2(n_518), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_427), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_433), .Y(n_429) );
INVx2_ASAP7_75t_L g586 ( .A(n_434), .Y(n_586) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_444), .Y(n_506) );
AO22x2_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_479), .B2(n_480), .Y(n_444) );
INVx2_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
XNOR2x1_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_461), .Y(n_448) );
NAND4xp25_ASAP7_75t_L g449 ( .A(n_450), .B(n_455), .C(n_458), .D(n_460), .Y(n_449) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .C(n_476), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_464), .B(n_469), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_467), .B(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_467), .B(n_577), .Y(n_576) );
INVx4_ASAP7_75t_L g639 ( .A(n_467), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_467), .B(n_687), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_467), .B(n_1049), .Y(n_1048) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx4_ASAP7_75t_L g544 ( .A(n_468), .Y(n_544) );
BUFx3_ASAP7_75t_L g625 ( .A(n_471), .Y(n_625) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g502 ( .A(n_475), .Y(n_502) );
INVx3_ASAP7_75t_SL g1021 ( .A(n_475), .Y(n_1021) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
HB1xp67_ASAP7_75t_SL g692 ( .A(n_480), .Y(n_692) );
INVx2_ASAP7_75t_L g719 ( .A(n_480), .Y(n_719) );
NOR2x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_495), .Y(n_481) );
NAND4xp25_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .C(n_490), .D(n_492), .Y(n_482) );
INVx5_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g745 ( .A(n_486), .Y(n_745) );
BUFx2_ASAP7_75t_L g762 ( .A(n_494), .Y(n_762) );
NAND4xp25_ASAP7_75t_SL g495 ( .A(n_496), .B(n_500), .C(n_501), .D(n_503), .Y(n_495) );
INVx2_ASAP7_75t_L g630 ( .A(n_505), .Y(n_630) );
XNOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_568), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
XNOR2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_545), .Y(n_510) );
NAND4xp75_ASAP7_75t_L g512 ( .A(n_513), .B(n_525), .C(n_530), .D(n_535), .Y(n_512) );
NOR2xp67_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_517), .B1(n_518), .B2(n_519), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_523), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_522), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
INVx2_ASAP7_75t_SL g636 ( .A(n_524), .Y(n_636) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_528), .Y(n_525) );
BUFx3_ASAP7_75t_L g648 ( .A(n_527), .Y(n_648) );
BUFx3_ASAP7_75t_L g652 ( .A(n_529), .Y(n_652) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_533), .Y(n_530) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g634 ( .A(n_538), .Y(n_634) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g662 ( .A(n_539), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_544), .B(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_544), .B(n_667), .Y(n_666) );
XOR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_567), .Y(n_545) );
NOR4xp75_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .C(n_553), .D(n_560), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_554), .B(n_557), .Y(n_553) );
OAI21x1_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_562), .B(n_564), .Y(n_560) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_563), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_595), .B1(n_613), .B2(n_614), .Y(n_568) );
INVx1_ASAP7_75t_L g613 ( .A(n_569), .Y(n_613) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g594 ( .A(n_573), .Y(n_594) );
NOR2x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_588), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_578), .C(n_587), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B1(n_584), .B2(n_586), .Y(n_579) );
CKINVDCx16_ASAP7_75t_R g580 ( .A(n_581), .Y(n_580) );
INVx4_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
CKINVDCx9p33_ASAP7_75t_R g584 ( .A(n_585), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .C(n_591), .D(n_592), .Y(n_588) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_597), .Y(n_615) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_608), .Y(n_599) );
NAND4xp25_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .C(n_603), .D(n_604), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .C(n_611), .D(n_612), .Y(n_608) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B1(n_689), .B2(n_770), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_655), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_641), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .C(n_631), .Y(n_622) );
BUFx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_640), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND4xp25_ASAP7_75t_SL g641 ( .A(n_642), .B(n_645), .C(n_649), .D(n_651), .Y(n_641) );
BUFx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
XNOR2x1_ASAP7_75t_L g656 ( .A(n_657), .B(n_673), .Y(n_656) );
XNOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .Y(n_657) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_668), .Y(n_659) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .C(n_664), .D(n_665), .Y(n_660) );
NAND4xp25_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .C(n_671), .D(n_672), .Y(n_668) );
XNOR2x1_ASAP7_75t_L g673 ( .A(n_674), .B(n_688), .Y(n_673) );
NAND4xp75_ASAP7_75t_L g674 ( .A(n_675), .B(n_679), .C(n_682), .D(n_685), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g770 ( .A(n_689), .Y(n_770) );
XNOR2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_721), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_716), .B2(n_720), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx2_ASAP7_75t_SL g720 ( .A(n_693), .Y(n_720) );
NAND4xp75_ASAP7_75t_SL g694 ( .A(n_695), .B(n_698), .C(n_701), .D(n_707), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx3_ASAP7_75t_L g1023 ( .A(n_706), .Y(n_1023) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_712), .B1(n_714), .B2(n_715), .Y(n_710) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B1(n_739), .B2(n_740), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
XOR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_738), .Y(n_723) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_725), .B(n_732), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .C(n_728), .D(n_730), .Y(n_725) );
NAND4xp25_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .C(n_735), .D(n_736), .Y(n_732) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND4xp75_ASAP7_75t_L g741 ( .A(n_742), .B(n_747), .C(n_755), .D(n_763), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_746), .Y(n_742) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NOR2x1_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .Y(n_747) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_761), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
BUFx3_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI21xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_769), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx3_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
HB1xp67_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND3xp33_ASAP7_75t_L g774 ( .A(n_775), .B(n_778), .C(n_779), .Y(n_774) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_775), .B(n_1035), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_775), .B(n_1036), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_775), .A2(n_779), .B(n_789), .Y(n_1060) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
AO21x1_ASAP7_75t_L g1058 ( .A1(n_776), .A2(n_1059), .B(n_1060), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
AND3x4_ASAP7_75t_L g786 ( .A(n_777), .B(n_787), .C(n_789), .Y(n_786) );
AND2x2_ASAP7_75t_L g794 ( .A(n_777), .B(n_795), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g1035 ( .A(n_778), .B(n_1036), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_779), .Y(n_1036) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_1004), .B1(n_1007), .B2(n_1033), .C(n_1037), .Y(n_780) );
AOI211x1_ASAP7_75t_SL g781 ( .A1(n_782), .A2(n_860), .B(n_874), .C(n_982), .Y(n_781) );
OAI211xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_803), .B(n_829), .C(n_849), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_798), .Y(n_783) );
INVx1_ASAP7_75t_L g834 ( .A(n_784), .Y(n_834) );
OR2x2_ASAP7_75t_L g852 ( .A(n_784), .B(n_835), .Y(n_852) );
AND2x2_ASAP7_75t_L g891 ( .A(n_784), .B(n_835), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_784), .B(n_799), .Y(n_910) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_792), .Y(n_784) );
AND2x4_ASAP7_75t_L g790 ( .A(n_787), .B(n_791), .Y(n_790) );
AND2x4_ASAP7_75t_L g808 ( .A(n_787), .B(n_794), .Y(n_808) );
AND2x4_ASAP7_75t_L g809 ( .A(n_787), .B(n_791), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_787), .B(n_791), .Y(n_818) );
AND2x2_ASAP7_75t_L g797 ( .A(n_791), .B(n_796), .Y(n_797) );
AND2x4_ASAP7_75t_L g801 ( .A(n_791), .B(n_796), .Y(n_801) );
AND2x2_ASAP7_75t_L g812 ( .A(n_791), .B(n_796), .Y(n_812) );
AND2x2_ASAP7_75t_L g793 ( .A(n_794), .B(n_796), .Y(n_793) );
AND2x2_ASAP7_75t_L g811 ( .A(n_794), .B(n_796), .Y(n_811) );
AND2x4_ASAP7_75t_L g822 ( .A(n_794), .B(n_796), .Y(n_822) );
NOR2x1_ASAP7_75t_R g846 ( .A(n_798), .B(n_847), .Y(n_846) );
AND2x2_ASAP7_75t_L g887 ( .A(n_798), .B(n_833), .Y(n_887) );
AND2x2_ASAP7_75t_L g905 ( .A(n_798), .B(n_834), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_798), .B(n_939), .Y(n_938) );
AND2x2_ASAP7_75t_L g952 ( .A(n_798), .B(n_891), .Y(n_952) );
AND2x2_ASAP7_75t_L g979 ( .A(n_798), .B(n_943), .Y(n_979) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_SL g832 ( .A(n_799), .Y(n_832) );
AND2x2_ASAP7_75t_L g843 ( .A(n_799), .B(n_844), .Y(n_843) );
OR2x2_ASAP7_75t_L g880 ( .A(n_799), .B(n_845), .Y(n_880) );
AND2x2_ASAP7_75t_L g942 ( .A(n_799), .B(n_943), .Y(n_942) );
OR2x2_ASAP7_75t_L g972 ( .A(n_799), .B(n_852), .Y(n_972) );
AND2x2_ASAP7_75t_L g984 ( .A(n_799), .B(n_834), .Y(n_984) );
AND2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
INVx2_ASAP7_75t_L g824 ( .A(n_801), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_804), .B(n_813), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_804), .B(n_905), .Y(n_904) );
NAND2xp67_ASAP7_75t_L g1002 ( .A(n_804), .B(n_830), .Y(n_1002) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
NOR2x1_ASAP7_75t_L g844 ( .A(n_805), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_SL g847 ( .A(n_805), .B(n_848), .Y(n_847) );
BUFx6f_ASAP7_75t_L g858 ( .A(n_805), .Y(n_858) );
INVx2_ASAP7_75t_L g879 ( .A(n_805), .Y(n_879) );
INVx1_ASAP7_75t_L g893 ( .A(n_805), .Y(n_893) );
AND2x2_ASAP7_75t_L g935 ( .A(n_805), .B(n_814), .Y(n_935) );
AND2x2_ASAP7_75t_L g941 ( .A(n_805), .B(n_942), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_805), .B(n_884), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_805), .B(n_905), .Y(n_962) );
AND2x2_ASAP7_75t_L g970 ( .A(n_805), .B(n_882), .Y(n_970) );
INVx4_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_806), .B(n_841), .Y(n_911) );
OR2x2_ASAP7_75t_L g915 ( .A(n_806), .B(n_831), .Y(n_915) );
AND2x2_ASAP7_75t_L g930 ( .A(n_806), .B(n_814), .Y(n_930) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_810), .Y(n_806) );
INVx3_ASAP7_75t_L g816 ( .A(n_808), .Y(n_816) );
INVx1_ASAP7_75t_L g917 ( .A(n_813), .Y(n_917) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_826), .Y(n_813) );
INVx2_ASAP7_75t_L g841 ( .A(n_814), .Y(n_841) );
INVx1_ASAP7_75t_L g882 ( .A(n_814), .Y(n_882) );
OR2x2_ASAP7_75t_L g924 ( .A(n_814), .B(n_826), .Y(n_924) );
AND2x2_ASAP7_75t_L g976 ( .A(n_814), .B(n_931), .Y(n_976) );
OR2x2_ASAP7_75t_L g814 ( .A(n_815), .B(n_820), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_816), .A2(n_817), .B1(n_818), .B2(n_819), .Y(n_815) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_816), .A2(n_818), .B1(n_865), .B2(n_866), .C(n_867), .Y(n_864) );
INVx1_ASAP7_75t_L g1006 ( .A(n_816), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_823), .B1(n_824), .B2(n_825), .Y(n_820) );
INVx3_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
OR2x2_ASAP7_75t_L g854 ( .A(n_826), .B(n_841), .Y(n_854) );
AND2x2_ASAP7_75t_L g859 ( .A(n_826), .B(n_841), .Y(n_859) );
HB1xp67_ASAP7_75t_L g894 ( .A(n_826), .Y(n_894) );
OR2x2_ASAP7_75t_L g898 ( .A(n_826), .B(n_870), .Y(n_898) );
AND2x2_ASAP7_75t_L g907 ( .A(n_826), .B(n_869), .Y(n_907) );
OR2x2_ASAP7_75t_L g926 ( .A(n_826), .B(n_871), .Y(n_926) );
AND2x2_ASAP7_75t_L g931 ( .A(n_826), .B(n_870), .Y(n_931) );
INVx2_ASAP7_75t_L g958 ( .A(n_826), .Y(n_958) );
AND2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_838), .B1(n_839), .B2(n_846), .Y(n_829) );
INVx1_ASAP7_75t_L g916 ( .A(n_830), .Y(n_916) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_833), .Y(n_830) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_831), .A2(n_850), .B1(n_853), .B2(n_855), .Y(n_849) );
AND2x4_ASAP7_75t_L g850 ( .A(n_831), .B(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g890 ( .A(n_831), .B(n_891), .Y(n_890) );
AND2x2_ASAP7_75t_L g903 ( .A(n_831), .B(n_835), .Y(n_903) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
AOI211xp5_ASAP7_75t_L g899 ( .A1(n_833), .A2(n_900), .B(n_901), .C(n_912), .Y(n_899) );
INVx1_ASAP7_75t_L g967 ( .A(n_833), .Y(n_967) );
AND2x2_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
OR2x2_ASAP7_75t_L g845 ( .A(n_834), .B(n_835), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_834), .B(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g943 ( .A(n_835), .Y(n_943) );
AOI222xp33_ASAP7_75t_L g991 ( .A1(n_835), .A2(n_859), .B1(n_992), .B2(n_993), .C1(n_995), .C2(n_996), .Y(n_991) );
AND2x2_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_842), .Y(n_838) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_839), .B(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g896 ( .A(n_840), .B(n_897), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_840), .B(n_903), .Y(n_902) );
A2O1A1Ixp33_ASAP7_75t_L g999 ( .A1(n_840), .A2(n_1000), .B(n_1001), .C(n_1003), .Y(n_999) );
NOR2xp67_ASAP7_75t_SL g1001 ( .A(n_840), .B(n_1002), .Y(n_1001) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g954 ( .A(n_841), .B(n_884), .Y(n_954) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx3_ASAP7_75t_SL g848 ( .A(n_845), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_848), .B(n_914), .Y(n_955) );
AOI221xp5_ASAP7_75t_L g983 ( .A1(n_848), .A2(n_900), .B1(n_984), .B2(n_985), .C(n_986), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_850), .B(n_878), .Y(n_877) );
INVx2_ASAP7_75t_SL g897 ( .A(n_850), .Y(n_897) );
AND2x2_ASAP7_75t_L g995 ( .A(n_850), .B(n_879), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_851), .B(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_852), .B(n_933), .Y(n_939) );
AND2x2_ASAP7_75t_L g900 ( .A(n_853), .B(n_883), .Y(n_900) );
AOI321xp33_ASAP7_75t_L g946 ( .A1(n_853), .A2(n_947), .A3(n_948), .B1(n_949), .B2(n_951), .C(n_953), .Y(n_946) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_859), .Y(n_856) );
AND2x2_ASAP7_75t_L g975 ( .A(n_857), .B(n_952), .Y(n_975) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g919 ( .A1(n_858), .A2(n_920), .B1(n_925), .B2(n_926), .C(n_927), .Y(n_919) );
OAI321xp33_ASAP7_75t_L g937 ( .A1(n_858), .A2(n_926), .A3(n_938), .B1(n_940), .B2(n_944), .C(n_946), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_858), .B(n_859), .Y(n_997) );
AND2x2_ASAP7_75t_L g951 ( .A(n_859), .B(n_952), .Y(n_951) );
INVxp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_868), .Y(n_861) );
OAI31xp33_ASAP7_75t_L g875 ( .A1(n_862), .A2(n_876), .A3(n_885), .B(n_888), .Y(n_875) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
AOI211xp5_ASAP7_75t_L g918 ( .A1(n_863), .A2(n_919), .B(n_937), .C(n_956), .Y(n_918) );
AOI222xp33_ASAP7_75t_L g963 ( .A1(n_863), .A2(n_907), .B1(n_964), .B2(n_965), .C1(n_968), .C2(n_973), .Y(n_963) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g950 ( .A(n_864), .Y(n_950) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_864), .B(n_883), .Y(n_998) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g884 ( .A(n_871), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
NAND4xp25_ASAP7_75t_L g874 ( .A(n_875), .B(n_918), .C(n_963), .D(n_974), .Y(n_874) );
AOI21xp33_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_880), .B(n_881), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_878), .B(n_890), .Y(n_960) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_879), .B(n_887), .Y(n_886) );
INVx1_ASAP7_75t_L g1000 ( .A(n_880), .Y(n_1000) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
INVx2_ASAP7_75t_L g945 ( .A(n_882), .Y(n_945) );
OAI322xp33_ASAP7_75t_L g986 ( .A1(n_882), .A2(n_933), .A3(n_943), .B1(n_966), .B2(n_987), .C1(n_988), .C2(n_990), .Y(n_986) );
INVx1_ASAP7_75t_L g973 ( .A(n_883), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g990 ( .A(n_883), .B(n_970), .Y(n_990) );
INVx2_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx3_ASAP7_75t_L g922 ( .A(n_884), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g985 ( .A(n_884), .B(n_924), .Y(n_985) );
NOR2xp33_ASAP7_75t_L g889 ( .A(n_887), .B(n_890), .Y(n_889) );
AOI321xp33_ASAP7_75t_L g974 ( .A1(n_887), .A2(n_950), .A3(n_958), .B1(n_975), .B2(n_976), .C(n_977), .Y(n_974) );
OAI221xp5_ASAP7_75t_SL g888 ( .A1(n_889), .A2(n_892), .B1(n_895), .B2(n_898), .C(n_899), .Y(n_888) );
INVx1_ASAP7_75t_L g925 ( .A(n_890), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_891), .B(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g933 ( .A(n_891), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_893), .B(n_924), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g908 ( .A(n_894), .B(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g994 ( .A(n_894), .Y(n_994) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
O2A1O1Ixp33_ASAP7_75t_L g953 ( .A1(n_898), .A2(n_950), .B(n_954), .C(n_955), .Y(n_953) );
A2O1A1Ixp33_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_904), .B(n_906), .C(n_908), .Y(n_901) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_907), .B(n_945), .Y(n_944) );
NOR2xp33_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
INVx1_ASAP7_75t_L g948 ( .A(n_910), .Y(n_948) );
AOI21xp33_ASAP7_75t_SL g912 ( .A1(n_913), .A2(n_916), .B(n_917), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OR2x2_ASAP7_75t_L g966 ( .A(n_915), .B(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g961 ( .A(n_921), .Y(n_961) );
AND2x2_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
INVx2_ASAP7_75t_L g936 ( .A(n_922), .Y(n_936) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
AOI21xp33_ASAP7_75t_L g977 ( .A1(n_925), .A2(n_978), .B(n_980), .Y(n_977) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_928), .A2(n_931), .B(n_932), .Y(n_927) );
INVxp67_ASAP7_75t_SL g928 ( .A(n_929), .Y(n_928) );
NOR3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_934), .C(n_936), .Y(n_932) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_945), .B(n_960), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_945), .B(n_966), .Y(n_965) );
INVx1_ASAP7_75t_L g987 ( .A(n_947), .Y(n_987) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g959 ( .A(n_950), .Y(n_959) );
OAI221xp5_ASAP7_75t_SL g982 ( .A1(n_950), .A2(n_983), .B1(n_991), .B2(n_998), .C(n_999), .Y(n_982) );
OAI22xp5_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_960), .B1(n_961), .B2(n_962), .Y(n_956) );
INVxp67_ASAP7_75t_L g1003 ( .A(n_957), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
CKINVDCx14_ASAP7_75t_R g989 ( .A(n_958), .Y(n_989) );
INVx1_ASAP7_75t_L g992 ( .A(n_962), .Y(n_992) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g969 ( .A(n_970), .B(n_971), .Y(n_969) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
CKINVDCx14_ASAP7_75t_R g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVxp67_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_1005), .Y(n_1004) );
HB1xp67_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
HB1xp67_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
XNOR2x1_ASAP7_75t_L g1011 ( .A(n_1012), .B(n_1032), .Y(n_1011) );
NAND4xp75_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1016), .C(n_1019), .D(n_1024), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1015), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_1017), .B(n_1018), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1022), .Y(n_1019) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1027), .Y(n_1024) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .Y(n_1028) );
INVx3_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
BUFx2_ASAP7_75t_SL g1038 ( .A(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1042), .Y(n_1056) );
INVxp33_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
NOR2x1_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1051), .Y(n_1043) );
NAND4xp25_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1046), .C(n_1047), .D(n_1050), .Y(n_1044) );
NAND4xp25_ASAP7_75t_SL g1051 ( .A(n_1052), .B(n_1053), .C(n_1054), .D(n_1055), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
endmodule