module fake_jpeg_3682_n_534 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_534);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx12f_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx9p33_ASAP7_75t_R g104 ( 
.A(n_55),
.Y(n_104)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_56),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_60),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_77),
.Y(n_116)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_66),
.Y(n_103)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_83),
.Y(n_117)
);

BUFx3_ASAP7_75t_SL g80 ( 
.A(n_19),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g145 ( 
.A(n_80),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_27),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

BUFx24_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx5_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_31),
.B(n_7),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_98),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_28),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_99),
.B(n_28),
.Y(n_154)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_97),
.A2(n_39),
.B1(n_26),
.B2(n_40),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_101),
.A2(n_100),
.B1(n_25),
.B2(n_35),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_50),
.A2(n_40),
.B1(n_20),
.B2(n_43),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_114),
.A2(n_20),
.B1(n_79),
.B2(n_73),
.Y(n_165)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

INVx6_ASAP7_75t_SL g130 ( 
.A(n_80),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_40),
.B1(n_28),
.B2(n_43),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_92),
.B1(n_91),
.B2(n_90),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_80),
.B(n_37),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_140),
.B(n_157),
.Y(n_208)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_51),
.Y(n_150)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_95),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_80),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_57),
.Y(n_160)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_116),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_164),
.B(n_166),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_165),
.A2(n_174),
.B1(n_141),
.B2(n_125),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_89),
.Y(n_166)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_168),
.Y(n_228)
);

OR2x4_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_66),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_169),
.A2(n_189),
.B1(n_195),
.B2(n_196),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_61),
.C(n_93),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_183),
.C(n_192),
.Y(n_217)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

CKINVDCx12_ASAP7_75t_R g172 ( 
.A(n_103),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_172),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_60),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_176),
.B(n_180),
.Y(n_222)
);

BUFx8_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_179),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_21),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_162),
.Y(n_182)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_113),
.B(n_81),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_109),
.B(n_31),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_184),
.B(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_112),
.Y(n_187)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_109),
.B(n_37),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_95),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_116),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_155),
.Y(n_194)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

CKINVDCx12_ASAP7_75t_R g195 ( 
.A(n_103),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_117),
.B(n_147),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_102),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_143),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_34),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_200),
.A2(n_203),
.B1(n_210),
.B2(n_211),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_110),
.B(n_34),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_25),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_205),
.B1(n_101),
.B2(n_155),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_134),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_136),
.A2(n_68),
.B1(n_58),
.B2(n_44),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_131),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_131),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_207),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_105),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

CKINVDCx12_ASAP7_75t_R g210 ( 
.A(n_145),
.Y(n_210)
);

NAND2x1_ASAP7_75t_SL g211 ( 
.A(n_137),
.B(n_25),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_239),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_230),
.B(n_235),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_126),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_234),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_174),
.A2(n_205),
.B1(n_114),
.B2(n_202),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_120),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_180),
.A2(n_141),
.B1(n_125),
.B2(n_159),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_244),
.B(n_248),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_107),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_169),
.Y(n_251)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_163),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g249 ( 
.A(n_223),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_249),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_171),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_250),
.B(n_254),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_275),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

INVx8_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_253),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_204),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_245),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_257),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_203),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_216),
.A2(n_170),
.B1(n_135),
.B2(n_149),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_264),
.B1(n_270),
.B2(n_276),
.Y(n_280)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_236),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_260),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_230),
.A2(n_183),
.B1(n_132),
.B2(n_108),
.Y(n_264)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_236),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_265),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_217),
.B(n_192),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_214),
.C(n_218),
.Y(n_285)
);

O2A1O1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_211),
.B(n_178),
.C(n_175),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_268),
.A2(n_221),
.B(n_226),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_269),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_225),
.A2(n_151),
.B1(n_182),
.B2(n_209),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_225),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_234),
.A2(n_159),
.B1(n_119),
.B2(n_118),
.Y(n_276)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_237),
.Y(n_310)
);

NOR2x1_ASAP7_75t_R g279 ( 
.A(n_244),
.B(n_178),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_194),
.B(n_122),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_232),
.B1(n_217),
.B2(n_229),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_286),
.B1(n_287),
.B2(n_301),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_261),
.A2(n_255),
.B1(n_273),
.B2(n_258),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_290),
.C(n_291),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_255),
.A2(n_229),
.B1(n_214),
.B2(n_241),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_255),
.A2(n_213),
.B1(n_215),
.B2(n_226),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_215),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_251),
.B(n_213),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_248),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g330 ( 
.A(n_296),
.B(n_298),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_272),
.B(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_299),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_269),
.A2(n_119),
.B1(n_181),
.B2(n_106),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_259),
.A2(n_156),
.B1(n_161),
.B2(n_106),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_272),
.A2(n_118),
.B1(n_173),
.B2(n_144),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_305),
.B1(n_309),
.B2(n_311),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_276),
.A2(n_275),
.B1(n_279),
.B2(n_264),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_266),
.B(n_246),
.Y(n_306)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

AOI22x1_ASAP7_75t_L g309 ( 
.A1(n_268),
.A2(n_237),
.B1(n_233),
.B2(n_227),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_266),
.A2(n_144),
.B1(n_163),
.B2(n_167),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_252),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_313),
.B(n_315),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_227),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_221),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_329),
.Y(n_349)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_319),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_293),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_322),
.Y(n_378)
);

AO22x1_ASAP7_75t_L g322 ( 
.A1(n_283),
.A2(n_274),
.B1(n_271),
.B2(n_278),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_285),
.C(n_282),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_326),
.C(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_324),
.Y(n_356)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_325),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_271),
.C(n_274),
.Y(n_326)
);

OR2x2_ASAP7_75t_SL g327 ( 
.A(n_292),
.B(n_249),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_327),
.A2(n_289),
.B(n_249),
.Y(n_352)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_328),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_311),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_289),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_334),
.Y(n_359)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_332),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_281),
.Y(n_335)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_335),
.Y(n_365)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_304),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_337),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_284),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_338),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_292),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_309),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_301),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_307),
.B(n_249),
.Y(n_342)
);

NOR3xp33_ASAP7_75t_SL g363 ( 
.A(n_342),
.B(n_343),
.C(n_238),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_305),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_298),
.B(n_278),
.C(n_233),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_240),
.C(n_197),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_314),
.A2(n_280),
.B1(n_295),
.B2(n_303),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_346),
.A2(n_376),
.B1(n_333),
.B2(n_329),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_334),
.A2(n_295),
.B(n_280),
.Y(n_347)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_350),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_338),
.B(n_343),
.Y(n_350)
);

NAND2xp67_ASAP7_75t_SL g385 ( 
.A(n_352),
.B(n_327),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_353),
.B(n_199),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_299),
.B(n_260),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_355),
.A2(n_367),
.B(n_371),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_340),
.A2(n_302),
.B1(n_294),
.B2(n_253),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_358),
.A2(n_362),
.B1(n_368),
.B2(n_377),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_337),
.A2(n_302),
.B1(n_294),
.B2(n_262),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_364),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_265),
.B(n_220),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_323),
.B(n_243),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_375),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_314),
.A2(n_321),
.B(n_322),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_325),
.A2(n_263),
.B1(n_262),
.B2(n_220),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_342),
.A2(n_206),
.B(n_207),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_335),
.C(n_332),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_322),
.A2(n_240),
.B(n_228),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_35),
.B(n_22),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_177),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_324),
.A2(n_277),
.B1(n_263),
.B2(n_187),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_185),
.B1(n_177),
.B2(n_167),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_365),
.Y(n_379)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_379),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_382),
.C(n_390),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_381),
.A2(n_383),
.B1(n_357),
.B2(n_356),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_320),
.C(n_326),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_345),
.A2(n_312),
.B1(n_319),
.B2(n_318),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_317),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_385),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_370),
.B(n_375),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_387),
.B(n_397),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_370),
.B(n_328),
.C(n_312),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_317),
.C(n_341),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_392),
.A2(n_399),
.B(n_406),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_372),
.B(n_341),
.C(n_185),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_393),
.B(n_396),
.C(n_364),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_359),
.B(n_354),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_394),
.B(n_400),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_228),
.C(n_168),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_367),
.B(n_146),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_398),
.Y(n_422)
);

AOI21xp33_ASAP7_75t_L g399 ( 
.A1(n_350),
.A2(n_146),
.B(n_30),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_361),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_401),
.Y(n_411)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_349),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_402),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_403),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_115),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_404),
.B(n_407),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_378),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_408),
.B(n_378),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_352),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_419),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_391),
.A2(n_346),
.B1(n_345),
.B2(n_357),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_414),
.B(n_431),
.Y(n_455)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_415),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_44),
.B1(n_39),
.B2(n_42),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_382),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_138),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_390),
.C(n_380),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_423),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_389),
.B(n_374),
.C(n_362),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_397),
.B(n_371),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_424),
.B(n_429),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_358),
.C(n_355),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_426),
.B(n_427),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_368),
.C(n_353),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_383),
.B(n_363),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_393),
.B(n_385),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_386),
.B(n_353),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_432),
.B(n_42),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_381),
.A2(n_376),
.B1(n_44),
.B2(n_39),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_403),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_430),
.A2(n_395),
.B(n_386),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_438),
.A2(n_457),
.B(n_454),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_433),
.A2(n_395),
.B1(n_403),
.B2(n_405),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_439),
.A2(n_78),
.B1(n_41),
.B2(n_3),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_406),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_440),
.B(n_446),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_441),
.B(n_443),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_418),
.B(n_44),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_115),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_444),
.B(n_448),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_445),
.A2(n_454),
.B1(n_433),
.B2(n_422),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_413),
.B(n_30),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_412),
.A2(n_42),
.B(n_30),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_447),
.A2(n_457),
.B(n_432),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_35),
.C(n_138),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_411),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_449),
.B(n_409),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_138),
.C(n_21),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_416),
.C(n_424),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_429),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_426),
.A2(n_22),
.B1(n_21),
.B2(n_87),
.Y(n_454)
);

AOI221xp5_ASAP7_75t_L g456 ( 
.A1(n_423),
.A2(n_22),
.B1(n_13),
.B2(n_2),
.C(n_3),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_456),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_45),
.B(n_19),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_465),
.Y(n_486)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_450),
.B(n_419),
.C(n_427),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_467),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_461),
.Y(n_480)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_462),
.Y(n_484)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_464),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_435),
.B(n_420),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_455),
.A2(n_416),
.B(n_87),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_466),
.A2(n_475),
.B(n_47),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_437),
.A2(n_78),
.B1(n_41),
.B2(n_2),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_470),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_453),
.B(n_9),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_447),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_472),
.B(n_8),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_47),
.C(n_41),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_473),
.B(n_474),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_435),
.B(n_47),
.C(n_1),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_439),
.C(n_441),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_SL g495 ( 
.A(n_478),
.B(n_489),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_452),
.Y(n_479)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_479),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_481),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_451),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_490),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_442),
.C(n_445),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_442),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_491),
.A2(n_494),
.B1(n_467),
.B2(n_466),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_8),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_492),
.B(n_13),
.Y(n_501)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_480),
.B(n_458),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_498),
.B(n_503),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_464),
.B(n_462),
.Y(n_499)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_499),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_501),
.B(n_504),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_481),
.B(n_471),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_471),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_493),
.A2(n_468),
.B1(n_474),
.B2(n_473),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_505),
.A2(n_494),
.B1(n_492),
.B2(n_488),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_486),
.B(n_5),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_506),
.B(n_507),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_485),
.B(n_478),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_47),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_508),
.B(n_484),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_511),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_479),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_482),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_497),
.B(n_47),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_514),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_502),
.B(n_9),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_496),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_522),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_516),
.A2(n_505),
.B(n_508),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_518),
.B(n_515),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_524),
.Y(n_527)
);

AOI322xp5_ASAP7_75t_L g525 ( 
.A1(n_519),
.A2(n_510),
.A3(n_513),
.B1(n_47),
.B2(n_4),
.C1(n_9),
.C2(n_10),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_525),
.A2(n_528),
.B(n_4),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g528 ( 
.A1(n_521),
.A2(n_3),
.A3(n_4),
.B1(n_10),
.B2(n_14),
.C1(n_0),
.C2(n_1),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_529),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_4),
.C(n_10),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_527),
.B(n_530),
.Y(n_532)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_532),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_10),
.Y(n_534)
);


endmodule