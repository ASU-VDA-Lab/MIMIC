module fake_jpeg_1258_n_612 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_612);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_612;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_6),
.B(n_13),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_61),
.Y(n_139)
);

INVx2_ASAP7_75t_R g62 ( 
.A(n_39),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_62),
.B(n_116),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_63),
.B(n_73),
.Y(n_151)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_9),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_78),
.Y(n_127)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_71),
.Y(n_153)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_77),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_9),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_81),
.Y(n_161)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_87),
.Y(n_168)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_90),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_92),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_94),
.Y(n_207)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_21),
.B(n_11),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_120),
.Y(n_144)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_38),
.Y(n_99)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_28),
.Y(n_101)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_46),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_102),
.B(n_111),
.Y(n_173)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_18),
.Y(n_104)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_105),
.Y(n_160)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx6f_ASAP7_75t_SL g110 ( 
.A(n_47),
.Y(n_110)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_46),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_41),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_112),
.B(n_117),
.Y(n_193)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_31),
.Y(n_113)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

CKINVDCx6p67_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_60),
.Y(n_117)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_119),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_21),
.B(n_8),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_18),
.Y(n_121)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_122),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_50),
.Y(n_123)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_23),
.Y(n_124)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_124),
.Y(n_201)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_125),
.B(n_35),
.Y(n_195)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_28),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_126),
.B(n_59),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_123),
.A2(n_51),
.B1(n_53),
.B2(n_43),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_131),
.A2(n_133),
.B1(n_164),
.B2(n_167),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_87),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_132),
.B(n_135),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_65),
.A2(n_60),
.B1(n_43),
.B2(n_57),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_88),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_78),
.B(n_43),
.C(n_57),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_15),
.C(n_16),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_60),
.B1(n_57),
.B2(n_51),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_143),
.A2(n_147),
.B1(n_174),
.B2(n_188),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_53),
.B1(n_59),
.B2(n_50),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_58),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_154),
.B(n_202),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_162),
.B(n_195),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_62),
.A2(n_50),
.B1(n_59),
.B2(n_27),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_74),
.A2(n_24),
.B1(n_26),
.B2(n_40),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_77),
.A2(n_24),
.B1(n_26),
.B2(n_40),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_178),
.B1(n_180),
.B2(n_190),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g174 ( 
.A1(n_84),
.A2(n_27),
.B1(n_19),
.B2(n_56),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_177),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_91),
.A2(n_19),
.B1(n_58),
.B2(n_56),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_61),
.A2(n_59),
.B1(n_50),
.B2(n_52),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_122),
.A2(n_107),
.B1(n_115),
.B2(n_94),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_92),
.A2(n_55),
.B1(n_44),
.B2(n_52),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_61),
.A2(n_35),
.B1(n_33),
.B2(n_44),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_205),
.B1(n_90),
.B2(n_82),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_89),
.B(n_55),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_89),
.B(n_12),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_134),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_79),
.A2(n_47),
.B1(n_32),
.B2(n_2),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_208),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_144),
.A2(n_100),
.B1(n_99),
.B2(n_109),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_210),
.B(n_251),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_127),
.B(n_0),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_211),
.B(n_214),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_157),
.B(n_116),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_215),
.Y(n_319)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_139),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_217),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_141),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_218),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_194),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_219),
.B(n_226),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_159),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

BUFx2_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_221),
.Y(n_291)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_174),
.Y(n_223)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_223),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_116),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_229),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_105),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_228),
.B(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_105),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_230),
.A2(n_234),
.B1(n_239),
.B2(n_279),
.Y(n_297)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_193),
.Y(n_231)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_231),
.Y(n_304)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_232),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_151),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_233),
.B(n_240),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_93),
.B1(n_114),
.B2(n_3),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_129),
.B(n_93),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_235),
.B(n_253),
.Y(n_292)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_237),
.Y(n_330)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_238),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_177),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_173),
.Y(n_240)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_169),
.Y(n_242)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_242),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_141),
.Y(n_243)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_143),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_244),
.A2(n_247),
.B1(n_270),
.B2(n_205),
.Y(n_287)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_168),
.Y(n_245)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_246),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_178),
.A2(n_7),
.B1(n_8),
.B2(n_12),
.Y(n_247)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_138),
.Y(n_248)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_248),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_7),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_164),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_256),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_7),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_185),
.Y(n_252)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_252),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_130),
.B(n_13),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_14),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_254),
.B(n_258),
.Y(n_309)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_255),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_149),
.B(n_14),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_261),
.C(n_150),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_140),
.B(n_14),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_180),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_260),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_206),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_146),
.B(n_15),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_262),
.B(n_265),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_142),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_263),
.B(n_267),
.Y(n_306)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_155),
.Y(n_264)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_264),
.Y(n_339)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_188),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_206),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_136),
.B(n_15),
.Y(n_267)
);

A2O1A1Ixp33_ASAP7_75t_L g268 ( 
.A1(n_156),
.A2(n_16),
.B(n_17),
.C(n_192),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_268),
.B(n_145),
.Y(n_325)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_271),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_152),
.A2(n_207),
.B1(n_187),
.B2(n_186),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_153),
.B(n_128),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_273),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_128),
.B(n_158),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_274),
.B(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_165),
.B(n_159),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g276 ( 
.A(n_134),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_277),
.Y(n_331)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_191),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_278),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_160),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_160),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_280),
.A2(n_150),
.B1(n_138),
.B2(n_172),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_287),
.A2(n_238),
.B1(n_277),
.B2(n_278),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_266),
.A2(n_152),
.B1(n_187),
.B2(n_186),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_296),
.A2(n_302),
.B1(n_310),
.B2(n_218),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_209),
.A2(n_131),
.B1(n_204),
.B2(n_199),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_298),
.A2(n_313),
.B1(n_324),
.B2(n_228),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_222),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_300),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_210),
.A2(n_176),
.B1(n_204),
.B2(n_199),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_249),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_307),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_305),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_249),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_223),
.A2(n_166),
.B1(n_207),
.B2(n_148),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_265),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_209),
.A2(n_176),
.B1(n_166),
.B2(n_148),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_251),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_315),
.B(n_276),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_241),
.B(n_172),
.C(n_163),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_322),
.B(n_329),
.C(n_333),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_250),
.A2(n_163),
.B1(n_138),
.B2(n_145),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_326),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_211),
.B(n_253),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_257),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_214),
.B(n_229),
.C(n_225),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_259),
.A2(n_212),
.B1(n_224),
.B2(n_228),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_213),
.B(n_236),
.Y(n_333)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_314),
.Y(n_340)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_295),
.A2(n_258),
.B1(n_262),
.B2(n_254),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_341),
.A2(n_345),
.B1(n_367),
.B2(n_373),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_235),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_342),
.B(n_363),
.C(n_374),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_333),
.B(n_251),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_343),
.B(n_344),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_300),
.B(n_257),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_346),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_348),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_309),
.B(n_261),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_309),
.B(n_232),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_350),
.B(n_371),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_304),
.B(n_321),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_351),
.B(n_380),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_294),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_368),
.Y(n_385)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_314),
.Y(n_353)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_355),
.A2(n_362),
.B1(n_375),
.B2(n_381),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_285),
.A2(n_268),
.B(n_221),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_357),
.A2(n_369),
.B(n_354),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_335),
.Y(n_360)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_360),
.Y(n_416)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_361),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_269),
.B1(n_245),
.B2(n_272),
.Y(n_362)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_299),
.Y(n_364)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_364),
.Y(n_392)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_283),
.Y(n_365)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_316),
.A2(n_237),
.B1(n_255),
.B2(n_264),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_331),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_286),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_291),
.Y(n_393)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_283),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_370),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_208),
.Y(n_371)
);

AO21x2_ASAP7_75t_L g372 ( 
.A1(n_298),
.A2(n_215),
.B(n_220),
.Y(n_372)
);

AO21x1_ASAP7_75t_L g395 ( 
.A1(n_372),
.A2(n_310),
.B(n_282),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_316),
.A2(n_243),
.B1(n_216),
.B2(n_242),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_279),
.C(n_280),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_316),
.A2(n_248),
.B1(n_252),
.B2(n_217),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_292),
.B(n_246),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_376),
.B(n_320),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_289),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_377),
.Y(n_387)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_312),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_378),
.B(n_382),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_311),
.B(n_288),
.C(n_292),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_281),
.C(n_301),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_295),
.A2(n_276),
.B1(n_326),
.B2(n_288),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_325),
.A2(n_306),
.B(n_284),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_383),
.A2(n_338),
.B(n_318),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_390),
.A2(n_398),
.B(n_400),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g437 ( 
.A(n_393),
.B(n_399),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_372),
.A2(n_296),
.B1(n_315),
.B2(n_307),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_394),
.A2(n_417),
.B1(n_423),
.B2(n_378),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_395),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_320),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_397),
.B(n_406),
.C(n_407),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_354),
.A2(n_297),
.B(n_308),
.Y(n_398)
);

HAxp5_ASAP7_75t_SL g399 ( 
.A(n_358),
.B(n_327),
.CON(n_399),
.SN(n_399)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_357),
.A2(n_303),
.B(n_323),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_349),
.A2(n_322),
.B(n_324),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_401),
.A2(n_398),
.B(n_422),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_363),
.B(n_366),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_281),
.Y(n_407)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_374),
.C(n_342),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_352),
.B(n_304),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_411),
.B(n_415),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_384),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_414),
.B(n_360),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_371),
.B(n_339),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_372),
.A2(n_281),
.B1(n_282),
.B2(n_301),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_381),
.A2(n_339),
.B(n_338),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_421),
.A2(n_422),
.B(n_293),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_372),
.A2(n_317),
.B1(n_334),
.B2(n_330),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_SL g483 ( 
.A(n_424),
.B(n_427),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_390),
.A2(n_356),
.B(n_383),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_409),
.Y(n_428)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_428),
.Y(n_463)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_402),
.Y(n_429)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_429),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_433),
.C(n_438),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_417),
.A2(n_349),
.B(n_368),
.Y(n_431)
);

OAI21xp33_ASAP7_75t_L g476 ( 
.A1(n_431),
.A2(n_439),
.B(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_418),
.A2(n_372),
.B1(n_345),
.B2(n_356),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_432),
.A2(n_452),
.B1(n_394),
.B2(n_420),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_348),
.C(n_356),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_402),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_440),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_421),
.A2(n_376),
.B(n_375),
.Y(n_435)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_436),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_397),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_403),
.A2(n_350),
.B(n_347),
.C(n_341),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_420),
.A2(n_400),
.B(n_395),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_414),
.B(n_382),
.Y(n_441)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_441),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_442),
.A2(n_444),
.B1(n_448),
.B2(n_450),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_385),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_443),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_418),
.A2(n_370),
.B1(n_365),
.B2(n_353),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_411),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_445),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_447),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_412),
.A2(n_340),
.B1(n_362),
.B2(n_364),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_412),
.A2(n_317),
.B1(n_359),
.B2(n_290),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_421),
.A2(n_335),
.B(n_318),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_454),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_386),
.A2(n_290),
.B1(n_336),
.B2(n_334),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_388),
.Y(n_453)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_453),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_337),
.B(n_336),
.Y(n_454)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_455),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_330),
.Y(n_457)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_405),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_407),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_462),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_425),
.B(n_404),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_425),
.B(n_410),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_464),
.B(n_466),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_430),
.B(n_386),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_442),
.A2(n_403),
.B1(n_408),
.B2(n_401),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_472),
.A2(n_486),
.B1(n_429),
.B2(n_454),
.Y(n_497)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_441),
.Y(n_475)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_475),
.Y(n_498)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_478),
.A2(n_456),
.B1(n_431),
.B2(n_448),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_415),
.C(n_409),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_479),
.B(n_482),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_432),
.A2(n_423),
.B1(n_389),
.B2(n_388),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_480),
.A2(n_456),
.B1(n_434),
.B2(n_435),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_427),
.B(n_387),
.C(n_413),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_426),
.B(n_387),
.C(n_413),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_485),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_426),
.A2(n_389),
.B1(n_395),
.B2(n_419),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_458),
.A2(n_396),
.B1(n_419),
.B2(n_416),
.Y(n_487)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_487),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_439),
.B(n_396),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_488),
.B(n_457),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g490 ( 
.A1(n_483),
.A2(n_449),
.B(n_424),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_490),
.A2(n_496),
.B(n_506),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_491),
.B(n_492),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_473),
.Y(n_492)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_494),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_467),
.A2(n_440),
.B(n_449),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_499),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_473),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_486),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_500),
.B(n_504),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_460),
.B(n_446),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_501),
.B(n_513),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_471),
.Y(n_502)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_502),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_445),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_437),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_505),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_467),
.A2(n_440),
.B(n_455),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_508),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g509 ( 
.A(n_469),
.B(n_443),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_509),
.B(n_517),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_472),
.A2(n_450),
.B1(n_446),
.B2(n_452),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_436),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_514),
.Y(n_540)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_475),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_516),
.Y(n_522)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_476),
.B(n_437),
.Y(n_517)
);

AO221x1_ASAP7_75t_L g525 ( 
.A1(n_497),
.A2(n_478),
.B1(n_480),
.B2(n_463),
.C(n_479),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_525),
.B(n_526),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_468),
.C(n_462),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_468),
.C(n_464),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_528),
.B(n_530),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_501),
.B(n_466),
.Y(n_530)
);

AO221x1_ASAP7_75t_L g532 ( 
.A1(n_509),
.A2(n_465),
.B1(n_471),
.B2(n_488),
.C(n_484),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_532),
.A2(n_539),
.B1(n_498),
.B2(n_515),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_511),
.B(n_470),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_533),
.B(n_535),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_491),
.B(n_477),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_459),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_537),
.B(n_538),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_493),
.B(n_459),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_510),
.B(n_391),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_526),
.C(n_493),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_541),
.B(n_543),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_538),
.B(n_537),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_542),
.B(n_545),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_540),
.C(n_520),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_496),
.Y(n_545)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_546),
.Y(n_567)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_529),
.B(n_506),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_547),
.B(n_551),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_540),
.B(n_514),
.C(n_507),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_554),
.C(n_556),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_518),
.A2(n_504),
.B(n_499),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_550),
.B(n_558),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_536),
.A2(n_510),
.B1(n_512),
.B2(n_519),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_527),
.A2(n_502),
.B1(n_498),
.B2(n_500),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_553),
.B(n_557),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_507),
.C(n_492),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_521),
.B(n_513),
.C(n_490),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_521),
.B(n_508),
.C(n_494),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_534),
.B(n_481),
.C(n_451),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_523),
.B(n_483),
.Y(n_559)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_559),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_554),
.B(n_522),
.Y(n_560)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_560),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_531),
.Y(n_561)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_561),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_531),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_565),
.A2(n_547),
.B1(n_545),
.B2(n_542),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_SL g569 ( 
.A1(n_559),
.A2(n_534),
.B(n_524),
.Y(n_569)
);

NAND3xp33_ASAP7_75t_SL g580 ( 
.A(n_569),
.B(n_573),
.C(n_552),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_557),
.A2(n_524),
.B(n_523),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_571),
.A2(n_569),
.B(n_561),
.Y(n_585)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_549),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_572),
.B(n_575),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_516),
.Y(n_573)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_558),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_563),
.B(n_544),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_576),
.B(n_577),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_574),
.B(n_555),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_580),
.B(n_565),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_566),
.A2(n_453),
.B1(n_541),
.B2(n_447),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_582),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_563),
.B(n_392),
.C(n_447),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_570),
.B(n_392),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_584),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_573),
.B(n_416),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_585),
.B(n_587),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_568),
.A2(n_337),
.B1(n_293),
.B2(n_319),
.Y(n_587)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_589),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_576),
.B(n_567),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_592),
.B(n_596),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_581),
.B(n_571),
.C(n_562),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_594),
.Y(n_600)
);

INVx6_ASAP7_75t_L g594 ( 
.A(n_578),
.Y(n_594)
);

OAI21xp33_ASAP7_75t_L g596 ( 
.A1(n_585),
.A2(n_564),
.B(n_560),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_590),
.A2(n_586),
.B(n_588),
.Y(n_598)
);

AO21x2_ASAP7_75t_L g605 ( 
.A1(n_598),
.A2(n_601),
.B(n_603),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g601 ( 
.A1(n_597),
.A2(n_582),
.B(n_562),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_596),
.B(n_587),
.Y(n_603)
);

AOI21x1_ASAP7_75t_L g604 ( 
.A1(n_599),
.A2(n_593),
.B(n_595),
.Y(n_604)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_604),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_600),
.B(n_594),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_606),
.B(n_607),
.Y(n_609)
);

AO21x2_ASAP7_75t_L g607 ( 
.A1(n_602),
.A2(n_591),
.B(n_601),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_609),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_L g611 ( 
.A1(n_610),
.A2(n_605),
.B(n_608),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_319),
.Y(n_612)
);


endmodule