module fake_ibex_980_n_751 (n_21, n_12, n_50, n_54, n_89, n_48, n_95, n_42, n_8, n_112, n_40, n_86, n_109, n_47, n_67, n_79, n_113, n_10, n_59, n_46, n_11, n_88, n_82, n_26, n_87, n_55, n_103, n_96, n_27, n_33, n_34, n_22, n_25, n_29, n_5, n_2, n_99, n_72, n_66, n_28, n_102, n_77, n_62, n_74, n_71, n_104, n_24, n_31, n_76, n_1, n_100, n_110, n_41, n_0, n_83, n_45, n_36, n_58, n_90, n_52, n_106, n_32, n_111, n_18, n_64, n_4, n_81, n_16, n_19, n_44, n_94, n_6, n_60, n_93, n_70, n_78, n_69, n_97, n_39, n_98, n_63, n_38, n_49, n_15, n_43, n_14, n_84, n_13, n_20, n_51, n_68, n_9, n_80, n_37, n_75, n_107, n_7, n_91, n_73, n_17, n_92, n_3, n_108, n_65, n_85, n_35, n_57, n_61, n_105, n_56, n_53, n_23, n_30, n_101, n_751);

input n_21;
input n_12;
input n_50;
input n_54;
input n_89;
input n_48;
input n_95;
input n_42;
input n_8;
input n_112;
input n_40;
input n_86;
input n_109;
input n_47;
input n_67;
input n_79;
input n_113;
input n_10;
input n_59;
input n_46;
input n_11;
input n_88;
input n_82;
input n_26;
input n_87;
input n_55;
input n_103;
input n_96;
input n_27;
input n_33;
input n_34;
input n_22;
input n_25;
input n_29;
input n_5;
input n_2;
input n_99;
input n_72;
input n_66;
input n_28;
input n_102;
input n_77;
input n_62;
input n_74;
input n_71;
input n_104;
input n_24;
input n_31;
input n_76;
input n_1;
input n_100;
input n_110;
input n_41;
input n_0;
input n_83;
input n_45;
input n_36;
input n_58;
input n_90;
input n_52;
input n_106;
input n_32;
input n_111;
input n_18;
input n_64;
input n_4;
input n_81;
input n_16;
input n_19;
input n_44;
input n_94;
input n_6;
input n_60;
input n_93;
input n_70;
input n_78;
input n_69;
input n_97;
input n_39;
input n_98;
input n_63;
input n_38;
input n_49;
input n_15;
input n_43;
input n_14;
input n_84;
input n_13;
input n_20;
input n_51;
input n_68;
input n_9;
input n_80;
input n_37;
input n_75;
input n_107;
input n_7;
input n_91;
input n_73;
input n_17;
input n_92;
input n_3;
input n_108;
input n_65;
input n_85;
input n_35;
input n_57;
input n_61;
input n_105;
input n_56;
input n_53;
input n_23;
input n_30;
input n_101;

output n_751;



endmodule