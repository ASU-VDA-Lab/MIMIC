module real_jpeg_32901_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_41, n_2, n_6, n_42, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_41;
input n_2;
input n_6;
input n_42;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_17;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_31;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_30;
wire n_16;
wire n_15;

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g13 ( 
.A1(n_1),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

OAI221xp5_ASAP7_75t_L g16 ( 
.A1(n_6),
.A2(n_17),
.B1(n_18),
.B2(n_34),
.C(n_35),
.Y(n_16)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_7),
.B(n_41),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_11),
.C(n_26),
.Y(n_25)
);

OAI211xp5_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_21),
.B(n_24),
.C(n_32),
.Y(n_20)
);

AOI211xp5_ASAP7_75t_SL g33 ( 
.A1(n_9),
.A2(n_21),
.B(n_24),
.C(n_32),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B(n_33),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.C(n_31),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_42),
.Y(n_28)
);


endmodule