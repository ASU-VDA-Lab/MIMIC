module fake_jpeg_5603_n_20 (n_0, n_3, n_2, n_1, n_20);

input n_0;
input n_3;
input n_2;
input n_1;

output n_20;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_4;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g4 ( 
.A(n_0),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g5 ( 
.A(n_0),
.Y(n_5)
);

INVx8_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_3),
.B(n_2),
.Y(n_7)
);

INVx4_ASAP7_75t_SL g8 ( 
.A(n_6),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

MAJIxp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_0),
.C(n_1),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_10),
.B(n_3),
.Y(n_11)
);

AOI221xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_13),
.B1(n_5),
.B2(n_8),
.C(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_5),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_14),
.A2(n_15),
.B1(n_4),
.B2(n_1),
.Y(n_17)
);

AOI22x1_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_15),
.A2(n_6),
.B1(n_4),
.B2(n_2),
.Y(n_16)
);

AOI31xp33_ASAP7_75t_L g18 ( 
.A1(n_16),
.A2(n_17),
.A3(n_4),
.B(n_1),
.Y(n_18)
);

NAND3xp33_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_0),
.C(n_1),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_19),
.A2(n_16),
.B(n_2),
.Y(n_20)
);


endmodule