module fake_jpeg_4132_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_7),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_6),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_21),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_11),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_20),
.C(n_14),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_17),
.C(n_15),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_46),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_33),
.A2(n_11),
.B(n_22),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_44),
.C(n_45),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_18),
.B1(n_13),
.B2(n_24),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_36),
.A2(n_18),
.B1(n_20),
.B2(n_14),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_15),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_25),
.B(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_51),
.B1(n_55),
.B2(n_10),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_48),
.A2(n_40),
.B1(n_45),
.B2(n_31),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_25),
.B1(n_30),
.B2(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_38),
.B1(n_40),
.B2(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_51),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_42),
.C(n_46),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.C(n_52),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_12),
.C(n_10),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_65),
.C(n_63),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_53),
.B1(n_2),
.B2(n_3),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_70),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_68),
.C(n_0),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_69),
.A2(n_66),
.A3(n_4),
.B1(n_6),
.B2(n_2),
.C(n_3),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_66),
.B(n_3),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_71),
.Y(n_77)
);


endmodule