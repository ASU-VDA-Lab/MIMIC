module fake_jpeg_18892_n_283 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_283);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_283;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_33),
.A2(n_27),
.B1(n_22),
.B2(n_21),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_29),
.B1(n_21),
.B2(n_22),
.Y(n_61)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_17),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_25),
.B(n_8),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_44),
.B(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_30),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_33),
.B1(n_27),
.B2(n_20),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_81)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_56),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_51),
.A2(n_54),
.B1(n_58),
.B2(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_30),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_62),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_40),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_21),
.B1(n_22),
.B2(n_19),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_30),
.B1(n_19),
.B2(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_39),
.B1(n_43),
.B2(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_34),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_34),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_29),
.B1(n_31),
.B2(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_75),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_70),
.Y(n_123)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_38),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_96),
.C(n_98),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_84),
.B1(n_104),
.B2(n_58),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_85),
.B1(n_18),
.B2(n_1),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_82),
.Y(n_128)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_31),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_26),
.B1(n_35),
.B2(n_24),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_26),
.B1(n_17),
.B2(n_42),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_57),
.A2(n_26),
.B1(n_35),
.B2(n_24),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_13),
.B(n_12),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_89),
.C(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_88),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_62),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_46),
.A2(n_26),
.B(n_35),
.C(n_24),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_95),
.B(n_96),
.C(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_45),
.B(n_28),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_28),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_26),
.B(n_37),
.C(n_23),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_37),
.B(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_103),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_28),
.C(n_37),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_23),
.B1(n_18),
.B2(n_17),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_2),
.CON(n_131),
.SN(n_131)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_28),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_121),
.B1(n_122),
.B2(n_124),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_71),
.A2(n_58),
.B1(n_64),
.B2(n_23),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_70),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_81),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_72),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_80),
.A2(n_84),
.B1(n_89),
.B2(n_72),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_75),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_126),
.A2(n_68),
.B(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_90),
.B1(n_98),
.B2(n_86),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_67),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_67),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_69),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_157),
.C(n_132),
.Y(n_174)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_88),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_141),
.A2(n_142),
.B(n_144),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_102),
.B(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_106),
.B(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_149),
.B(n_150),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_105),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_108),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_159),
.Y(n_181)
);

HAxp5_ASAP7_75t_SL g154 ( 
.A(n_127),
.B(n_5),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_112),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_116),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_161),
.Y(n_172)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_118),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_97),
.B(n_92),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_123),
.A2(n_77),
.B(n_100),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_126),
.Y(n_187)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_153),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_136),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_178),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_156),
.A2(n_110),
.B1(n_130),
.B2(n_119),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_183),
.B1(n_146),
.B2(n_135),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_101),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_145),
.A2(n_114),
.B1(n_78),
.B2(n_100),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_134),
.B1(n_86),
.B2(n_163),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_179),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_146),
.B1(n_135),
.B2(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_182),
.A2(n_148),
.B1(n_147),
.B2(n_117),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_126),
.B1(n_120),
.B2(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_106),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_186),
.B(n_188),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_187),
.A2(n_141),
.B(n_150),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_137),
.B(n_133),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_114),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_124),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_192),
.B(n_194),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_145),
.B(n_162),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_160),
.B(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_168),
.B1(n_208),
.B2(n_166),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_185),
.B(n_144),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_212),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_205),
.B1(n_170),
.B2(n_183),
.Y(n_215)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_129),
.B(n_77),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_178),
.Y(n_218)
);

AOI32xp33_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_129),
.A3(n_101),
.B1(n_134),
.B2(n_86),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_209),
.A2(n_169),
.B(n_172),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_180),
.B(n_129),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_186),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_180),
.B1(n_182),
.B2(n_173),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_215),
.A2(n_211),
.B1(n_204),
.B2(n_195),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_174),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_221),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_223),
.B1(n_203),
.B2(n_209),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_168),
.B1(n_166),
.B2(n_172),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_224),
.A2(n_228),
.B1(n_201),
.B2(n_196),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_188),
.C(n_175),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_195),
.C(n_202),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_192),
.A2(n_175),
.B1(n_167),
.B2(n_165),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_232),
.A2(n_236),
.B1(n_215),
.B2(n_224),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_234),
.C(n_221),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_191),
.C(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_240),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_216),
.A2(n_204),
.B(n_200),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_244),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_243),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_242),
.Y(n_252)
);

NOR3xp33_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_179),
.C(n_207),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_206),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_211),
.B(n_167),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_165),
.A3(n_164),
.B1(n_193),
.B2(n_171),
.C1(n_76),
.C2(n_14),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_219),
.Y(n_249)
);

AOI31xp67_ASAP7_75t_SL g247 ( 
.A1(n_242),
.A2(n_229),
.A3(n_226),
.B(n_222),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_253),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_238),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_254),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_251),
.A2(n_255),
.B1(n_238),
.B2(n_237),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_164),
.B(n_213),
.Y(n_254)
);

XNOR2x1_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_213),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_217),
.C(n_171),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_243),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_261),
.Y(n_269)
);

AOI31xp33_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_252),
.A3(n_240),
.B(n_231),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_260),
.A2(n_244),
.B(n_7),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_253),
.A2(n_232),
.B1(n_249),
.B2(n_254),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_SL g271 ( 
.A1(n_263),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_264),
.A2(n_250),
.B(n_255),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_246),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_76),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_256),
.C(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_268),
.A2(n_271),
.B1(n_262),
.B2(n_263),
.Y(n_272)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_272),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_261),
.B(n_10),
.C(n_12),
.D(n_16),
.Y(n_274)
);

XOR2x2_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_10),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_9),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_12),
.C(n_273),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_276),
.B(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_281),
.Y(n_283)
);


endmodule