module fake_ibex_1060_n_1046 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_201, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_166, n_195, n_163, n_26, n_188, n_200, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_202, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_207, n_54, n_19, n_1046);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_201;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_207;
input n_54;
input n_19;

output n_1046;

wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_1031;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_510;
wire n_845;
wire n_947;
wire n_972;
wire n_981;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_698;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_708;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_306;
wire n_400;
wire n_736;
wire n_550;
wire n_732;
wire n_673;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_538;
wire n_464;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_1001;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_1038;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_648;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_589;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_839;
wire n_768;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_651;
wire n_581;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_354;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_899;
wire n_843;
wire n_1019;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_379;
wire n_320;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_268;
wire n_440;
wire n_955;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_912;
wire n_890;
wire n_874;
wire n_921;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_231;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_180),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_13),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_99),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_49),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_50),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_14),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_130),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_64),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_59),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_118),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_56),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_147),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_10),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_20),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_175),
.Y(n_236)
);

NOR2xp67_ASAP7_75t_L g237 ( 
.A(n_83),
.B(n_169),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_133),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_112),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_107),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_51),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_72),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_151),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_53),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_94),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_77),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_43),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_28),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_69),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_20),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_110),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_27),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_80),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_27),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_79),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_171),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_19),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_141),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_136),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_137),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_155),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_55),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_63),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_199),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_70),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_67),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_76),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_164),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_10),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_54),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_71),
.B(n_102),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_93),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_100),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_140),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_46),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_166),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_149),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_37),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_2),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_114),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_39),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_154),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_108),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_142),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_65),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_58),
.Y(n_293)
);

BUFx10_ASAP7_75t_L g294 ( 
.A(n_60),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_146),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_82),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_95),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_60),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_143),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_157),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_204),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_84),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_109),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_123),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_59),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_53),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_22),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_202),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_194),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_163),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_196),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_68),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_177),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_152),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_125),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_21),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_144),
.Y(n_318)
);

BUFx2_ASAP7_75t_SL g319 ( 
.A(n_78),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_191),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_173),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_33),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_135),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_18),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_62),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_85),
.B(n_51),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_150),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_178),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_170),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_113),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_87),
.B(n_26),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_201),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_91),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_121),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_124),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_29),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_81),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_195),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_56),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_207),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_73),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_167),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_61),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_132),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_126),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_229),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_293),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_254),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_345),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_324),
.B(n_0),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_260),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_342),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_298),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_345),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_345),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_0),
.Y(n_356)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_304),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_229),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_322),
.B(n_1),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_209),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_223),
.B(n_2),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_274),
.B(n_3),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_238),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_238),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_305),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_269),
.Y(n_366)
);

OAI21x1_ASAP7_75t_L g367 ( 
.A1(n_269),
.A2(n_105),
.B(n_206),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_296),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_276),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_282),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_312),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_213),
.B(n_8),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_345),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_211),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g375 ( 
.A(n_304),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g376 ( 
.A1(n_286),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g377 ( 
.A1(n_296),
.A2(n_106),
.B(n_205),
.Y(n_377)
);

AOI22x1_ASAP7_75t_SL g378 ( 
.A1(n_286),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_303),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_317),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

BUFx8_ASAP7_75t_SL g383 ( 
.A(n_210),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_279),
.B(n_15),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_214),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_243),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_254),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_215),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_243),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_254),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_224),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_242),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_16),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_313),
.B(n_17),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

BUFx12f_ASAP7_75t_L g397 ( 
.A(n_294),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_228),
.B(n_18),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_230),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_399)
);

OAI22x1_ASAP7_75t_R g400 ( 
.A1(n_210),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_247),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_232),
.B(n_234),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_314),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_294),
.B(n_25),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_310),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_254),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_315),
.B(n_26),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_222),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_256),
.Y(n_411)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_295),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_259),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_222),
.A2(n_231),
.B1(n_236),
.B2(n_226),
.Y(n_414)
);

CKINVDCx8_ASAP7_75t_R g415 ( 
.A(n_319),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_226),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_262),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_231),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_250),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_267),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_277),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_315),
.B(n_34),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_295),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_253),
.Y(n_426)
);

INVx6_ASAP7_75t_L g427 ( 
.A(n_295),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_295),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_285),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_288),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_236),
.Y(n_431)
);

INVx6_ASAP7_75t_L g432 ( 
.A(n_311),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_353),
.A2(n_248),
.B1(n_264),
.B2(n_263),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_384),
.B(n_212),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_348),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_384),
.B(n_216),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_349),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_383),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_394),
.B(n_251),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_349),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_393),
.B(n_217),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_349),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_393),
.B(n_218),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_374),
.B(n_275),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_394),
.B(n_300),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_354),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_357),
.B(n_394),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_405),
.B(n_394),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_355),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_383),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_370),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_395),
.Y(n_457)
);

INVxp33_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_370),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g460 ( 
.A(n_419),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_257),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_418),
.A2(n_306),
.B1(n_339),
.B2(n_307),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_355),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_350),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_360),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_346),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_360),
.Y(n_470)
);

INVx5_ASAP7_75t_L g471 ( 
.A(n_427),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_369),
.A2(n_248),
.B1(n_264),
.B2(n_263),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_346),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_392),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_352),
.B(n_208),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_386),
.B(n_220),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_358),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_358),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_363),
.A2(n_364),
.B1(n_368),
.B2(n_366),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_363),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_364),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_373),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_356),
.B(n_221),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_373),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_403),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_366),
.Y(n_487)
);

NAND3xp33_ASAP7_75t_L g488 ( 
.A(n_406),
.B(n_253),
.C(n_344),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_351),
.B(n_225),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

AND2x2_ASAP7_75t_SL g494 ( 
.A(n_377),
.B(n_227),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_387),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_371),
.B(n_219),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_397),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_404),
.B(n_233),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_390),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_396),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_L g502 ( 
.A1(n_365),
.A2(n_273),
.B1(n_271),
.B2(n_270),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_375),
.Y(n_503)
);

NOR2x1_ASAP7_75t_L g504 ( 
.A(n_385),
.B(n_343),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_401),
.B(n_239),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_375),
.B(n_326),
.Y(n_506)
);

AND2x6_ASAP7_75t_L g507 ( 
.A(n_401),
.B(n_240),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_402),
.A2(n_258),
.B1(n_340),
.B2(n_281),
.Y(n_508)
);

INVx2_ASAP7_75t_SL g509 ( 
.A(n_388),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_391),
.B(n_411),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_390),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_SL g512 ( 
.A1(n_399),
.A2(n_329),
.B1(n_245),
.B2(n_244),
.Y(n_512)
);

BUFx6f_ASAP7_75t_SL g513 ( 
.A(n_413),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

INVx4_ASAP7_75t_SL g515 ( 
.A(n_427),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_417),
.B(n_241),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_416),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_362),
.Y(n_519)
);

NAND2xp33_ASAP7_75t_L g520 ( 
.A(n_420),
.B(n_235),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_421),
.B(n_429),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_430),
.B(n_249),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_428),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_416),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_L g527 ( 
.A(n_372),
.B(n_341),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_380),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_428),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_381),
.B(n_246),
.Y(n_531)
);

INVx3_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_410),
.B(n_331),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_428),
.Y(n_535)
);

NOR2x1p5_ASAP7_75t_L g536 ( 
.A(n_347),
.B(n_252),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_367),
.Y(n_538)
);

CKINVDCx6p67_ASAP7_75t_R g539 ( 
.A(n_347),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_432),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_431),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_359),
.B(n_255),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_412),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_377),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_412),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_412),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_425),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_425),
.Y(n_549)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_431),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_422),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_414),
.B(n_261),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_400),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_377),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_376),
.B(n_265),
.Y(n_556)
);

OR2x6_ASAP7_75t_L g557 ( 
.A(n_378),
.B(n_237),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_361),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_466),
.B(n_268),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_509),
.B(n_272),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_280),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_283),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_L g563 ( 
.A1(n_521),
.A2(n_299),
.B(n_321),
.C(n_320),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_555),
.A2(n_278),
.B(n_297),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_474),
.B(n_486),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_519),
.B(n_302),
.Y(n_566)
);

A2O1A1Ixp33_ASAP7_75t_L g567 ( 
.A1(n_521),
.A2(n_523),
.B(n_516),
.C(n_445),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_519),
.B(n_266),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_539),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_498),
.B(n_35),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_545),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_456),
.A2(n_459),
.B1(n_460),
.B2(n_458),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_434),
.B(n_35),
.Y(n_573)
);

AND2x6_ASAP7_75t_SL g574 ( 
.A(n_557),
.B(n_271),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_531),
.B(n_284),
.Y(n_577)
);

A2O1A1Ixp33_ASAP7_75t_L g578 ( 
.A1(n_516),
.A2(n_289),
.B(n_287),
.C(n_337),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_543),
.B(n_499),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_483),
.B(n_290),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_462),
.B(n_291),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_543),
.B(n_292),
.Y(n_582)
);

INVx8_ASAP7_75t_L g583 ( 
.A(n_513),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_513),
.B(n_301),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_465),
.A2(n_338),
.B1(n_335),
.B2(n_327),
.Y(n_585)
);

O2A1O1Ixp33_ASAP7_75t_L g586 ( 
.A1(n_463),
.A2(n_327),
.B(n_334),
.C(n_328),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_510),
.B(n_316),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_476),
.B(n_318),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_525),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_475),
.B(n_461),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_502),
.B(n_333),
.C(n_323),
.Y(n_591)
);

O2A1O1Ixp5_ASAP7_75t_L g592 ( 
.A1(n_435),
.A2(n_330),
.B(n_311),
.C(n_122),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_532),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_461),
.B(n_330),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_532),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_468),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_449),
.B(n_36),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_472),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_473),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_484),
.B(n_40),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_503),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_558),
.B(n_66),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_477),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_478),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_480),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_554),
.B(n_41),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_435),
.B(n_75),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_525),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_484),
.B(n_42),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_530),
.B(n_488),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_534),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_487),
.Y(n_613)
);

BUFx24_ASAP7_75t_SL g614 ( 
.A(n_508),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_491),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_508),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_616)
);

A2O1A1Ixp33_ASAP7_75t_L g617 ( 
.A1(n_523),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_493),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_437),
.B(n_86),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_512),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_437),
.B(n_444),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_530),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_504),
.B(n_50),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_444),
.B(n_52),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_447),
.B(n_52),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_497),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_442),
.B(n_88),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_447),
.B(n_89),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_452),
.B(n_54),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_452),
.B(n_55),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_517),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_450),
.B(n_57),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_556),
.A2(n_58),
.B1(n_90),
.B2(n_92),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_467),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_501),
.Y(n_635)
);

BUFx5_ASAP7_75t_L g636 ( 
.A(n_494),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_520),
.B(n_97),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_507),
.A2(n_98),
.B1(n_101),
.B2(n_103),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_518),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_527),
.B(n_104),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_522),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_538),
.A2(n_111),
.B(n_115),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_490),
.A2(n_116),
.B(n_117),
.C(n_119),
.Y(n_643)
);

BUFx12f_ASAP7_75t_L g644 ( 
.A(n_440),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_467),
.B(n_128),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_505),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_506),
.B(n_129),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_455),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g649 ( 
.A(n_526),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_507),
.A2(n_131),
.B1(n_134),
.B2(n_138),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_538),
.B(n_139),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_470),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_540),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_479),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_533),
.A2(n_145),
.B1(n_148),
.B2(n_153),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_479),
.B(n_156),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_553),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_161),
.Y(n_658)
);

AND2x6_ASAP7_75t_SL g659 ( 
.A(n_557),
.B(n_533),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_545),
.B(n_162),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_545),
.B(n_172),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_496),
.A2(n_174),
.B1(n_179),
.B2(n_183),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_453),
.B(n_184),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_553),
.A2(n_185),
.B(n_186),
.C(n_189),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_579),
.B(n_536),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_576),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_566),
.B(n_533),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_576),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_572),
.A2(n_502),
.B1(n_557),
.B2(n_541),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_622),
.B(n_601),
.Y(n_670)
);

NOR2xp67_ASAP7_75t_L g671 ( 
.A(n_634),
.B(n_540),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_573),
.A2(n_549),
.B1(n_548),
.B2(n_547),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_597),
.B(n_515),
.Y(n_673)
);

OAI22xp5_ASAP7_75t_L g674 ( 
.A1(n_567),
.A2(n_548),
.B1(n_547),
.B2(n_546),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_559),
.B(n_542),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_583),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_568),
.B(n_544),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_590),
.B(n_471),
.Y(n_678)
);

OAI21x1_ASAP7_75t_L g679 ( 
.A1(n_651),
.A2(n_454),
.B(n_529),
.Y(n_679)
);

AOI221xp5_ASAP7_75t_L g680 ( 
.A1(n_591),
.A2(n_586),
.B1(n_598),
.B2(n_614),
.C(n_585),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_571),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_631),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_L g683 ( 
.A1(n_660),
.A2(n_464),
.B(n_524),
.Y(n_683)
);

NOR2x1_ASAP7_75t_L g684 ( 
.A(n_570),
.B(n_451),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_602),
.A2(n_651),
.B(n_661),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_654),
.A2(n_471),
.B1(n_535),
.B2(n_469),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_649),
.B(n_190),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_621),
.B(n_192),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_661),
.A2(n_448),
.B(n_514),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_583),
.Y(n_690)
);

OAI21xp5_ASAP7_75t_L g691 ( 
.A1(n_592),
.A2(n_656),
.B(n_563),
.Y(n_691)
);

A2O1A1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_619),
.A2(n_511),
.B(n_443),
.C(n_439),
.Y(n_692)
);

A2O1A1Ixp33_ASAP7_75t_L g693 ( 
.A1(n_628),
.A2(n_441),
.B(n_495),
.C(n_492),
.Y(n_693)
);

OAI21xp33_ASAP7_75t_L g694 ( 
.A1(n_582),
.A2(n_560),
.B(n_587),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g695 ( 
.A1(n_656),
.A2(n_438),
.B(n_485),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_583),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_596),
.A2(n_436),
.B(n_433),
.C(n_500),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_642),
.A2(n_436),
.B(n_433),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_594),
.A2(n_446),
.B(n_482),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g700 ( 
.A1(n_607),
.A2(n_446),
.B(n_482),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_561),
.A2(n_562),
.B(n_588),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_L g703 ( 
.A1(n_607),
.A2(n_489),
.B(n_500),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_606),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_644),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_606),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_600),
.A2(n_609),
.B1(n_625),
.B2(n_624),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_646),
.A2(n_577),
.B(n_581),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_599),
.B(n_603),
.Y(n_709)
);

OR2x6_ASAP7_75t_SL g710 ( 
.A(n_569),
.B(n_648),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_604),
.B(n_605),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_612),
.B(n_613),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_SL g713 ( 
.A(n_636),
.B(n_657),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_645),
.B(n_580),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_615),
.B(n_618),
.Y(n_715)
);

BUFx2_ASAP7_75t_L g716 ( 
.A(n_574),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_626),
.A2(n_641),
.B(n_639),
.C(n_635),
.Y(n_717)
);

BUFx12f_ASAP7_75t_L g718 ( 
.A(n_659),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_632),
.B(n_633),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_663),
.A2(n_610),
.B(n_630),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_589),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_578),
.B(n_608),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_663),
.A2(n_629),
.B(n_640),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_647),
.Y(n_724)
);

O2A1O1Ixp33_ASAP7_75t_L g725 ( 
.A1(n_617),
.A2(n_616),
.B(n_620),
.C(n_623),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_616),
.Y(n_726)
);

CKINVDCx16_ASAP7_75t_R g727 ( 
.A(n_658),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_643),
.A2(n_664),
.B(n_627),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_593),
.Y(n_729)
);

NOR3xp33_ASAP7_75t_L g730 ( 
.A(n_657),
.B(n_653),
.C(n_637),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_611),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_595),
.Y(n_732)
);

CKINVDCx10_ASAP7_75t_R g733 ( 
.A(n_655),
.Y(n_733)
);

CKINVDCx10_ASAP7_75t_R g734 ( 
.A(n_662),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_638),
.B(n_650),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_565),
.B(n_434),
.C(n_502),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_565),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_579),
.B(n_537),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_579),
.B(n_537),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_564),
.A2(n_555),
.B(n_602),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_579),
.B(n_537),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_575),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_565),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_621),
.A2(n_567),
.B(n_579),
.C(n_564),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_652),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_652),
.B(n_622),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_583),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_679),
.A2(n_700),
.B(n_683),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_742),
.B(n_732),
.Y(n_749)
);

A2O1A1Ixp33_ASAP7_75t_L g750 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_750)
);

OAI21x1_ASAP7_75t_L g751 ( 
.A1(n_698),
.A2(n_695),
.B(n_699),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_737),
.B(n_687),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_698),
.A2(n_695),
.B(n_689),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_676),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_730),
.B(n_680),
.C(n_691),
.Y(n_755)
);

BUFx2_ASAP7_75t_SL g756 ( 
.A(n_676),
.Y(n_756)
);

AOI211x1_ASAP7_75t_L g757 ( 
.A1(n_672),
.A2(n_667),
.B(n_665),
.C(n_712),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_737),
.B(n_743),
.Y(n_758)
);

AO21x1_ASAP7_75t_L g759 ( 
.A1(n_713),
.A2(n_691),
.B(n_719),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_710),
.Y(n_760)
);

AOI221x1_ASAP7_75t_L g761 ( 
.A1(n_728),
.A2(n_720),
.B1(n_707),
.B2(n_703),
.C(n_722),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_707),
.A2(n_726),
.B(n_708),
.C(n_717),
.Y(n_763)
);

AO31x2_ASAP7_75t_L g764 ( 
.A1(n_674),
.A2(n_686),
.A3(n_692),
.B(n_693),
.Y(n_764)
);

AO31x2_ASAP7_75t_L g765 ( 
.A1(n_674),
.A2(n_686),
.A3(n_697),
.B(n_688),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_736),
.B(n_669),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_696),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_706),
.B(n_704),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_715),
.A2(n_724),
.B1(n_675),
.B2(n_727),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_701),
.B(n_670),
.Y(n_770)
);

BUFx4_ASAP7_75t_SL g771 ( 
.A(n_705),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_696),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_745),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_732),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_746),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_690),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_733),
.A2(n_734),
.B1(n_666),
.B2(n_668),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_718),
.A2(n_716),
.B1(n_684),
.B2(n_677),
.Y(n_778)
);

AO31x2_ASAP7_75t_L g779 ( 
.A1(n_678),
.A2(n_721),
.A3(n_731),
.B(n_729),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_671),
.B(n_673),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_744),
.A2(n_707),
.A3(n_685),
.B(n_740),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_747),
.Y(n_782)
);

A2O1A1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_783)
);

AOI22xp5_ASAP7_75t_L g784 ( 
.A1(n_737),
.A2(n_565),
.B1(n_434),
.B2(n_414),
.Y(n_784)
);

OAI21x1_ASAP7_75t_SL g785 ( 
.A1(n_702),
.A2(n_711),
.B(n_709),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_738),
.B(n_739),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_700),
.A2(n_685),
.B(n_735),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_726),
.A2(n_739),
.B1(n_741),
.B2(n_738),
.Y(n_788)
);

A2O1A1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_738),
.B(n_739),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_738),
.B(n_739),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_682),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_738),
.B(n_739),
.Y(n_793)
);

AOI21xp33_ASAP7_75t_L g794 ( 
.A1(n_665),
.A2(n_526),
.B(n_517),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_738),
.B(n_739),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_744),
.A2(n_707),
.A3(n_685),
.B(n_740),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_738),
.B(n_739),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_738),
.B(n_739),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_726),
.A2(n_434),
.B1(n_598),
.B2(n_573),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_738),
.B(n_739),
.Y(n_801)
);

INVx4_ASAP7_75t_L g802 ( 
.A(n_676),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_738),
.Y(n_803)
);

OAI21x1_ASAP7_75t_SL g804 ( 
.A1(n_702),
.A2(n_711),
.B(n_709),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_726),
.A2(n_739),
.B1(n_741),
.B2(n_738),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_737),
.A2(n_565),
.B1(n_434),
.B2(n_414),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_705),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_738),
.B(n_739),
.Y(n_809)
);

O2A1O1Ixp5_ASAP7_75t_L g810 ( 
.A1(n_719),
.A2(n_735),
.B(n_728),
.C(n_714),
.Y(n_810)
);

AO31x2_ASAP7_75t_L g811 ( 
.A1(n_744),
.A2(n_707),
.A3(n_685),
.B(n_740),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_738),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_737),
.B(n_565),
.Y(n_813)
);

BUFx4f_ASAP7_75t_SL g814 ( 
.A(n_705),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_726),
.A2(n_739),
.B1(n_741),
.B2(n_738),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_745),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_738),
.B(n_739),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_738),
.B(n_739),
.Y(n_818)
);

AOI211x1_ASAP7_75t_L g819 ( 
.A1(n_672),
.A2(n_598),
.B(n_614),
.C(n_667),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_738),
.B(n_739),
.Y(n_820)
);

AO31x2_ASAP7_75t_L g821 ( 
.A1(n_744),
.A2(n_707),
.A3(n_685),
.B(n_740),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_681),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_738),
.Y(n_823)
);

OR2x6_ASAP7_75t_L g824 ( 
.A(n_676),
.B(n_696),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_738),
.B(n_739),
.Y(n_826)
);

AO31x2_ASAP7_75t_L g827 ( 
.A1(n_744),
.A2(n_707),
.A3(n_685),
.B(n_740),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_726),
.A2(n_739),
.B1(n_741),
.B2(n_738),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_738),
.B(n_739),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_737),
.B(n_550),
.Y(n_830)
);

AOI221x1_ASAP7_75t_L g831 ( 
.A1(n_730),
.A2(n_691),
.B1(n_728),
.B2(n_723),
.C(n_695),
.Y(n_831)
);

CKINVDCx11_ASAP7_75t_R g832 ( 
.A(n_710),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_737),
.A2(n_565),
.B1(n_434),
.B2(n_414),
.Y(n_833)
);

BUFx8_ASAP7_75t_L g834 ( 
.A(n_705),
.Y(n_834)
);

AOI221x1_ASAP7_75t_L g835 ( 
.A1(n_730),
.A2(n_691),
.B1(n_728),
.B2(n_723),
.C(n_695),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_738),
.B(n_739),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_738),
.B(n_739),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_738),
.B(n_739),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_702),
.A2(n_725),
.B(n_694),
.C(n_744),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_738),
.B(n_739),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_754),
.Y(n_841)
);

OA21x2_ASAP7_75t_L g842 ( 
.A1(n_831),
.A2(n_835),
.B(n_748),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_803),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_755),
.A2(n_810),
.B(n_783),
.Y(n_844)
);

NAND2x1p5_ASAP7_75t_L g845 ( 
.A(n_754),
.B(n_767),
.Y(n_845)
);

BUFx2_ASAP7_75t_L g846 ( 
.A(n_762),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_792),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_786),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_767),
.B(n_802),
.Y(n_849)
);

OA21x2_ASAP7_75t_L g850 ( 
.A1(n_751),
.A2(n_761),
.B(n_753),
.Y(n_850)
);

BUFx2_ASAP7_75t_L g851 ( 
.A(n_836),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_812),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_785),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_802),
.B(n_782),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_790),
.B(n_791),
.Y(n_855)
);

AO31x2_ASAP7_75t_L g856 ( 
.A1(n_750),
.A2(n_799),
.A3(n_789),
.B(n_839),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_806),
.A2(n_825),
.B(n_804),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_824),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_763),
.A2(n_805),
.B(n_788),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_781),
.Y(n_860)
);

OAI21x1_ASAP7_75t_SL g861 ( 
.A1(n_815),
.A2(n_828),
.B(n_829),
.Y(n_861)
);

BUFx8_ASAP7_75t_L g862 ( 
.A(n_772),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_795),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_771),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_756),
.B(n_824),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_L g866 ( 
.A1(n_766),
.A2(n_752),
.B(n_800),
.Y(n_866)
);

OAI22xp33_ASAP7_75t_L g867 ( 
.A1(n_797),
.A2(n_840),
.B1(n_838),
.B2(n_837),
.Y(n_867)
);

OAI21x1_ASAP7_75t_SL g868 ( 
.A1(n_798),
.A2(n_801),
.B(n_826),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_758),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_809),
.A2(n_817),
.B(n_818),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_813),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_793),
.B(n_820),
.Y(n_872)
);

OAI21x1_ASAP7_75t_L g873 ( 
.A1(n_780),
.A2(n_827),
.B(n_796),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_768),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_757),
.Y(n_875)
);

NAND3xp33_ASAP7_75t_L g876 ( 
.A(n_819),
.B(n_769),
.C(n_830),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_834),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_784),
.B(n_807),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_814),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_816),
.Y(n_880)
);

OA21x2_ASAP7_75t_L g881 ( 
.A1(n_765),
.A2(n_827),
.B(n_811),
.Y(n_881)
);

OA21x2_ASAP7_75t_L g882 ( 
.A1(n_811),
.A2(n_821),
.B(n_764),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_834),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_833),
.A2(n_777),
.B1(n_775),
.B2(n_778),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_777),
.B(n_776),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_770),
.A2(n_794),
.B1(n_760),
.B2(n_808),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_749),
.A2(n_773),
.B(n_779),
.Y(n_887)
);

CKINVDCx6p67_ASAP7_75t_R g888 ( 
.A(n_832),
.Y(n_888)
);

CKINVDCx11_ASAP7_75t_R g889 ( 
.A(n_774),
.Y(n_889)
);

AO21x2_ASAP7_75t_L g890 ( 
.A1(n_822),
.A2(n_759),
.B(n_787),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_785),
.Y(n_891)
);

NOR2xp67_ASAP7_75t_L g892 ( 
.A(n_754),
.B(n_676),
.Y(n_892)
);

INVx11_ASAP7_75t_L g893 ( 
.A(n_834),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_786),
.B(n_836),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_771),
.Y(n_895)
);

NAND2x1p5_ASAP7_75t_L g896 ( 
.A(n_754),
.B(n_767),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_803),
.B(n_823),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_771),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_868),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_845),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_853),
.Y(n_901)
);

OR2x6_ASAP7_75t_L g902 ( 
.A(n_861),
.B(n_891),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_845),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_875),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_873),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_860),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_855),
.B(n_870),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_855),
.B(n_870),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_884),
.B(n_863),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_876),
.A2(n_859),
.B(n_866),
.C(n_894),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_852),
.Y(n_911)
);

AO21x2_ASAP7_75t_L g912 ( 
.A1(n_857),
.A2(n_859),
.B(n_844),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_887),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_887),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_896),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_869),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_896),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_850),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_844),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_889),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_871),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_918),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_912),
.B(n_882),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_912),
.B(n_907),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_907),
.B(n_882),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_912),
.B(n_908),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_908),
.B(n_881),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_919),
.B(n_867),
.Y(n_928)
);

OAI211xp5_ASAP7_75t_L g929 ( 
.A1(n_900),
.A2(n_866),
.B(n_849),
.C(n_878),
.Y(n_929)
);

OAI221xp5_ASAP7_75t_L g930 ( 
.A1(n_915),
.A2(n_884),
.B1(n_865),
.B2(n_851),
.C(n_897),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_905),
.B(n_890),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_901),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_909),
.B(n_856),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_902),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_915),
.A2(n_872),
.B1(n_874),
.B2(n_848),
.Y(n_935)
);

AND2x4_ASAP7_75t_SL g936 ( 
.A(n_899),
.B(n_865),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_916),
.B(n_921),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_915),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_906),
.B(n_842),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_931),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_925),
.B(n_913),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_924),
.B(n_913),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_932),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_933),
.B(n_904),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_922),
.Y(n_945)
);

INVx2_ASAP7_75t_SL g946 ( 
.A(n_936),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_933),
.B(n_910),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_924),
.B(n_914),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_938),
.B(n_915),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_928),
.B(n_911),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_932),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_924),
.B(n_926),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_934),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_925),
.B(n_914),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_945),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_943),
.Y(n_956)
);

NAND3xp33_ASAP7_75t_L g957 ( 
.A(n_947),
.B(n_930),
.C(n_929),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_952),
.B(n_926),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_940),
.B(n_926),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_943),
.Y(n_960)
);

NOR2x1_ASAP7_75t_L g961 ( 
.A(n_949),
.B(n_929),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_940),
.B(n_927),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_952),
.B(n_927),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_946),
.Y(n_964)
);

NAND2xp67_ASAP7_75t_SL g965 ( 
.A(n_942),
.B(n_939),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_952),
.B(n_927),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_951),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_951),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_950),
.B(n_937),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_952),
.B(n_923),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_950),
.B(n_937),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_956),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_969),
.B(n_947),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_955),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_956),
.Y(n_975)
);

OAI31xp33_ASAP7_75t_L g976 ( 
.A1(n_957),
.A2(n_930),
.A3(n_885),
.B(n_936),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_958),
.B(n_942),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_971),
.B(n_941),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_960),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_963),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_959),
.B(n_940),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_958),
.B(n_941),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_960),
.Y(n_983)
);

AOI21xp33_ASAP7_75t_SL g984 ( 
.A1(n_965),
.A2(n_898),
.B(n_864),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_961),
.B(n_946),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_963),
.B(n_948),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_967),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_967),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_966),
.B(n_954),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_989),
.Y(n_990)
);

AOI21xp33_ASAP7_75t_SL g991 ( 
.A1(n_976),
.A2(n_895),
.B(n_946),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_973),
.A2(n_970),
.B(n_966),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_986),
.B(n_970),
.Y(n_993)
);

AOI22xp5_ASAP7_75t_L g994 ( 
.A1(n_985),
.A2(n_959),
.B1(n_962),
.B2(n_961),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_972),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_974),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_986),
.B(n_959),
.Y(n_997)
);

OAI22xp33_ASAP7_75t_L g998 ( 
.A1(n_980),
.A2(n_964),
.B1(n_954),
.B2(n_953),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_977),
.B(n_978),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_974),
.Y(n_1000)
);

OAI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_989),
.A2(n_953),
.B1(n_928),
.B2(n_937),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_972),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_978),
.A2(n_959),
.B1(n_962),
.B2(n_948),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_981),
.B(n_962),
.Y(n_1004)
);

NAND4xp25_ASAP7_75t_SL g1005 ( 
.A(n_991),
.B(n_984),
.C(n_982),
.D(n_977),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_994),
.B(n_981),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_992),
.A2(n_981),
.B1(n_962),
.B2(n_982),
.Y(n_1007)
);

AOI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_998),
.A2(n_883),
.B(n_877),
.C(n_920),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_1003),
.A2(n_979),
.B(n_975),
.Y(n_1009)
);

OAI32xp33_ASAP7_75t_L g1010 ( 
.A1(n_990),
.A2(n_965),
.A3(n_920),
.B1(n_900),
.B2(n_903),
.Y(n_1010)
);

AOI221xp5_ASAP7_75t_L g1011 ( 
.A1(n_998),
.A2(n_988),
.B1(n_987),
.B2(n_983),
.C(n_975),
.Y(n_1011)
);

AOI31xp33_ASAP7_75t_L g1012 ( 
.A1(n_1001),
.A2(n_893),
.A3(n_888),
.B(n_935),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_SL g1013 ( 
.A1(n_1012),
.A2(n_1001),
.B(n_1004),
.Y(n_1013)
);

AOI221xp5_ASAP7_75t_L g1014 ( 
.A1(n_1005),
.A2(n_1002),
.B1(n_995),
.B2(n_999),
.C(n_996),
.Y(n_1014)
);

OAI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_1009),
.A2(n_1006),
.B(n_1007),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_1008),
.A2(n_865),
.B(n_843),
.C(n_920),
.Y(n_1016)
);

AOI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_996),
.B1(n_1000),
.B2(n_1004),
.C(n_979),
.Y(n_1017)
);

OAI21xp33_ASAP7_75t_L g1018 ( 
.A1(n_1010),
.A2(n_997),
.B(n_993),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1011),
.B(n_1000),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_1005),
.B(n_880),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_1016),
.A2(n_854),
.B(n_879),
.Y(n_1021)
);

AOI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_1015),
.A2(n_944),
.B1(n_846),
.B2(n_847),
.C(n_968),
.Y(n_1022)
);

AOI211xp5_ASAP7_75t_L g1023 ( 
.A1(n_1013),
.A2(n_892),
.B(n_886),
.C(n_928),
.Y(n_1023)
);

NAND3xp33_ASAP7_75t_SL g1024 ( 
.A(n_1014),
.B(n_1017),
.C(n_1020),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_SL g1025 ( 
.A(n_1018),
.B(n_858),
.C(n_879),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_L g1026 ( 
.A(n_1019),
.B(n_858),
.C(n_841),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1026),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_1025),
.B(n_841),
.Y(n_1028)
);

AOI211xp5_ASAP7_75t_L g1029 ( 
.A1(n_1024),
.A2(n_1023),
.B(n_1022),
.C(n_1021),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_1025),
.Y(n_1030)
);

OR2x2_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_944),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1023),
.Y(n_1032)
);

INVxp33_ASAP7_75t_L g1033 ( 
.A(n_1028),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1032),
.B(n_936),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_968),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1027),
.Y(n_1036)
);

OAI221xp5_ASAP7_75t_L g1037 ( 
.A1(n_1029),
.A2(n_935),
.B1(n_917),
.B2(n_900),
.C(n_903),
.Y(n_1037)
);

OR2x2_ASAP7_75t_L g1038 ( 
.A(n_1036),
.B(n_1030),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_1035),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1038),
.Y(n_1040)
);

CKINVDCx14_ASAP7_75t_R g1041 ( 
.A(n_1040),
.Y(n_1041)
);

AO22x2_ASAP7_75t_L g1042 ( 
.A1(n_1041),
.A2(n_1039),
.B1(n_1033),
.B2(n_1034),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_1042),
.B(n_1037),
.C(n_862),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1043),
.B(n_1028),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1044),
.B(n_862),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_1045),
.A2(n_889),
.B1(n_917),
.B2(n_903),
.Y(n_1046)
);


endmodule