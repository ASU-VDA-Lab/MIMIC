module real_jpeg_14393_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx10_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_61),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_4),
.A2(n_53),
.B1(n_61),
.B2(n_63),
.Y(n_169)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_7),
.A2(n_48),
.B1(n_49),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_7),
.A2(n_61),
.B1(n_63),
.B2(n_68),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_8),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_8),
.A2(n_38),
.B1(n_61),
.B2(n_63),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_11),
.A2(n_34),
.B1(n_35),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_51),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_11),
.A2(n_51),
.B1(n_61),
.B2(n_63),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_13),
.A2(n_48),
.B1(n_49),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_13),
.A2(n_34),
.B1(n_35),
.B2(n_65),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_14),
.A2(n_61),
.B1(n_63),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_36),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_15),
.B(n_59),
.C(n_61),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_15),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_15),
.A2(n_91),
.B1(n_112),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_15),
.B(n_101),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_121),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_20),
.B(n_95),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.C(n_84),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_21),
.B(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_40),
.C(n_69),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_36),
.B2(n_37),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_23),
.A2(n_31),
.B(n_35),
.C(n_83),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.CON(n_23),
.SN(n_23)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_24),
.A2(n_25),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_32),
.C(n_34),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g134 ( 
.A(n_27),
.B(n_35),
.CON(n_134),
.SN(n_134)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_27),
.B(n_91),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_27),
.B(n_117),
.Y(n_177)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_29),
.A2(n_33),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND3xp33_ASAP7_75t_L g135 ( 
.A(n_35),
.B(n_46),
.C(n_49),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_37),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_54),
.B2(n_69),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_42),
.A2(n_52),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_43),
.A2(n_87),
.B1(n_101),
.B2(n_134),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_45),
.A2(n_48),
.B(n_134),
.C(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_49),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_48),
.B(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_64),
.B(n_66),
.Y(n_54)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_55),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_55),
.A2(n_117),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_55),
.A2(n_117),
.B1(n_139),
.B2(n_164),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_59),
.B1(n_61),
.B2(n_63),
.Y(n_60)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_60),
.A2(n_120),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_60),
.B(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_61),
.Y(n_63)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_63),
.B(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_70),
.A2(n_71),
.B1(n_84),
.B2(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_81),
.B2(n_82),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_74),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_115),
.B(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_74),
.A2(n_75),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_75),
.B(n_131),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_79),
.Y(n_113)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_84),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.C(n_90),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_85),
.B(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_94),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_91),
.A2(n_112),
.B1(n_167),
.B2(n_175),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_108),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_106),
.B2(n_107),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_112),
.A2(n_169),
.B(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B(n_119),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_199),
.B(n_204),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_153),
.B(n_198),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_141),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_126),
.B(n_141),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_136),
.C(n_137),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_127),
.A2(n_128),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_129),
.B(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_137),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_140),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_142),
.B(n_147),
.C(n_151),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_192),
.B(n_197),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_181),
.B(n_191),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_170),
.B(n_180),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_176),
.B(n_179),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_189),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_196),
.Y(n_197)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_203),
.Y(n_204)
);


endmodule