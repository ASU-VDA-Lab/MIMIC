module fake_aes_4094_n_17 (n_1, n_2, n_4, n_3, n_5, n_0, n_17);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
NAND2xp5_ASAP7_75t_SL g7 ( .A(n_5), .B(n_1), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_2), .B(n_0), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_2), .B(n_1), .Y(n_9) );
BUFx6f_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
AND2x2_ASAP7_75t_L g11 ( .A(n_6), .B(n_3), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
OR2x2_ASAP7_75t_SL g13 ( .A(n_12), .B(n_7), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_10), .B(n_4), .Y(n_14) );
AOI22xp33_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_10), .B1(n_11), .B2(n_13), .Y(n_15) );
INVx2_ASAP7_75t_SL g16 ( .A(n_15), .Y(n_16) );
AOI221x1_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_10), .B1(n_11), .B2(n_14), .C(n_8), .Y(n_17) );
endmodule