module real_jpeg_4444_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_11;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_1),
.A2(n_24),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_2),
.Y(n_76)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_4),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_4),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_5),
.B(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_5),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_5),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_5),
.A2(n_74),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_5),
.A2(n_122),
.B(n_125),
.C(n_129),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_5),
.B(n_45),
.C(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_5),
.A2(n_74),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_5),
.B(n_16),
.Y(n_185)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_6),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_8),
.A2(n_34),
.B1(n_37),
.B2(n_38),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_8),
.A2(n_20),
.B1(n_37),
.B2(n_84),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_8),
.A2(n_37),
.B1(n_96),
.B2(n_101),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_137),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_135),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_88),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_12),
.B(n_88),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_51),
.C(n_64),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_13),
.A2(n_14),
.B1(n_51),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_32),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_23),
.Y(n_15)
);

NOR2x1_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_16),
.B(n_33),
.Y(n_91)
);

AO22x1_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_16)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_18),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_21),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_39),
.Y(n_92)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_26),
.Y(n_142)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_27),
.Y(n_150)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_28),
.Y(n_152)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_39),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_48),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_42),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_51),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_52),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_63),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_107)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_65),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_77),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_79),
.B(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_72),
.B(n_79),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_78),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_79),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_83),
.B(n_163),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_120),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_104),
.Y(n_93)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_100),
.Y(n_103)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_130),
.B1(n_131),
.B2(n_134),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_156),
.B(n_188),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_153),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_153),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_141),
.B1(n_145),
.B2(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_171),
.B(n_187),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_158),
.B(n_160),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_179),
.Y(n_178)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_183),
.Y(n_182)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_180),
.B(n_186),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_185),
.Y(n_186)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);


endmodule