module fake_jpeg_28355_n_311 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_311);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_311;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_30),
.Y(n_44)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_32),
.Y(n_67)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_49),
.B(n_31),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_32),
.C(n_34),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_32),
.B(n_34),
.C(n_36),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_61),
.Y(n_101)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_60),
.B(n_79),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_19),
.B1(n_29),
.B2(n_25),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_63),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_71),
.Y(n_103)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_70),
.C(n_67),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_67),
.B(n_75),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g70 ( 
.A1(n_44),
.A2(n_38),
.B1(n_36),
.B2(n_40),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_40),
.B1(n_47),
.B2(n_42),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_36),
.B1(n_40),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_55),
.B1(n_52),
.B2(n_61),
.Y(n_90)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_73),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_36),
.B1(n_40),
.B2(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_81),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_20),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_38),
.A3(n_21),
.B1(n_33),
.B2(n_35),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_26),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_85),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_84),
.A2(n_97),
.B1(n_58),
.B2(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_95),
.Y(n_114)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_93),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_58),
.B1(n_69),
.B2(n_56),
.Y(n_127)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_91),
.B(n_99),
.Y(n_116)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_76),
.A2(n_37),
.B1(n_34),
.B2(n_55),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_66),
.B(n_34),
.C(n_38),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_72),
.C(n_38),
.Y(n_121)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_0),
.B(n_1),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_110),
.B(n_94),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_48),
.B1(n_26),
.B2(n_23),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_38),
.B1(n_56),
.B2(n_57),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_113),
.B(n_118),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_76),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_115),
.B(n_119),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_86),
.B1(n_85),
.B2(n_111),
.Y(n_140)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_98),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_128),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_48),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_96),
.B(n_23),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_124),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_23),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_29),
.B1(n_73),
.B2(n_77),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_75),
.B(n_71),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_127),
.B1(n_134),
.B2(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_64),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_137),
.B(n_128),
.Y(n_144)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_63),
.B1(n_75),
.B2(n_37),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_75),
.B1(n_37),
.B2(n_57),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_104),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_136),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_45),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_163),
.B1(n_24),
.B2(n_28),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_151),
.B(n_158),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_97),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_146),
.B(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_25),
.B(n_16),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_111),
.B1(n_86),
.B2(n_89),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_152),
.A2(n_117),
.B1(n_133),
.B2(n_132),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g154 ( 
.A(n_119),
.B(n_20),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_157),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_88),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_114),
.A2(n_92),
.B(n_19),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_89),
.B1(n_93),
.B2(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_166),
.B1(n_127),
.B2(n_112),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_105),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_168),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_114),
.A2(n_92),
.B(n_19),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_164),
.B(n_165),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_29),
.B1(n_25),
.B2(n_16),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_24),
.B(n_28),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_121),
.A2(n_16),
.B(n_27),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_83),
.B1(n_109),
.B2(n_37),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_27),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_167),
.A2(n_22),
.B(n_17),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g168 ( 
.A1(n_126),
.A2(n_20),
.A3(n_21),
.B1(n_27),
.B2(n_22),
.C1(n_35),
.C2(n_33),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_126),
.B(n_9),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_17),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_170),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_171),
.A2(n_178),
.B1(n_179),
.B2(n_198),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_161),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_177),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_199),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_135),
.B1(n_138),
.B2(n_109),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_37),
.B1(n_52),
.B2(n_21),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_161),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_52),
.B1(n_24),
.B2(n_28),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_35),
.C(n_33),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_185),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_182),
.B(n_183),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_35),
.C(n_31),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_18),
.Y(n_186)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_18),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_156),
.B(n_35),
.C(n_18),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_197),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_192),
.B(n_15),
.Y(n_226)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_18),
.C(n_17),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_166),
.A2(n_22),
.B1(n_17),
.B2(n_15),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_150),
.B1(n_142),
.B2(n_143),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_153),
.B(n_9),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_15),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_144),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_215),
.B1(n_217),
.B2(n_220),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_154),
.C(n_162),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_196),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_158),
.B(n_184),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_195),
.B(n_198),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_214),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_139),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_171),
.A2(n_142),
.B1(n_143),
.B2(n_165),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_139),
.B1(n_151),
.B2(n_169),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_200),
.A2(n_163),
.B1(n_167),
.B2(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_174),
.A2(n_15),
.B1(n_8),
.B2(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_2),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_189),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_7),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_191),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_203),
.B(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_173),
.B1(n_190),
.B2(n_199),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_228),
.A2(n_207),
.B1(n_204),
.B2(n_216),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_236),
.Y(n_255)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_235),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_223),
.A2(n_189),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_240),
.Y(n_247)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_184),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_239),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_181),
.C(n_180),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_202),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_197),
.C(n_185),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_195),
.C(n_8),
.Y(n_242)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_253),
.B1(n_12),
.B2(n_3),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_214),
.C(n_210),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_261),
.C(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_227),
.B(n_219),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_11),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_228),
.A2(n_207),
.B1(n_218),
.B2(n_211),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_243),
.A2(n_206),
.B(n_219),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_14),
.B(n_12),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_230),
.A2(n_226),
.B1(n_3),
.B2(n_4),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_7),
.C(n_13),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_262),
.B(n_273),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_239),
.C(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_275),
.C(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_269),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_236),
.B(n_242),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_265),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_229),
.B(n_233),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_267),
.B(n_272),
.Y(n_277)
);

AOI21x1_ASAP7_75t_SL g267 ( 
.A1(n_246),
.A2(n_2),
.B(n_3),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_7),
.B(n_13),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_268),
.B(n_2),
.Y(n_283)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_257),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

INVx11_ASAP7_75t_L g278 ( 
.A(n_271),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_4),
.B(n_5),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_274),
.A2(n_259),
.B1(n_253),
.B2(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_250),
.C(n_256),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_280),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_277),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_256),
.B1(n_255),
.B2(n_5),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_269),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_275),
.C(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_262),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_290),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_280),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_295),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_278),
.B(n_281),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_285),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_268),
.Y(n_295)
);

AOI21x1_ASAP7_75t_L g299 ( 
.A1(n_295),
.A2(n_278),
.B(n_267),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_294),
.B(n_288),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_285),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_298),
.A2(n_293),
.B(n_291),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_302),
.A2(n_296),
.B(n_297),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_304),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_306),
.A2(n_303),
.B(n_284),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_307),
.A2(n_305),
.B(n_5),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_4),
.C(n_6),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_309),
.B(n_6),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_6),
.Y(n_311)
);


endmodule