module real_aes_7545_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_140;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g109 ( .A(n_0), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g457 ( .A1(n_1), .A2(n_147), .B(n_159), .C(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g266 ( .A(n_2), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_3), .A2(n_174), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_4), .B(n_170), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g173 ( .A1(n_5), .A2(n_174), .B(n_175), .Y(n_173) );
AND2x6_ASAP7_75t_L g147 ( .A(n_6), .B(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_7), .A2(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g106 ( .A(n_8), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_8), .B(n_40), .Y(n_127) );
INVx1_ASAP7_75t_L g473 ( .A(n_9), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_10), .B(n_180), .Y(n_461) );
INVx1_ASAP7_75t_L g182 ( .A(n_11), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_12), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
INVx1_ASAP7_75t_L g248 ( .A(n_14), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_15), .A2(n_183), .B(n_249), .C(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_16), .B(n_170), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_17), .B(n_193), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_18), .B(n_174), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_19), .B(n_515), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_20), .A2(n_150), .B(n_234), .C(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_21), .B(n_170), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_22), .B(n_180), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_23), .A2(n_246), .B(n_247), .C(n_249), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_24), .B(n_180), .Y(n_523) );
CKINVDCx16_ASAP7_75t_R g532 ( .A(n_25), .Y(n_532) );
INVx1_ASAP7_75t_L g522 ( .A(n_26), .Y(n_522) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_27), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_28), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_29), .B(n_180), .Y(n_267) );
INVx1_ASAP7_75t_L g511 ( .A(n_30), .Y(n_511) );
INVx1_ASAP7_75t_L g158 ( .A(n_31), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_32), .A2(n_100), .B1(n_114), .B2(n_729), .Y(n_99) );
INVx2_ASAP7_75t_L g152 ( .A(n_33), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_34), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_35), .A2(n_184), .B(n_234), .C(n_500), .Y(n_499) );
INVxp67_ASAP7_75t_L g512 ( .A(n_36), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g203 ( .A1(n_37), .A2(n_147), .B(n_159), .C(n_204), .Y(n_203) );
CKINVDCx14_ASAP7_75t_R g498 ( .A(n_38), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_39), .A2(n_159), .B(n_521), .C(n_525), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_40), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g156 ( .A(n_41), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_42), .A2(n_179), .B(n_209), .C(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_43), .B(n_180), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_44), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_45), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_46), .Y(n_128) );
INVx1_ASAP7_75t_L g488 ( .A(n_47), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g162 ( .A(n_48), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_49), .B(n_174), .Y(n_236) );
AOI222xp33_ASAP7_75t_SL g129 ( .A1(n_50), .A2(n_59), .B1(n_130), .B2(n_715), .C1(n_716), .C2(n_720), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_51), .A2(n_150), .B1(n_153), .B2(n_159), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_52), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_53), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g178 ( .A1(n_54), .A2(n_179), .B(n_181), .C(n_184), .Y(n_178) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_55), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_56), .Y(n_223) );
INVx1_ASAP7_75t_L g176 ( .A(n_57), .Y(n_176) );
INVx1_ASAP7_75t_L g148 ( .A(n_58), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_59), .Y(n_715) );
INVx1_ASAP7_75t_L g143 ( .A(n_60), .Y(n_143) );
INVx1_ASAP7_75t_SL g501 ( .A(n_61), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_62), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_63), .B(n_170), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_64), .A2(n_447), .B1(n_717), .B2(n_726), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_64), .Y(n_726) );
INVx1_ASAP7_75t_L g535 ( .A(n_65), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_SL g192 ( .A1(n_66), .A2(n_184), .B(n_193), .C(n_194), .Y(n_192) );
INVxp67_ASAP7_75t_L g195 ( .A(n_67), .Y(n_195) );
INVx1_ASAP7_75t_L g113 ( .A(n_68), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_69), .A2(n_174), .B(n_469), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_70), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_71), .Y(n_167) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_72), .A2(n_174), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g216 ( .A(n_73), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_74), .A2(n_242), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g480 ( .A(n_75), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g519 ( .A(n_76), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_L g217 ( .A1(n_77), .A2(n_147), .B(n_159), .C(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_78), .A2(n_174), .B(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g483 ( .A(n_79), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_80), .B(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx1_ASAP7_75t_L g459 ( .A(n_82), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_83), .B(n_193), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_84), .A2(n_147), .B(n_159), .C(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g110 ( .A(n_85), .Y(n_110) );
OR2x2_ASAP7_75t_L g124 ( .A(n_85), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g714 ( .A(n_85), .B(n_126), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_86), .A2(n_159), .B(n_534), .C(n_537), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_87), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g270 ( .A(n_88), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_89), .A2(n_147), .B(n_159), .C(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_90), .Y(n_238) );
INVx1_ASAP7_75t_L g191 ( .A(n_91), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g244 ( .A(n_92), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_93), .B(n_206), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_94), .B(n_172), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_95), .B(n_172), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_96), .B(n_113), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_97), .A2(n_174), .B(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g491 ( .A(n_98), .Y(n_491) );
BUFx4f_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
INVx3_ASAP7_75t_SL g729 ( .A(n_103), .Y(n_729) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_109), .B(n_110), .C(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g126 ( .A(n_109), .B(n_127), .Y(n_126) );
OR2x2_ASAP7_75t_L g446 ( .A(n_110), .B(n_126), .Y(n_446) );
NOR2x2_ASAP7_75t_L g722 ( .A(n_110), .B(n_125), .Y(n_722) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_129), .B1(n_723), .B2(n_724), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g723 ( .A(n_118), .Y(n_723) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_121), .A2(n_725), .B(n_727), .Y(n_724) );
NOR2xp33_ASAP7_75t_SL g121 ( .A(n_122), .B(n_128), .Y(n_121) );
INVx1_ASAP7_75t_SL g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g728 ( .A(n_124), .Y(n_728) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_444), .B1(n_447), .B2(n_714), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_SL g716 ( .A1(n_132), .A2(n_444), .B1(n_717), .B2(n_718), .Y(n_716) );
AND3x1_ASAP7_75t_L g132 ( .A(n_133), .B(n_369), .C(n_418), .Y(n_132) );
NOR3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_276), .C(n_314), .Y(n_133) );
OAI222xp33_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_197), .B1(n_251), .B2(n_257), .C1(n_271), .C2(n_274), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_168), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_136), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_136), .B(n_319), .Y(n_410) );
BUFx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g287 ( .A(n_137), .B(n_188), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_137), .B(n_169), .Y(n_295) );
AND2x2_ASAP7_75t_L g330 ( .A(n_137), .B(n_307), .Y(n_330) );
OR2x2_ASAP7_75t_L g354 ( .A(n_137), .B(n_169), .Y(n_354) );
OR2x2_ASAP7_75t_L g362 ( .A(n_137), .B(n_261), .Y(n_362) );
AND2x2_ASAP7_75t_L g365 ( .A(n_137), .B(n_188), .Y(n_365) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
OR2x2_ASAP7_75t_L g259 ( .A(n_138), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g273 ( .A(n_138), .B(n_188), .Y(n_273) );
AND2x2_ASAP7_75t_L g323 ( .A(n_138), .B(n_261), .Y(n_323) );
AND2x2_ASAP7_75t_L g336 ( .A(n_138), .B(n_169), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_138), .B(n_422), .Y(n_443) );
AO21x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_145), .B(n_166), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_139), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_139), .A2(n_262), .B(n_269), .Y(n_261) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_SL g187 ( .A(n_141), .B(n_142), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_149), .B1(n_162), .B2(n_163), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g175 ( .A1(n_146), .A2(n_176), .B(n_177), .C(n_178), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_146), .A2(n_177), .B(n_191), .C(n_192), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_146), .A2(n_177), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g469 ( .A1(n_146), .A2(n_177), .B(n_470), .C(n_471), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g479 ( .A1(n_146), .A2(n_177), .B(n_480), .C(n_481), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_SL g487 ( .A1(n_146), .A2(n_177), .B(n_488), .C(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_146), .A2(n_177), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_146), .A2(n_177), .B(n_508), .C(n_509), .Y(n_507) );
INVx1_ASAP7_75t_L g537 ( .A(n_146), .Y(n_537) );
INVx4_ASAP7_75t_SL g146 ( .A(n_147), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g163 ( .A(n_147), .B(n_164), .Y(n_163) );
AND2x4_ASAP7_75t_L g174 ( .A(n_147), .B(n_164), .Y(n_174) );
BUFx3_ASAP7_75t_L g525 ( .A(n_147), .Y(n_525) );
INVx2_ASAP7_75t_L g268 ( .A(n_150), .Y(n_268) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g160 ( .A(n_152), .Y(n_160) );
INVx1_ASAP7_75t_L g165 ( .A(n_152), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g153 ( .A1(n_154), .A2(n_156), .B1(n_157), .B2(n_158), .Y(n_153) );
INVx2_ASAP7_75t_L g157 ( .A(n_154), .Y(n_157) );
INVx4_ASAP7_75t_L g246 ( .A(n_154), .Y(n_246) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
AND2x2_ASAP7_75t_L g164 ( .A(n_155), .B(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx3_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
INVx1_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
INVx2_ASAP7_75t_L g460 ( .A(n_157), .Y(n_460) );
INVx5_ASAP7_75t_L g177 ( .A(n_159), .Y(n_177) );
AND2x6_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
BUFx3_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_163), .A2(n_216), .B(n_217), .Y(n_215) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_163), .A2(n_263), .B(n_264), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g455 ( .A1(n_163), .A2(n_456), .B(n_457), .Y(n_455) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_163), .A2(n_187), .B(n_519), .C(n_520), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_163), .A2(n_532), .B(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g513 ( .A(n_165), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g361 ( .A1(n_168), .A2(n_362), .B(n_363), .C(n_366), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_168), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_168), .B(n_306), .Y(n_428) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_188), .Y(n_168) );
AND2x2_ASAP7_75t_SL g272 ( .A(n_169), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g286 ( .A(n_169), .Y(n_286) );
AND2x2_ASAP7_75t_L g313 ( .A(n_169), .B(n_307), .Y(n_313) );
INVx1_ASAP7_75t_SL g321 ( .A(n_169), .Y(n_321) );
AND2x2_ASAP7_75t_L g344 ( .A(n_169), .B(n_345), .Y(n_344) );
BUFx2_ASAP7_75t_L g422 ( .A(n_169), .Y(n_422) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_173), .B(n_186), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_171), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_171), .B(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_171), .B(n_527), .Y(n_526) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_171), .A2(n_531), .B(n_538), .Y(n_530) );
INVx4_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_172), .A2(n_189), .B(n_196), .Y(n_188) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_172), .Y(n_477) );
BUFx2_ASAP7_75t_L g242 ( .A(n_174), .Y(n_242) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx4_ASAP7_75t_L g234 ( .A(n_180), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_183), .B(n_195), .Y(n_194) );
INVx5_ASAP7_75t_L g206 ( .A(n_183), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_183), .B(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g224 ( .A(n_187), .Y(n_224) );
INVx2_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_187), .A2(n_241), .B(n_250), .Y(n_240) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_187), .A2(n_468), .B(n_474), .Y(n_467) );
BUFx2_ASAP7_75t_L g258 ( .A(n_188), .Y(n_258) );
INVx1_ASAP7_75t_L g320 ( .A(n_188), .Y(n_320) );
INVx3_ASAP7_75t_L g345 ( .A(n_188), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_197), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_225), .Y(n_197) );
INVx1_ASAP7_75t_L g341 ( .A(n_198), .Y(n_341) );
OAI32xp33_ASAP7_75t_L g347 ( .A1(n_198), .A2(n_286), .A3(n_348), .B1(n_349), .B2(n_350), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_198), .A2(n_352), .B1(n_355), .B2(n_360), .Y(n_351) );
INVx4_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g289 ( .A(n_199), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g367 ( .A(n_199), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g437 ( .A(n_199), .B(n_383), .Y(n_437) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
AND2x2_ASAP7_75t_L g252 ( .A(n_200), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
INVx1_ASAP7_75t_L g301 ( .A(n_200), .Y(n_301) );
OR2x2_ASAP7_75t_L g309 ( .A(n_200), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g316 ( .A(n_200), .B(n_290), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_200), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g337 ( .A(n_200), .B(n_255), .Y(n_337) );
INVx3_ASAP7_75t_L g359 ( .A(n_200), .Y(n_359) );
AND2x2_ASAP7_75t_L g384 ( .A(n_200), .B(n_256), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_200), .B(n_349), .Y(n_432) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_212), .Y(n_200) );
AOI21xp5_ASAP7_75t_SL g201 ( .A1(n_202), .A2(n_203), .B(n_211), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_207), .B(n_208), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_206), .A2(n_266), .B(n_267), .C(n_268), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_206), .A2(n_246), .B1(n_511), .B2(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_206), .A2(n_522), .B(n_523), .C(n_524), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_208), .A2(n_219), .B(n_220), .Y(n_218) );
O2A1O1Ixp5_ASAP7_75t_L g458 ( .A1(n_208), .A2(n_459), .B(n_460), .C(n_461), .Y(n_458) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_208), .A2(n_460), .B(n_535), .C(n_536), .Y(n_534) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx1_ASAP7_75t_L g221 ( .A(n_211), .Y(n_221) );
INVx2_ASAP7_75t_L g256 ( .A(n_214), .Y(n_256) );
AND2x2_ASAP7_75t_L g388 ( .A(n_214), .B(n_226), .Y(n_388) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_221), .B(n_222), .Y(n_214) );
INVx1_ASAP7_75t_L g505 ( .A(n_221), .Y(n_505) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_221), .A2(n_558), .B(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_224), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_224), .B(n_270), .Y(n_269) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_224), .A2(n_455), .B(n_462), .Y(n_454) );
INVx2_ASAP7_75t_L g430 ( .A(n_225), .Y(n_430) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_239), .Y(n_225) );
INVx1_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_226), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_226), .B(n_256), .Y(n_310) );
AND2x2_ASAP7_75t_L g368 ( .A(n_226), .B(n_291), .Y(n_368) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g254 ( .A(n_227), .Y(n_254) );
AND2x2_ASAP7_75t_L g281 ( .A(n_227), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_227), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_227), .B(n_256), .Y(n_356) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_237), .Y(n_227) );
INVx1_ASAP7_75t_L g515 ( .A(n_228), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_228), .B(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_236), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_235), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_234), .B(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_239), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g303 ( .A(n_239), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_239), .B(n_256), .Y(n_349) );
AND2x2_ASAP7_75t_L g358 ( .A(n_239), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g383 ( .A(n_239), .Y(n_383) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g255 ( .A(n_240), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g291 ( .A(n_240), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_246), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_246), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_246), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g419 ( .A1(n_251), .A2(n_261), .B1(n_420), .B2(n_423), .Y(n_419) );
INVx1_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
OAI21xp5_ASAP7_75t_SL g442 ( .A1(n_253), .A2(n_364), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_254), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g401 ( .A(n_254), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_255), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g328 ( .A(n_255), .B(n_281), .Y(n_328) );
INVx2_ASAP7_75t_L g284 ( .A(n_256), .Y(n_284) );
INVx1_ASAP7_75t_L g334 ( .A(n_256), .Y(n_334) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_257), .A2(n_409), .B1(n_426), .B2(n_429), .C(n_431), .Y(n_425) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_258), .B(n_307), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_259), .B(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g350 ( .A(n_259), .B(n_296), .Y(n_350) );
INVx3_ASAP7_75t_SL g391 ( .A(n_259), .Y(n_391) );
AND2x2_ASAP7_75t_L g335 ( .A(n_260), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g364 ( .A(n_260), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_260), .B(n_273), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_260), .B(n_319), .Y(n_405) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g307 ( .A(n_261), .Y(n_307) );
OAI322xp33_ASAP7_75t_L g402 ( .A1(n_261), .A2(n_333), .A3(n_355), .B1(n_403), .B2(n_405), .C1(n_406), .C2(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI21xp33_ASAP7_75t_L g426 ( .A1(n_272), .A2(n_275), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_SL g352 ( .A(n_273), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g374 ( .A(n_273), .B(n_286), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_273), .B(n_313), .Y(n_389) );
INVxp67_ASAP7_75t_L g340 ( .A(n_275), .Y(n_340) );
AOI211xp5_ASAP7_75t_L g346 ( .A1(n_275), .A2(n_347), .B(n_351), .C(n_361), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_285), .B1(n_288), .B2(n_292), .C(n_297), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g300 ( .A(n_284), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g417 ( .A(n_284), .Y(n_417) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_285), .A2(n_434), .B1(n_439), .B2(n_440), .C(n_442), .Y(n_433) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_286), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_SL g333 ( .A(n_286), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_286), .B(n_364), .Y(n_371) );
AND2x2_ASAP7_75t_L g413 ( .A(n_286), .B(n_391), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_287), .B(n_312), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g408 ( .A1(n_287), .A2(n_299), .B1(n_409), .B2(n_410), .Y(n_408) );
OR2x2_ASAP7_75t_L g439 ( .A(n_287), .B(n_307), .Y(n_439) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g416 ( .A(n_290), .Y(n_416) );
AND2x2_ASAP7_75t_L g441 ( .A(n_290), .B(n_384), .Y(n_441) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_SL g293 ( .A(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g305 ( .A(n_295), .B(n_306), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_304), .B1(n_308), .B2(n_311), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_302), .Y(n_299) );
INVx1_ASAP7_75t_L g372 ( .A(n_300), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_300), .B(n_340), .Y(n_407) );
AOI322xp5_ASAP7_75t_L g331 ( .A1(n_302), .A2(n_332), .A3(n_334), .B1(n_335), .B2(n_337), .C1(n_338), .C2(n_342), .Y(n_331) );
INVxp67_ASAP7_75t_L g325 ( .A(n_303), .Y(n_325) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_305), .A2(n_310), .B1(n_327), .B2(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_306), .B(n_319), .Y(n_406) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_307), .B(n_345), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_307), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g403 ( .A(n_309), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NAND3xp33_ASAP7_75t_SL g314 ( .A(n_315), .B(n_331), .C(n_346), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_322), .B2(n_324), .C(n_326), .Y(n_315) );
AND2x2_ASAP7_75t_L g322 ( .A(n_318), .B(n_323), .Y(n_322) );
INVx3_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g332 ( .A(n_323), .B(n_333), .Y(n_332) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_325), .Y(n_404) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_330), .B(n_344), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_333), .B(n_391), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_334), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g409 ( .A(n_337), .Y(n_409) );
AND2x2_ASAP7_75t_L g424 ( .A(n_337), .B(n_401), .Y(n_424) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_348), .A2(n_419), .B(n_425), .C(n_433), .Y(n_418) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_388), .Y(n_387) );
NAND2x1_ASAP7_75t_SL g429 ( .A(n_359), .B(n_430), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g399 ( .A(n_362), .Y(n_399) );
INVx1_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
AND2x2_ASAP7_75t_L g398 ( .A(n_368), .B(n_384), .Y(n_398) );
NOR5xp2_ASAP7_75t_L g369 ( .A(n_370), .B(n_385), .C(n_402), .D(n_408), .E(n_411), .Y(n_369) );
OAI221xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_373), .B2(n_375), .C(n_377), .Y(n_370) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_374), .B(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_384), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g400 ( .A(n_384), .B(n_401), .Y(n_400) );
OAI221xp5_ASAP7_75t_SL g385 ( .A1(n_386), .A2(n_389), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B1(n_399), .B2(n_400), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g438 ( .A(n_398), .Y(n_438) );
AOI211xp5_ASAP7_75t_SL g411 ( .A1(n_412), .A2(n_414), .B(n_416), .C(n_417), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
CKINVDCx14_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g717 ( .A(n_447), .Y(n_717) );
OR2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_669), .Y(n_447) );
NAND5xp2_ASAP7_75t_L g448 ( .A(n_449), .B(n_581), .C(n_619), .D(n_640), .E(n_657), .Y(n_448) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_553), .C(n_574), .Y(n_449) );
OAI221xp5_ASAP7_75t_SL g450 ( .A1(n_451), .A2(n_493), .B1(n_516), .B2(n_540), .C(n_544), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_464), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_453), .B(n_542), .Y(n_561) );
OR2x2_ASAP7_75t_L g588 ( .A(n_453), .B(n_476), .Y(n_588) );
AND2x2_ASAP7_75t_L g602 ( .A(n_453), .B(n_476), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_453), .B(n_467), .Y(n_616) );
AND2x2_ASAP7_75t_L g654 ( .A(n_453), .B(n_618), .Y(n_654) );
AND2x2_ASAP7_75t_L g683 ( .A(n_453), .B(n_593), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_453), .B(n_565), .Y(n_700) );
INVx4_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g580 ( .A(n_454), .B(n_475), .Y(n_580) );
BUFx3_ASAP7_75t_L g605 ( .A(n_454), .Y(n_605) );
AND2x2_ASAP7_75t_L g634 ( .A(n_454), .B(n_476), .Y(n_634) );
AND3x2_ASAP7_75t_L g647 ( .A(n_454), .B(n_648), .C(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g570 ( .A(n_464), .Y(n_570) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_475), .Y(n_464) );
AOI32xp33_ASAP7_75t_L g625 ( .A1(n_465), .A2(n_577), .A3(n_626), .B1(n_629), .B2(n_630), .Y(n_625) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g552 ( .A(n_466), .B(n_475), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_466), .B(n_580), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_466), .B(n_602), .Y(n_630) );
OR2x2_ASAP7_75t_L g636 ( .A(n_466), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_466), .B(n_591), .Y(n_661) );
OR2x2_ASAP7_75t_L g679 ( .A(n_466), .B(n_504), .Y(n_679) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_L g543 ( .A(n_467), .B(n_485), .Y(n_543) );
INVx2_ASAP7_75t_L g565 ( .A(n_467), .Y(n_565) );
OR2x2_ASAP7_75t_L g587 ( .A(n_467), .B(n_485), .Y(n_587) );
AND2x2_ASAP7_75t_L g592 ( .A(n_467), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_467), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g648 ( .A(n_467), .B(n_542), .Y(n_648) );
INVx1_ASAP7_75t_SL g699 ( .A(n_475), .Y(n_699) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
INVx1_ASAP7_75t_SL g542 ( .A(n_476), .Y(n_542) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_476), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_476), .B(n_628), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_476), .B(n_565), .C(n_683), .Y(n_694) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_484), .Y(n_476) );
OA21x2_ASAP7_75t_L g485 ( .A1(n_477), .A2(n_486), .B(n_492), .Y(n_485) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_477), .A2(n_496), .B(n_502), .Y(n_495) );
INVx2_ASAP7_75t_L g593 ( .A(n_485), .Y(n_593) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_485), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
INVx1_ASAP7_75t_L g629 ( .A(n_494), .Y(n_629) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g547 ( .A(n_495), .B(n_529), .Y(n_547) );
INVx2_ASAP7_75t_L g564 ( .A(n_495), .Y(n_564) );
AND2x2_ASAP7_75t_L g569 ( .A(n_495), .B(n_530), .Y(n_569) );
AND2x2_ASAP7_75t_L g584 ( .A(n_495), .B(n_517), .Y(n_584) );
AND2x2_ASAP7_75t_L g596 ( .A(n_495), .B(n_568), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_503), .B(n_612), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_503), .B(n_569), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_503), .B(n_688), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_503), .B(n_563), .Y(n_691) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g528 ( .A(n_504), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_504), .B(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g573 ( .A(n_504), .B(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g599 ( .A(n_504), .B(n_529), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_504), .B(n_639), .Y(n_638) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_506), .B(n_514), .Y(n_504) );
INVx1_ASAP7_75t_L g558 ( .A(n_506), .Y(n_558) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_510), .B(n_513), .Y(n_509) );
INVx2_ASAP7_75t_L g524 ( .A(n_513), .Y(n_524) );
INVx1_ASAP7_75t_L g559 ( .A(n_514), .Y(n_559) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_528), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_517), .B(n_550), .Y(n_549) );
AND2x4_ASAP7_75t_L g563 ( .A(n_517), .B(n_564), .Y(n_563) );
INVx3_ASAP7_75t_SL g568 ( .A(n_517), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_517), .B(n_555), .Y(n_621) );
OR2x2_ASAP7_75t_L g631 ( .A(n_517), .B(n_557), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_517), .B(n_599), .Y(n_659) );
OR2x2_ASAP7_75t_L g689 ( .A(n_517), .B(n_529), .Y(n_689) );
AND2x2_ASAP7_75t_L g693 ( .A(n_517), .B(n_530), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_517), .B(n_569), .Y(n_706) );
AND2x2_ASAP7_75t_L g713 ( .A(n_517), .B(n_595), .Y(n_713) );
OR2x6_ASAP7_75t_L g517 ( .A(n_518), .B(n_526), .Y(n_517) );
INVx1_ASAP7_75t_SL g656 ( .A(n_528), .Y(n_656) );
AND2x2_ASAP7_75t_L g595 ( .A(n_529), .B(n_557), .Y(n_595) );
AND2x2_ASAP7_75t_L g609 ( .A(n_529), .B(n_564), .Y(n_609) );
AND2x2_ASAP7_75t_L g612 ( .A(n_529), .B(n_568), .Y(n_612) );
INVx1_ASAP7_75t_L g639 ( .A(n_529), .Y(n_639) );
INVx2_ASAP7_75t_SL g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g551 ( .A(n_530), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g710 ( .A1(n_541), .A2(n_587), .B(n_711), .C(n_712), .Y(n_710) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_543), .B(n_560), .Y(n_575) );
AND2x2_ASAP7_75t_L g601 ( .A(n_543), .B(n_602), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_545), .A2(n_548), .B(n_552), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_546), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g572 ( .A(n_547), .B(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_547), .B(n_568), .Y(n_613) );
AND2x2_ASAP7_75t_L g704 ( .A(n_547), .B(n_555), .Y(n_704) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g577 ( .A(n_551), .B(n_564), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_551), .B(n_562), .Y(n_578) );
OAI322xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_561), .A3(n_562), .B1(n_565), .B2(n_566), .C1(n_570), .C2(n_571), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_560), .Y(n_554) );
AND2x2_ASAP7_75t_L g665 ( .A(n_555), .B(n_577), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_555), .B(n_629), .Y(n_711) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g608 ( .A(n_557), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g674 ( .A(n_561), .B(n_587), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_562), .B(n_656), .Y(n_655) );
INVx3_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_563), .B(n_595), .Y(n_652) );
AND2x2_ASAP7_75t_L g598 ( .A(n_564), .B(n_568), .Y(n_598) );
AND2x2_ASAP7_75t_L g606 ( .A(n_565), .B(n_607), .Y(n_606) );
A2O1A1Ixp33_ASAP7_75t_L g703 ( .A1(n_565), .A2(n_644), .B(n_704), .C(n_705), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_566), .A2(n_579), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_568), .B(n_595), .Y(n_635) );
AND2x2_ASAP7_75t_L g641 ( .A(n_568), .B(n_609), .Y(n_641) );
AND2x2_ASAP7_75t_L g675 ( .A(n_568), .B(n_577), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_569), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_SL g685 ( .A(n_569), .Y(n_685) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_573), .A2(n_601), .B1(n_603), .B2(n_608), .Y(n_600) );
OAI22xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_576), .B1(n_578), .B2(n_579), .Y(n_574) );
OAI22xp33_ASAP7_75t_L g610 ( .A1(n_575), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_610) );
INVxp67_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_580), .A2(n_682), .B1(n_684), .B2(n_686), .C(n_690), .Y(n_681) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_585), .B(n_589), .C(n_610), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
OR2x2_ASAP7_75t_L g651 ( .A(n_587), .B(n_604), .Y(n_651) );
INVx1_ASAP7_75t_L g702 ( .A(n_587), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_588), .A2(n_590), .B1(n_594), .B2(n_597), .C(n_600), .Y(n_589) );
INVx2_ASAP7_75t_SL g644 ( .A(n_588), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g709 ( .A(n_591), .Y(n_709) );
AND2x2_ASAP7_75t_L g633 ( .A(n_592), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g618 ( .A(n_593), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g680 ( .A(n_596), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_604), .B(n_706), .Y(n_705) );
CKINVDCx16_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g649 ( .A(n_607), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g619 ( .A1(n_608), .A2(n_620), .B(n_622), .C(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g697 ( .A(n_611), .Y(n_697) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_615), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx2_ASAP7_75t_L g628 ( .A(n_618), .Y(n_628) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI222xp33_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_631), .B1(n_632), .B2(n_635), .C1(n_636), .C2(n_638), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g664 ( .A(n_628), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_631), .B(n_685), .Y(n_684) );
NAND2xp33_ASAP7_75t_SL g662 ( .A(n_632), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g637 ( .A(n_634), .Y(n_637) );
AND2x2_ASAP7_75t_L g701 ( .A(n_634), .B(n_702), .Y(n_701) );
OR2x2_ASAP7_75t_L g667 ( .A(n_637), .B(n_664), .Y(n_667) );
INVx1_ASAP7_75t_L g696 ( .A(n_638), .Y(n_696) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_642), .B(n_645), .C(n_650), .Y(n_640) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_644), .B(n_664), .Y(n_663) );
INVx2_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AOI322xp5_ASAP7_75t_L g695 ( .A1(n_647), .A2(n_675), .A3(n_680), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_701), .Y(n_695) );
AND2x2_ASAP7_75t_L g682 ( .A(n_648), .B(n_683), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_653), .B2(n_655), .Y(n_650) );
INVxp33_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .B1(n_662), .B2(n_665), .C(n_666), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
NAND5xp2_ASAP7_75t_L g669 ( .A(n_670), .B(n_681), .C(n_695), .D(n_703), .E(n_707), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_675), .B(n_676), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVxp33_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g707 ( .A1(n_683), .A2(n_708), .B(n_709), .C(n_710), .Y(n_707) );
AOI31xp33_ASAP7_75t_L g690 ( .A1(n_685), .A2(n_691), .A3(n_692), .B(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g708 ( .A(n_706), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g719 ( .A(n_714), .Y(n_719) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
endmodule