module real_jpeg_16091_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_216;
wire n_202;
wire n_128;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_0),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_18)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_178),
.B1(n_181),
.B2(n_184),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_2),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_3),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_4),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_5),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_5),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_5),
.A2(n_107),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g363 ( 
.A1(n_5),
.A2(n_107),
.B1(n_364),
.B2(n_369),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_6),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_7),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_7),
.Y(n_89)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_7),
.Y(n_120)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_7),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_7),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_7),
.Y(n_278)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_7),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_7),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_8),
.A2(n_134),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_8),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_8),
.A2(n_138),
.B1(n_256),
.B2(n_259),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_8),
.A2(n_138),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_9),
.A2(n_58),
.B1(n_62),
.B2(n_63),
.Y(n_57)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_9),
.A2(n_62),
.B1(n_99),
.B2(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_9),
.A2(n_62),
.B1(n_289),
.B2(n_294),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_9),
.A2(n_62),
.B1(n_339),
.B2(n_340),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_11),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_186),
.A3(n_190),
.B1(n_191),
.B2(n_195),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_11),
.B(n_37),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_11),
.B(n_83),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_11),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_11),
.B(n_143),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_11),
.A2(n_56),
.B1(n_372),
.B2(n_374),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g379 ( 
.A1(n_11),
.A2(n_380),
.A3(n_382),
.B1(n_383),
.B2(n_387),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g131 ( 
.A(n_13),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_13),
.Y(n_158)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_14),
.A2(n_162),
.B1(n_168),
.B2(n_172),
.Y(n_161)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_14),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_14),
.A2(n_172),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_16),
.A2(n_145),
.B1(n_146),
.B2(n_148),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_16),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_16),
.A2(n_145),
.B1(n_216),
.B2(n_219),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_263),
.B1(n_418),
.B2(n_419),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_22),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_262),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_222),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_24),
.B(n_222),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_150),
.C(n_200),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_25),
.B(n_415),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_65),
.Y(n_25)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_26),
.B(n_66),
.C(n_114),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_50),
.B1(n_57),
.B2(n_64),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_27),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_37),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_36),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_32),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_37),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_243)
);

AO22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_43),
.B2(n_47),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_42),
.Y(n_205)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_42),
.Y(n_377)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_46),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_46),
.Y(n_258)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_55),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_56),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_56),
.B(n_277),
.Y(n_276)
);

OAI21xp33_ASAP7_75t_SL g286 ( 
.A1(n_56),
.A2(n_276),
.B(n_287),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_56),
.A2(n_154),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_56),
.B(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_57),
.Y(n_244)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_60),
.Y(n_197)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_63),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_114),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_94),
.B1(n_105),
.B2(n_113),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_67),
.A2(n_94),
.B1(n_113),
.B2(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_67),
.A2(n_113),
.B1(n_202),
.B2(n_371),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_83),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_77),
.B2(n_80),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_76),
.Y(n_260)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_83)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_85),
.Y(n_287)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_86),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_86),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_87),
.Y(n_316)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_92),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_104),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx2_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_98),
.A2(n_104),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_98),
.A2(n_104),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_98),
.A2(n_104),
.B1(n_282),
.B2(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_103),
.Y(n_381)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_105),
.Y(n_253)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_110),
.Y(n_373)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_112),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_113),
.B(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_133),
.B(n_142),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_115),
.A2(n_127),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_116),
.B(n_144),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_116),
.A2(n_143),
.B1(n_286),
.B2(n_288),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_116),
.A2(n_143),
.B1(n_288),
.B2(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_116),
.A2(n_403),
.B(n_404),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_121),
.B1(n_123),
.B2(n_126),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_120),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_126),
.Y(n_270)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_127),
.B(n_133),
.Y(n_404)
);

OA22x2_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_127)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_128),
.Y(n_301)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_128),
.Y(n_346)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_129),
.Y(n_275)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_130),
.Y(n_311)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_131),
.Y(n_283)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_131),
.Y(n_312)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_143),
.B(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_146),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_149),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_150),
.A2(n_151),
.B1(n_200),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_185),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_152),
.B(n_185),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_161),
.B1(n_173),
.B2(n_177),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_153),
.A2(n_177),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_153),
.A2(n_324),
.B1(n_329),
.B2(n_330),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_153),
.A2(n_226),
.B(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_154),
.B(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_154),
.A2(n_299),
.B(n_305),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_154),
.A2(n_325),
.B1(n_338),
.B2(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_159),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_156),
.Y(n_340)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_157),
.Y(n_304)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_158),
.Y(n_273)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_161),
.A2(n_210),
.B(n_214),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_176),
.Y(n_337)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_200),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.C(n_208),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_201),
.B(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_209),
.Y(n_408)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_210),
.Y(n_352)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_213),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_241),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_240),
.Y(n_223)
);

XOR2x2_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_230),
.Y(n_309)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_231),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_261),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_251),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B(n_254),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_257),
.Y(n_390)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_263),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_411),
.B(n_417),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_397),
.B(n_410),
.Y(n_264)
);

OAI21x1_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_357),
.B(n_396),
.Y(n_265)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_321),
.B(n_356),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_297),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_268),
.B(n_297),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_284),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_269),
.A2(n_284),
.B1(n_285),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_269),
.Y(n_333)
);

OAI32xp33_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.A3(n_274),
.B1(n_276),
.B2(n_279),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_278),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_293),
.Y(n_386)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_313),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_298),
.B(n_314),
.C(n_320),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_299),
.Y(n_329)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_320),
.Y(n_313)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_315),
.Y(n_362)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_334),
.B(n_355),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_332),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_332),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_335),
.A2(n_350),
.B(n_354),
.Y(n_334)
);

NOR2x1_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_341),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_347),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_353),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_353),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_358),
.B(n_359),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_378),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_370),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_370),
.C(n_378),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_363),
.Y(n_403)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_367),
.Y(n_382)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_394),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_394),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_398),
.B(n_399),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_405),
.B1(n_406),
.B2(n_409),
.Y(n_399)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_401),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_402),
.B(n_405),
.C(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_412),
.B(n_414),
.Y(n_417)
);


endmodule