module fake_aes_6407_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
INVx1_ASAP7_75t_SL g15 ( .A(n_10), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_4), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_5), .Y(n_17) );
INVx4_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_12), .Y(n_19) );
AOI21xp5_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_9), .B(n_6), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_12), .A2(n_0), .B(n_1), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_21), .B(n_17), .Y(n_23) );
NOR3xp33_ASAP7_75t_SL g24 ( .A(n_22), .B(n_17), .C(n_11), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_18), .B(n_13), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_23), .Y(n_27) );
NAND2x1p5_ASAP7_75t_L g28 ( .A(n_25), .B(n_18), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_24), .B1(n_12), .B2(n_19), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
OAI211xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_12), .B(n_20), .C(n_28), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g32 ( .A(n_29), .B(n_0), .Y(n_32) );
CKINVDCx5p33_ASAP7_75t_R g33 ( .A(n_32), .Y(n_33) );
NOR2x1_ASAP7_75t_L g34 ( .A(n_31), .B(n_12), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g36 ( .A(n_34), .Y(n_36) );
AOI22xp5_ASAP7_75t_SL g37 ( .A1(n_36), .A2(n_2), .B1(n_5), .B2(n_35), .Y(n_37) );
endmodule