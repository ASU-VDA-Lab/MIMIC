module fake_jpeg_3857_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_32),
.B(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_42),
.B1(n_19),
.B2(n_21),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

AO22x1_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_46),
.B1(n_58),
.B2(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_32),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_53),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_23),
.B1(n_22),
.B2(n_28),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_27),
.B1(n_23),
.B2(n_22),
.Y(n_70)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_55),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_62),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_71),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_44),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_20),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_73),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_84),
.B1(n_30),
.B2(n_26),
.Y(n_95)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_43),
.B(n_31),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_26),
.B1(n_47),
.B2(n_53),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_43),
.A2(n_41),
.B1(n_42),
.B2(n_39),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_90),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_77),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_91),
.A2(n_42),
.B(n_49),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx4_ASAP7_75t_SL g93 ( 
.A(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_71),
.B1(n_78),
.B2(n_64),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_55),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_98),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_70),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_101),
.A2(n_52),
.B1(n_56),
.B2(n_66),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_83),
.B(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_103),
.B(n_64),
.Y(n_116)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_104),
.B(n_66),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_73),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_72),
.B(n_82),
.C(n_76),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_37),
.B(n_39),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_44),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_114),
.A2(n_126),
.B(n_120),
.Y(n_132)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_102),
.Y(n_145)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_125),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_87),
.B1(n_88),
.B2(n_93),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_56),
.B1(n_41),
.B2(n_39),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_122),
.A2(n_52),
.B1(n_106),
.B2(n_100),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_101),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_96),
.B(n_106),
.C(n_94),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_132),
.B(n_148),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_138),
.C(n_147),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_133),
.A2(n_144),
.B1(n_121),
.B2(n_148),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_145),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_127),
.A2(n_106),
.B1(n_87),
.B2(n_37),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_17),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_17),
.B(n_35),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_149),
.B(n_125),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_102),
.B(n_67),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_117),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_111),
.B(n_123),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_35),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_160),
.B1(n_37),
.B2(n_36),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_146),
.B1(n_129),
.B2(n_115),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_110),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_131),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_168),
.B(n_170),
.CI(n_172),
.CON(n_181),
.SN(n_181)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_109),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_134),
.B1(n_130),
.B2(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_130),
.B1(n_112),
.B2(n_67),
.Y(n_175)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_130),
.C(n_112),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_35),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_92),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_178),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_156),
.B1(n_164),
.B2(n_155),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_92),
.B1(n_36),
.B2(n_51),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

XNOR2x1_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_152),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_171),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_191),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_33),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_36),
.B1(n_3),
.B2(n_5),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_36),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_179),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_199),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_165),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_203),
.B(n_205),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_152),
.C(n_170),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_166),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_204),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_160),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_207),
.B(n_173),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_195),
.A2(n_189),
.B1(n_180),
.B2(n_154),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_186),
.B(n_190),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_211),
.A2(n_215),
.B(n_219),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.C(n_220),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_167),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_154),
.B1(n_159),
.B2(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_201),
.B1(n_194),
.B2(n_197),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_162),
.C(n_175),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_205),
.C(n_198),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_199),
.B(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_164),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_230),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_202),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_225),
.B(n_229),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_200),
.B(n_201),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_1),
.C(n_6),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_227),
.A2(n_222),
.B1(n_7),
.B2(n_8),
.Y(n_238)
);

OAI321xp33_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_206),
.A3(n_181),
.B1(n_169),
.B2(n_196),
.C(n_184),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_192),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_228),
.A2(n_217),
.B1(n_220),
.B2(n_181),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_214),
.B1(n_3),
.B2(n_5),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_235),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_238),
.B(n_8),
.Y(n_241)
);

AOI31xp33_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_1),
.A3(n_6),
.B(n_7),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_1),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_6),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_234),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_7),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_241),
.B(n_244),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_9),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_236),
.Y(n_246)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_246),
.A2(n_12),
.B(n_9),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

AOI322xp5_ASAP7_75t_L g248 ( 
.A1(n_243),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_232),
.C2(n_241),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_245),
.C(n_11),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_249),
.B(n_11),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_12),
.Y(n_253)
);


endmodule