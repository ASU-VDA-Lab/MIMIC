module fake_jpeg_19701_n_325 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx8_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_24),
.B(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_15),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_28),
.A2(n_23),
.B1(n_22),
.B2(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_34),
.B(n_12),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_44),
.B1(n_29),
.B2(n_16),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_21),
.C(n_11),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_26),
.B1(n_32),
.B2(n_43),
.Y(n_57)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_55),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_29),
.B1(n_32),
.B2(n_26),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_58),
.B1(n_35),
.B2(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_59),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_35),
.B1(n_40),
.B2(n_39),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_37),
.A2(n_28),
.B1(n_33),
.B2(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_20),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_61),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_50),
.A2(n_45),
.B1(n_38),
.B2(n_43),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_77),
.B1(n_57),
.B2(n_38),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_28),
.B1(n_40),
.B2(n_39),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_71),
.B1(n_58),
.B2(n_63),
.Y(n_91)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_35),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_51),
.CI(n_62),
.CON(n_92),
.SN(n_92)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_84),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_39),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_36),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_52),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_92),
.Y(n_118)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_96),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_51),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_103),
.B(n_97),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_89),
.A2(n_94),
.B1(n_72),
.B2(n_66),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_57),
.C(n_51),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_89),
.C(n_91),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_104),
.B1(n_65),
.B2(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_51),
.B1(n_53),
.B2(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_95),
.B(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_76),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_69),
.A2(n_64),
.B1(n_54),
.B2(n_48),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_66),
.B1(n_36),
.B2(n_27),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_54),
.Y(n_103)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_72),
.B1(n_78),
.B2(n_50),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_64),
.B1(n_48),
.B2(n_45),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_16),
.B(n_22),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_19),
.B(n_14),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_75),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_106),
.A2(n_111),
.B(n_113),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_107),
.A2(n_108),
.B1(n_30),
.B2(n_27),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_80),
.B1(n_72),
.B2(n_74),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_87),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_112),
.B(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_101),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_124),
.B1(n_135),
.B2(n_36),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_34),
.B(n_14),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_88),
.B(n_92),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_127),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_131),
.C(n_104),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_74),
.B1(n_84),
.B2(n_73),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_41),
.C(n_49),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_92),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_78),
.B1(n_66),
.B2(n_70),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_134),
.B1(n_36),
.B2(n_49),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_78),
.B1(n_66),
.B2(n_70),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_88),
.B(n_95),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_146),
.B(n_158),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_137),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_87),
.B1(n_104),
.B2(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_138),
.A2(n_142),
.B1(n_167),
.B2(n_168),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_139),
.B(n_106),
.Y(n_182)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_125),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_92),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_149),
.Y(n_190)
);

AO22x1_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_88),
.B1(n_107),
.B2(n_111),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_15),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_161),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_15),
.B(n_23),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_109),
.B(n_22),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_122),
.B1(n_116),
.B2(n_135),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_162),
.A2(n_170),
.B1(n_49),
.B2(n_30),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_23),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_13),
.B(n_18),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_130),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_164),
.A2(n_171),
.B(n_113),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_41),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_169),
.C(n_115),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_19),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_166),
.A2(n_13),
.B1(n_18),
.B2(n_30),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_108),
.A2(n_19),
.B1(n_33),
.B2(n_31),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_41),
.C(n_49),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_41),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_179),
.B(n_187),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_188),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_SL g183 ( 
.A(n_143),
.B(n_113),
.C(n_115),
.Y(n_183)
);

HB1xp67_ASAP7_75t_SL g222 ( 
.A(n_183),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_184),
.A2(n_200),
.B1(n_168),
.B2(n_173),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_138),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_185),
.A2(n_194),
.B1(n_166),
.B2(n_163),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_165),
.C(n_169),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_49),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_195),
.Y(n_207)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_144),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_11),
.B1(n_21),
.B2(n_13),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_196),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_25),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_136),
.A2(n_13),
.B1(n_12),
.B2(n_25),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_25),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_199),
.B(n_156),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_212),
.B1(n_219),
.B2(n_180),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_218),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_200),
.A2(n_141),
.B(n_145),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_206),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_141),
.B(n_145),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_150),
.B1(n_147),
.B2(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_172),
.B(n_161),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_164),
.Y(n_217)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

OAI22x1_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_149),
.B1(n_159),
.B2(n_148),
.Y(n_219)
);

AO22x1_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_149),
.B1(n_167),
.B2(n_163),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_154),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_224),
.Y(n_245)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_155),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_187),
.C(n_182),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_230),
.C(n_234),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_176),
.C(n_188),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_231),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_193),
.B1(n_199),
.B2(n_151),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_212),
.B1(n_219),
.B2(n_201),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_174),
.C(n_152),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_198),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_236),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_205),
.B(n_185),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_194),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_158),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_202),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_21),
.C(n_11),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_224),
.C(n_206),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_262),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_204),
.B1(n_217),
.B2(n_221),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_253),
.A2(n_254),
.B1(n_264),
.B2(n_242),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_247),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_259),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_237),
.Y(n_258)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_201),
.C(n_208),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_265),
.C(n_241),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_263),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_220),
.Y(n_262)
);

OAI21xp33_ASAP7_75t_SL g263 ( 
.A1(n_246),
.A2(n_220),
.B(n_207),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_228),
.A2(n_207),
.B1(n_213),
.B2(n_21),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_11),
.C(n_18),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_233),
.C(n_236),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_232),
.C(n_227),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_246),
.B1(n_226),
.B2(n_240),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_235),
.C(n_226),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_274),
.B(n_251),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_18),
.C(n_13),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_280),
.A2(n_13),
.B1(n_7),
.B2(n_10),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_268),
.A2(n_250),
.B1(n_265),
.B2(n_252),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_279),
.A2(n_251),
.B1(n_7),
.B2(n_8),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_283),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_7),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_284),
.B(n_286),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_4),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_10),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_270),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_266),
.A2(n_9),
.B(n_8),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_278),
.B(n_275),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_9),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_4),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_277),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_297),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_2),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_302),
.Y(n_310)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_304),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_288),
.A2(n_290),
.B(n_282),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_293),
.B(n_287),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_18),
.C(n_5),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);

O2A1O1Ixp33_ASAP7_75t_SL g316 ( 
.A1(n_306),
.A2(n_294),
.B(n_295),
.C(n_6),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_297),
.C(n_304),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_307),
.B(n_313),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_311),
.C(n_310),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_314),
.B(n_306),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_319),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_4),
.B(n_5),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_4),
.CI(n_5),
.CON(n_324),
.SN(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_5),
.Y(n_325)
);


endmodule