module fake_jpeg_451_n_558 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_558);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_558;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_509;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_13),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_10),
.B(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_17),
.B(n_1),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_62),
.Y(n_160)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_69),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_36),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_70),
.B(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_76),
.Y(n_158)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_19),
.B(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_82),
.Y(n_139)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_45),
.B(n_9),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_19),
.B(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_98),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

BUFx4f_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_22),
.Y(n_89)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_47),
.B(n_18),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_33),
.Y(n_100)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_9),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_102),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_47),
.B(n_9),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_104),
.Y(n_117)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_23),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_38),
.B(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_105),
.B(n_27),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_46),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_34),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_86),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_118),
.B(n_122),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_120),
.A2(n_129),
.B1(n_144),
.B2(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_40),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_41),
.B1(n_39),
.B2(n_42),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_81),
.A2(n_41),
.B1(n_20),
.B2(n_35),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_86),
.A2(n_20),
.B1(n_35),
.B2(n_43),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_73),
.A2(n_49),
.B(n_22),
.C(n_44),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_80),
.B(n_49),
.C(n_83),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_59),
.B(n_40),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_154),
.B(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_155),
.B(n_167),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_65),
.B(n_28),
.Y(n_157)
);

OR2x4_ASAP7_75t_L g162 ( 
.A(n_69),
.B(n_22),
.Y(n_162)
);

OR2x2_ASAP7_75t_SL g222 ( 
.A(n_162),
.B(n_0),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_62),
.A2(n_54),
.B1(n_32),
.B2(n_50),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_163),
.A2(n_44),
.B1(n_48),
.B2(n_56),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_63),
.B(n_28),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_169),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_170),
.B(n_186),
.Y(n_260)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_172),
.B(n_174),
.Y(n_225)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_179),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_117),
.A2(n_151),
.B1(n_143),
.B2(n_136),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_176),
.A2(n_197),
.B(n_214),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_177),
.A2(n_193),
.B(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_178),
.B(n_120),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_114),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_72),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_180),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_27),
.B1(n_106),
.B2(n_85),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_181),
.A2(n_194),
.B1(n_218),
.B2(n_219),
.Y(n_242)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_183),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_121),
.A2(n_20),
.B1(n_35),
.B2(n_51),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_185),
.B(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_140),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_140),
.A2(n_51),
.B1(n_34),
.B2(n_32),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_123),
.C(n_152),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_161),
.C(n_159),
.Y(n_229)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_133),
.Y(n_191)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_191),
.Y(n_272)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_129),
.B(n_148),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_74),
.B1(n_92),
.B2(n_88),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_133),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_196),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_139),
.A2(n_76),
.B1(n_75),
.B2(n_50),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_130),
.B(n_94),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_109),
.B(n_90),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_200),
.B(n_203),
.Y(n_267)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_111),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_137),
.A2(n_51),
.B1(n_50),
.B2(n_23),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_204),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_165),
.B1(n_170),
.B2(n_198),
.Y(n_250)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_111),
.Y(n_208)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_209),
.Y(n_261)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_125),
.Y(n_210)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_210),
.Y(n_269)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_113),
.Y(n_211)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_211),
.Y(n_262)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_213),
.B(n_216),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_115),
.A2(n_44),
.B1(n_48),
.B2(n_2),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_115),
.A2(n_44),
.B1(n_48),
.B2(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_220),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_138),
.A2(n_44),
.B1(n_1),
.B2(n_3),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_11),
.B1(n_1),
.B2(n_4),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_132),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_221),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_222),
.B(n_170),
.Y(n_239)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_108),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_224),
.Y(n_263)
);

BUFx4f_ASAP7_75t_SL g224 ( 
.A(n_142),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_229),
.B(n_6),
.C(n_7),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_230),
.B(n_195),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_153),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_249),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_239),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_205),
.B(n_132),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_244),
.B(n_246),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_197),
.A2(n_164),
.B1(n_158),
.B2(n_134),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_245),
.A2(n_250),
.B1(n_264),
.B2(n_182),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_202),
.B(n_176),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_134),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_164),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_252),
.B(n_270),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_188),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_268),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_206),
.A2(n_146),
.B1(n_145),
.B2(n_138),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_190),
.B(n_145),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_180),
.B(n_108),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_146),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_243),
.Y(n_304)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_274),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_231),
.B(n_224),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_277),
.B(n_282),
.Y(n_320)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_180),
.C(n_198),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_278),
.B(n_307),
.C(n_254),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_240),
.A2(n_193),
.B1(n_177),
.B2(n_191),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_279),
.A2(n_283),
.B1(n_287),
.B2(n_293),
.Y(n_324)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_272),
.Y(n_280)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_280),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_240),
.A2(n_196),
.B1(n_220),
.B2(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_260),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_284),
.B(n_291),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_230),
.A2(n_209),
.B1(n_168),
.B2(n_171),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_285),
.A2(n_290),
.B1(n_295),
.B2(n_301),
.Y(n_338)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_286),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_201),
.B1(n_192),
.B2(n_207),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_265),
.Y(n_288)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_245),
.A2(n_173),
.B1(n_183),
.B2(n_212),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_213),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_233),
.A2(n_208),
.B1(n_223),
.B2(n_186),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_294),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_224),
.B1(n_210),
.B2(n_217),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_247),
.A2(n_11),
.B(n_1),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_296),
.A2(n_232),
.B(n_238),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_225),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_297),
.B(n_312),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_260),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_298),
.B(n_304),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_249),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_315),
.B1(n_234),
.B2(n_254),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_242),
.A2(n_17),
.B1(n_6),
.B2(n_7),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_302),
.Y(n_347)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_266),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_231),
.B(n_5),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_305),
.B(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_306),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_6),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_310),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_239),
.A2(n_12),
.B(n_13),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_SL g326 ( 
.A1(n_309),
.A2(n_314),
.B(n_284),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_267),
.B(n_14),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_311),
.Y(n_357)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_258),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_14),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_14),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_236),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_264),
.A2(n_15),
.B1(n_267),
.B2(n_247),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_263),
.B1(n_269),
.B2(n_266),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_225),
.B(n_15),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_317),
.B(n_318),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_228),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_229),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_321),
.B(n_355),
.C(n_311),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_270),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_326),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_251),
.B1(n_237),
.B2(n_235),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_330),
.B1(n_341),
.B2(n_346),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_288),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_329),
.B(n_334),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_288),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_302),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_335),
.B(n_337),
.Y(n_375)
);

AO22x1_ASAP7_75t_SL g337 ( 
.A1(n_282),
.A2(n_234),
.B1(n_261),
.B2(n_248),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_277),
.A2(n_273),
.B1(n_268),
.B2(n_263),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_342),
.A2(n_343),
.B1(n_298),
.B2(n_300),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_316),
.A2(n_271),
.B1(n_255),
.B2(n_269),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_345),
.B(n_291),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_283),
.A2(n_271),
.B1(n_255),
.B2(n_256),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_302),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_352),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_281),
.B(n_256),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g366 ( 
.A(n_350),
.B(n_289),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_351),
.A2(n_315),
.B1(n_314),
.B2(n_309),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_304),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_293),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_356),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_248),
.C(n_259),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_296),
.A2(n_232),
.B(n_238),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_282),
.A2(n_241),
.B1(n_262),
.B2(n_259),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_359),
.A2(n_290),
.B1(n_285),
.B2(n_318),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_367),
.B1(n_379),
.B2(n_381),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_332),
.B(n_297),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_361),
.B(n_373),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_319),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_362),
.B(n_395),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_289),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_371),
.C(n_377),
.Y(n_411)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_366),
.B(n_325),
.Y(n_406)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_352),
.A2(n_341),
.B1(n_357),
.B2(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_348),
.Y(n_372)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_372),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_331),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_331),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_374),
.B(n_390),
.Y(n_426)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_348),
.Y(n_376)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_376),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_345),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_320),
.A2(n_312),
.B1(n_295),
.B2(n_299),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_384),
.C(n_386),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_320),
.A2(n_343),
.B1(n_342),
.B2(n_324),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_291),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_344),
.Y(n_385)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_385),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_292),
.C(n_307),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_387),
.A2(n_338),
.B1(n_327),
.B2(n_359),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_320),
.A2(n_301),
.B1(n_287),
.B2(n_308),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_388),
.A2(n_394),
.B1(n_346),
.B2(n_330),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_389),
.A2(n_327),
.B(n_335),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_319),
.B(n_310),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_391),
.Y(n_410)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_392),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_322),
.B(n_306),
.C(n_274),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_333),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_324),
.A2(n_314),
.B1(n_294),
.B2(n_317),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_336),
.Y(n_395)
);

XOR2x2_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_333),
.Y(n_397)
);

XNOR2x1_ASAP7_75t_SL g444 ( 
.A(n_397),
.B(n_364),
.Y(n_444)
);

NOR2xp67_ASAP7_75t_R g398 ( 
.A(n_369),
.B(n_333),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_402),
.B(n_406),
.Y(n_441)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_393),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_415),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_322),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_405),
.B(n_409),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_356),
.B(n_351),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_408),
.A2(n_419),
.B(n_428),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_371),
.B(n_358),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_412),
.A2(n_416),
.B1(n_387),
.B2(n_395),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_413),
.A2(n_379),
.B1(n_375),
.B2(n_360),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_382),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_381),
.A2(n_338),
.B1(n_325),
.B2(n_349),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_337),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_427),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_382),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_378),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_337),
.Y(n_422)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_422),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_366),
.B(n_339),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_423),
.B(n_372),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_294),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_383),
.A2(n_334),
.B(n_329),
.Y(n_428)
);

FAx1_ASAP7_75t_SL g429 ( 
.A(n_386),
.B(n_339),
.CI(n_340),
.CON(n_429),
.SN(n_429)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_369),
.Y(n_432)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_431),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_401),
.Y(n_435)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_370),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_445),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_439),
.A2(n_447),
.B1(n_396),
.B2(n_347),
.Y(n_478)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_410),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_411),
.B(n_424),
.C(n_409),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_424),
.C(n_397),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_449),
.Y(n_468)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_425),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_426),
.B(n_392),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_446),
.B(n_458),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_413),
.A2(n_375),
.B1(n_388),
.B2(n_389),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g448 ( 
.A(n_422),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_448),
.A2(n_456),
.B1(n_408),
.B2(n_420),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_411),
.B(n_394),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_450),
.B(n_452),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_416),
.B(n_376),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_455),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_457),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_407),
.B(n_368),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_405),
.B(n_340),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_402),
.B(n_303),
.Y(n_458)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_456),
.A2(n_419),
.B1(n_398),
.B2(n_429),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_460),
.A2(n_432),
.B1(n_447),
.B2(n_439),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_455),
.A2(n_404),
.B1(n_400),
.B2(n_417),
.Y(n_461)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_463),
.B(n_471),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g464 ( 
.A(n_451),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_464),
.B(n_433),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_429),
.B(n_427),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_442),
.B(n_423),
.C(n_406),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_449),
.B(n_404),
.Y(n_473)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_438),
.B(n_418),
.C(n_410),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_457),
.C(n_454),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_478),
.A2(n_479),
.B1(n_444),
.B2(n_430),
.Y(n_496)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_433),
.B(n_347),
.CI(n_331),
.CON(n_479),
.SN(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_438),
.B(n_280),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_443),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_482),
.A2(n_484),
.B1(n_491),
.B2(n_500),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_435),
.B1(n_434),
.B2(n_453),
.Y(n_484)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_486),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_495),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_499),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_494),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_434),
.B1(n_450),
.B2(n_437),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_473),
.B(n_477),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_462),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_496),
.A2(n_481),
.B1(n_479),
.B2(n_470),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_445),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_498),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_286),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_443),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_465),
.A2(n_441),
.B1(n_241),
.B2(n_262),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_491),
.B(n_496),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_501),
.A2(n_509),
.B(n_441),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_494),
.B(n_463),
.C(n_480),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_503),
.B(n_506),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_484),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_504),
.A2(n_510),
.B1(n_515),
.B2(n_507),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_468),
.C(n_471),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_492),
.A2(n_475),
.B(n_466),
.Y(n_509)
);

INVx11_ASAP7_75t_L g510 ( 
.A(n_493),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_483),
.B(n_468),
.C(n_478),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_512),
.B(n_513),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_482),
.A2(n_475),
.B1(n_481),
.B2(n_472),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_460),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_226),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_486),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_517),
.B(n_487),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_505),
.B(n_485),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_518),
.B(n_519),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_505),
.B(n_462),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_520),
.B(n_523),
.Y(n_539)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_509),
.A2(n_500),
.B(n_479),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_522),
.B(n_526),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_502),
.B(n_241),
.Y(n_523)
);

XNOR2x1_ASAP7_75t_SL g524 ( 
.A(n_514),
.B(n_470),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_524),
.B(n_506),
.C(n_517),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_525),
.A2(n_501),
.B1(n_504),
.B2(n_511),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_502),
.B(n_226),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_527),
.B(n_532),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_253),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_531),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_253),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_15),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_533),
.B(n_529),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_516),
.Y(n_537)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_537),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_540),
.B(n_519),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_528),
.B(n_513),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_541),
.A2(n_511),
.B(n_515),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_544),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_539),
.B(n_521),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_545),
.B(n_547),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_535),
.B(n_507),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_548),
.A2(n_536),
.B(n_541),
.Y(n_550)
);

AOI21xp5_ASAP7_75t_SL g553 ( 
.A1(n_550),
.A2(n_551),
.B(n_552),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_546),
.A2(n_542),
.B(n_534),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_553),
.B(n_554),
.C(n_534),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_549),
.B(n_503),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_508),
.C(n_524),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_556),
.A2(n_538),
.B(n_510),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_557),
.B(n_531),
.Y(n_558)
);


endmodule