module real_jpeg_31762_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_469;
wire n_98;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_0),
.Y(n_242)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_0),
.Y(n_327)
);

BUFx12f_ASAP7_75t_L g417 ( 
.A(n_0),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_1),
.A2(n_70),
.B1(n_229),
.B2(n_233),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g315 ( 
.A1(n_1),
.A2(n_70),
.B1(n_316),
.B2(n_321),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_2),
.Y(n_133)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_89),
.B1(n_199),
.B2(n_201),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_3),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_3),
.A2(n_201),
.B1(n_252),
.B2(n_254),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_4),
.A2(n_102),
.B1(n_103),
.B2(n_107),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_4),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_4),
.A2(n_102),
.B1(n_334),
.B2(n_336),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g449 ( 
.A1(n_4),
.A2(n_102),
.B1(n_450),
.B2(n_452),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_4),
.A2(n_102),
.B1(n_471),
.B2(n_474),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_5),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_5),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_5),
.B(n_111),
.Y(n_395)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_5),
.A2(n_429),
.A3(n_432),
.B1(n_437),
.B2(n_443),
.Y(n_428)
);

OAI21xp33_ASAP7_75t_L g507 ( 
.A1(n_5),
.A2(n_75),
.B(n_508),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_5),
.A2(n_371),
.B1(n_558),
.B2(n_562),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_6),
.A2(n_34),
.B1(n_183),
.B2(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_6),
.A2(n_34),
.B1(n_270),
.B2(n_274),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g398 ( 
.A1(n_6),
.A2(n_34),
.B1(n_399),
.B2(n_402),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_135),
.B1(n_136),
.B2(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_7),
.A2(n_135),
.B1(n_375),
.B2(n_378),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g463 ( 
.A1(n_7),
.A2(n_135),
.B1(n_464),
.B2(n_466),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_7),
.A2(n_135),
.B1(n_536),
.B2(n_539),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_8),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_8),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_9),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_10),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_93),
.B1(n_96),
.B2(n_99),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_11),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_11),
.A2(n_99),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_12),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_12),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_176),
.B1(n_220),
.B2(n_223),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_12),
.A2(n_176),
.B1(n_362),
.B2(n_364),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_12),
.A2(n_176),
.B1(n_421),
.B2(n_426),
.Y(n_420)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_14),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_14),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_14),
.A2(n_35),
.B1(n_87),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_14),
.A2(n_87),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_15),
.A2(n_20),
.B(n_582),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_15),
.B(n_583),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_16),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_17),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_18),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_18),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_18),
.Y(n_163)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_18),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_286),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_283),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_244),
.Y(n_23)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_24),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_192),
.C(n_213),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_25),
.B(n_290),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_100),
.C(n_143),
.Y(n_25)
);

XNOR2x1_ASAP7_75t_L g344 ( 
.A(n_26),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_74),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_27),
.B(n_74),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_38),
.B1(n_65),
.B2(n_73),
.Y(n_27)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_28),
.Y(n_366)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_33),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_37),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_38),
.A2(n_73),
.B1(n_203),
.B2(n_208),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_38),
.A2(n_65),
.B1(n_73),
.B2(n_208),
.Y(n_243)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_38),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_38),
.A2(n_449),
.B(n_453),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.Y(n_38)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_39),
.Y(n_257)
);

OAI22x1_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_50),
.Y(n_39)
);

INVx4_ASAP7_75t_L g473 ( 
.A(n_40),
.Y(n_473)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_42),
.Y(n_427)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_42),
.Y(n_465)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_48),
.Y(n_323)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_49),
.Y(n_495)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_59),
.B2(n_62),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g490 ( 
.A(n_57),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_64),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_64),
.Y(n_538)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_69),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_72),
.Y(n_204)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_72),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_72),
.Y(n_363)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_73),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_77),
.B1(n_83),
.B2(n_92),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_75),
.A2(n_92),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_75),
.A2(n_398),
.B(n_403),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_75),
.A2(n_470),
.B(n_508),
.Y(n_531)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OA21x2_ASAP7_75t_L g194 ( 
.A1(n_76),
.A2(n_195),
.B(n_198),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_76),
.A2(n_84),
.B1(n_315),
.B2(n_324),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_76),
.B(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_76),
.A2(n_404),
.B1(n_462),
.B2(n_469),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_80),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g404 ( 
.A(n_77),
.Y(n_404)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_79),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_79),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_79),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_79),
.Y(n_550)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_82),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_82),
.Y(n_485)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g468 ( 
.A(n_91),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_93),
.B(n_515),
.Y(n_514)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_98),
.Y(n_401)
);

AOI22x1_ASAP7_75t_L g345 ( 
.A1(n_100),
.A2(n_144),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_100),
.Y(n_347)
);

AO22x1_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_111),
.B1(n_123),
.B2(n_134),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_101),
.B(n_123),
.Y(n_225)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_110),
.Y(n_224)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_110),
.Y(n_277)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_110),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_111),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_111),
.B(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_111),
.B(n_134),
.Y(n_330)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_124),
.Y(n_123)
);

AOI22x1_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_115),
.Y(n_261)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_121),
.Y(n_310)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

NAND2x1_ASAP7_75t_L g278 ( 
.A(n_123),
.B(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_123),
.B(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_128),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_133),
.Y(n_313)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g304 ( 
.A(n_138),
.Y(n_304)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_142),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_144),
.Y(n_346)
);

OAI21x1_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_171),
.B(n_180),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_145),
.A2(n_333),
.B(n_341),
.Y(n_332)
);

OA21x2_ASAP7_75t_L g556 ( 
.A1(n_145),
.A2(n_341),
.B(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_146),
.A2(n_182),
.B1(n_191),
.B2(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_146),
.A2(n_228),
.B1(n_259),
.B2(n_263),
.Y(n_258)
);

AOI22x1_ASAP7_75t_L g373 ( 
.A1(n_146),
.A2(n_263),
.B1(n_374),
.B2(n_379),
.Y(n_373)
);

NAND2xp33_ASAP7_75t_SL g394 ( 
.A(n_146),
.B(n_172),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_160),
.Y(n_146)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_152),
.B1(n_155),
.B2(n_157),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_149),
.Y(n_446)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_150),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_156),
.Y(n_451)
);

INVx5_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_159),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B1(n_167),
.B2(n_170),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_162),
.Y(n_377)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_162),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_163),
.Y(n_299)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_163),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_163),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_166),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_172),
.B(n_191),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_190),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_188),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_189),
.Y(n_431)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_190),
.A2(n_393),
.B(n_394),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_190),
.B(n_371),
.Y(n_533)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_192),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_202),
.B2(n_212),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_193),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_194),
.B(n_202),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_198),
.Y(n_240)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_203),
.Y(n_249)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_206),
.Y(n_497)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_207),
.Y(n_365)
);

INVx1_ASAP7_75t_SL g539 ( 
.A(n_209),
.Y(n_539)
);

INVx4_ASAP7_75t_SL g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_215),
.B(n_291),
.Y(n_290)
);

XNOR2x1_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_238),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_226),
.B1(n_227),
.B2(n_237),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_225),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_218),
.B(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx4_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_223),
.Y(n_370)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_281),
.C(n_282),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_239),
.B(n_243),
.Y(n_342)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_280),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_265),
.Y(n_245)
);

NAND2x1_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_264),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_258),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_258),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_257),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_250),
.A2(n_257),
.B1(n_361),
.B2(n_366),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_250),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_250),
.B(n_361),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_250),
.A2(n_553),
.B1(n_554),
.B2(n_555),
.Y(n_552)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_257),
.B(n_361),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_257),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_279),
.Y(n_265)
);

NAND2x1_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_278),
.Y(n_267)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_278),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

AO21x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_348),
.B(n_580),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_292),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_289),
.B(n_292),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_342),
.C(n_343),
.Y(n_292)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_328),
.C(n_331),
.Y(n_293)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_358),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_314),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_295),
.B(n_314),
.Y(n_389)
);

AOI32xp33_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_300),
.A3(n_302),
.B1(n_305),
.B2(n_309),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx11_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_305),
.Y(n_372)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_R g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_315),
.B(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_327),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_358)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_333),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_342),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_354),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_349),
.A2(n_405),
.B(n_577),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_355),
.B(n_382),
.Y(n_350)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_351),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

MAJx2_ASAP7_75t_L g577 ( 
.A(n_356),
.B(n_578),
.C(n_579),
.Y(n_577)
);

MAJx2_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_359),
.C(n_380),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_384),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_359),
.A2(n_380),
.B1(n_381),
.B2(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_359),
.Y(n_385)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_367),
.C(n_373),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_373),
.Y(n_388)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_367),
.B(n_388),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_370),
.A2(n_371),
.B(n_372),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_371),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_371),
.B(n_435),
.Y(n_482)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_371),
.A2(n_482),
.B(n_501),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_371),
.B(n_516),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_371),
.B(n_522),
.Y(n_521)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_374),
.Y(n_393)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_377),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_383),
.B(n_386),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_389),
.C(n_390),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_409),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_389),
.A2(n_390),
.B1(n_391),
.B2(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_389),
.Y(n_410)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.C(n_396),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_395),
.B(n_397),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_R g414 ( 
.A(n_398),
.B(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_398),
.A2(n_419),
.B(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_457),
.B(n_575),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_408),
.Y(n_576)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_412),
.B(n_576),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_447),
.C(n_454),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_413),
.A2(n_447),
.B1(n_448),
.B2(n_570),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_413),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_418),
.B(n_428),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx8_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

OAI21xp33_ASAP7_75t_SL g523 ( 
.A1(n_419),
.A2(n_463),
.B(n_524),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_420),
.B(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_425),
.Y(n_478)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_428),
.B(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_440),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_449),
.Y(n_555)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_453),
.B(n_499),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_455),
.B(n_569),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_566),
.B(n_574),
.Y(n_457)
);

O2A1O1Ixp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_528),
.B(n_541),
.C(n_542),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_505),
.B(n_527),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_479),
.Y(n_460)
);

NOR2xp67_ASAP7_75t_L g527 ( 
.A(n_461),
.B(n_479),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_498),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_480),
.B(n_498),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_483),
.B1(n_491),
.B2(n_496),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_484),
.B(n_486),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_486),
.B(n_497),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

OAI21xp33_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_520),
.B(n_526),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_514),
.Y(n_506)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx2_ASAP7_75t_SL g518 ( 
.A(n_519),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_523),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_521),
.B(n_523),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_522),
.A2(n_535),
.B(n_540),
.Y(n_534)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_529),
.B(n_530),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_531),
.B(n_544),
.C(n_545),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_533),
.B(n_534),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_533),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_534),
.Y(n_544)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_535),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_537),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_546),
.Y(n_542)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_543),
.B(n_546),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_551),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_547),
.Y(n_572)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_556),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_552),
.B(n_556),
.C(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_567),
.B(n_573),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_571),
.Y(n_567)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_571),
.Y(n_574)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);


endmodule