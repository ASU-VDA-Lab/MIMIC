module fake_jpeg_15162_n_168 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_51),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_62),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_68),
.Y(n_73)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_75),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_56),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_52),
.B(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_43),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_60),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_68),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_79),
.Y(n_99)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_56),
.B1(n_40),
.B2(n_57),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_82),
.A2(n_57),
.B1(n_54),
.B2(n_53),
.Y(n_104)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_43),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_92),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_71),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_93),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_0),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_98),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_71),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_85),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_75),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_109),
.B1(n_2),
.B2(n_4),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_110),
.B1(n_6),
.B2(n_8),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_0),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_1),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_49),
.C(n_47),
.Y(n_108)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_44),
.B1(n_42),
.B2(n_50),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_126),
.Y(n_133)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_124),
.B(n_107),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_123),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_133),
.B(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_94),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_140),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_116),
.B1(n_99),
.B2(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_91),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_148),
.B(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_144),
.B1(n_113),
.B2(n_131),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_150),
.A2(n_146),
.B1(n_147),
.B2(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_148),
.B(n_106),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_152),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_153),
.B(n_150),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_151),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_154),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_14),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_15),
.B(n_16),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_17),
.B(n_18),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_162),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_163),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_164),
.B(n_21),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_22),
.B(n_23),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_24),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_167),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_168)
);


endmodule