module fake_jpeg_17559_n_36 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_36);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_32;

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_16),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_27)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_6),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_19),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_21),
.B(n_18),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_28),
.B(n_24),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_22),
.C(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_31),
.C(n_27),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_23),
.A3(n_26),
.B1(n_11),
.B2(n_12),
.C1(n_15),
.C2(n_9),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_10),
.B(n_23),
.Y(n_36)
);


endmodule