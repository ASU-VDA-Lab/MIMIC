module fake_jpeg_17399_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

BUFx5_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

INVx8_ASAP7_75t_SL g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_31),
.B(n_15),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_35),
.C(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_1),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_37),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_34),
.B1(n_43),
.B2(n_50),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_62),
.B1(n_58),
.B2(n_52),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_66),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_2),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_3),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_5),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_58),
.A2(n_18),
.B1(n_29),
.B2(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_61),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_4),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_83),
.B(n_30),
.Y(n_88)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_8),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_22),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_13),
.C(n_14),
.Y(n_81)
);

A2O1A1O1Ixp25_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_17),
.B(n_19),
.C(n_20),
.D(n_21),
.Y(n_83)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_88),
.Y(n_91)
);

OAI322xp33_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_82),
.A3(n_80),
.B1(n_89),
.B2(n_87),
.C1(n_85),
.C2(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_90),
.B1(n_89),
.B2(n_81),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_90),
.Y(n_94)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_83),
.B(n_78),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_25),
.Y(n_98)
);


endmodule