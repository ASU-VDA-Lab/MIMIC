module fake_jpeg_20779_n_116 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_116);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_31),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_8),
.B(n_34),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_45),
.Y(n_53)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_56),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_36),
.Y(n_66)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_64),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_50),
.B1(n_45),
.B2(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_69),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_0),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_50),
.B1(n_49),
.B2(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_48),
.B1(n_44),
.B2(n_39),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_82),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_40),
.B(n_38),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_78),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_77),
.B(n_81),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_1),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_1),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_2),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_3),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_3),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_15),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_73),
.B1(n_78),
.B2(n_82),
.Y(n_92)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_11),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_12),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_13),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_100),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.C(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_105),
.A2(n_100),
.B1(n_101),
.B2(n_87),
.Y(n_108)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

AO221x1_ASAP7_75t_L g109 ( 
.A1(n_107),
.A2(n_108),
.B1(n_89),
.B2(n_91),
.C(n_106),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_91),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_97),
.Y(n_111)
);

AOI31xp67_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_19),
.A3(n_21),
.B(n_24),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_25),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_26),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_27),
.B(n_28),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_30),
.Y(n_116)
);


endmodule