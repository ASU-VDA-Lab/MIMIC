module fake_jpeg_3604_n_38 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AOI21xp33_ASAP7_75t_L g7 ( 
.A1(n_4),
.A2(n_3),
.B(n_0),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_5),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_2),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_2),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_20),
.C(n_21),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_5),
.B(n_6),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_6),
.C(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_12),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.C(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_17),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_31)
);

AOI21x1_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_33),
.B(n_34),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_26),
.C(n_30),
.Y(n_36)
);

OAI311xp33_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_10),
.A3(n_13),
.B1(n_8),
.C1(n_0),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_10),
.B1(n_30),
.B2(n_29),
.Y(n_34)
);

AOI322xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_25),
.A3(n_33),
.B1(n_31),
.B2(n_32),
.C1(n_34),
.C2(n_27),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_35),
.Y(n_38)
);


endmodule