module fake_jpeg_17610_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_24),
.B(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_23),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_34),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_65),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_17),
.B1(n_29),
.B2(n_26),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_59),
.A2(n_71),
.B1(n_73),
.B2(n_61),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_38),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_41),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_33),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_33),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_29),
.B1(n_26),
.B2(n_21),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_21),
.B(n_31),
.C(n_30),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_25),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_47),
.A2(n_22),
.B1(n_18),
.B2(n_32),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_74),
.B(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_80),
.B(n_81),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_83),
.B(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_25),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_4),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_57),
.B(n_4),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_32),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_22),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_18),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_5),
.B1(n_49),
.B2(n_66),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_4),
.Y(n_95)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_69),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_103),
.A2(n_79),
.B(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_66),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_108),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_51),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_51),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_98),
.B(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_64),
.B1(n_5),
.B2(n_8),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_81),
.B1(n_95),
.B2(n_85),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_55),
.B(n_8),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_118),
.A2(n_94),
.B(n_77),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_127),
.B(n_130),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_98),
.C(n_85),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_132),
.C(n_104),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_76),
.B(n_74),
.C(n_91),
.Y(n_125)
);

OAI211xp5_ASAP7_75t_SL g149 ( 
.A1(n_125),
.A2(n_117),
.B(n_109),
.C(n_105),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_75),
.B(n_86),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_128),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_93),
.Y(n_129)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_134),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_103),
.B1(n_115),
.B2(n_117),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_75),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_55),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_123),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_114),
.C(n_107),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_136),
.C(n_120),
.Y(n_156)
);

A2O1A1O1Ixp25_ASAP7_75t_L g143 ( 
.A1(n_124),
.A2(n_107),
.B(n_112),
.C(n_118),
.D(n_115),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_130),
.A3(n_125),
.B1(n_97),
.B2(n_109),
.Y(n_161)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_148),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_149),
.A2(n_135),
.B(n_120),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_142),
.B(n_126),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_152),
.B(n_156),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_149),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_119),
.C(n_122),
.Y(n_160)
);

FAx1_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_141),
.CI(n_143),
.CON(n_162),
.SN(n_162)
);

AOI321xp33_ASAP7_75t_L g168 ( 
.A1(n_161),
.A2(n_144),
.A3(n_139),
.B1(n_147),
.B2(n_145),
.C(n_137),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_160),
.C(n_156),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_151),
.B(n_146),
.C(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_163),
.B(n_159),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_150),
.B(n_144),
.C(n_139),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_157),
.B(n_155),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_153),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_97),
.B1(n_10),
.B2(n_11),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_165),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_174),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_154),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_178),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_169),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_165),
.B(n_152),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_176),
.B(n_166),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_7),
.B(n_12),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_183),
.C(n_12),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_179),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_184),
.B(n_185),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_13),
.Y(n_187)
);


endmodule