module real_jpeg_7530_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_1),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_1),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_1),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_1),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_2),
.A2(n_29),
.B1(n_47),
.B2(n_50),
.Y(n_46)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_2),
.A2(n_50),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_2),
.A2(n_50),
.B1(n_147),
.B2(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_2),
.A2(n_50),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_2),
.A2(n_266),
.B(n_269),
.C(n_272),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_2),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_2),
.B(n_99),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_2),
.B(n_308),
.C(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_2),
.B(n_89),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_2),
.B(n_80),
.C(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_2),
.B(n_31),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_3),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_80),
.B1(n_91),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_3),
.A2(n_91),
.B1(n_164),
.B2(n_168),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_4),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_4),
.A2(n_28),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_4),
.A2(n_28),
.B1(n_118),
.B2(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_4),
.A2(n_28),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_5),
.Y(n_103)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_5),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_5),
.Y(n_167)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_7),
.Y(n_179)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_7),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_8),
.Y(n_398)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g271 ( 
.A(n_9),
.Y(n_271)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_11),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_13),
.Y(n_101)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_13),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_13),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_13),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_393),
.B(n_396),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_191),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_190),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_19),
.B(n_136),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_125),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_123),
.B2(n_124),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_52),
.B2(n_53),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_23),
.A2(n_24),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_23),
.A2(n_24),
.B1(n_153),
.B2(n_346),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_24),
.B(n_201),
.C(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_24),
.B(n_153),
.C(n_264),
.Y(n_263)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_46),
.B2(n_51),
.Y(n_24)
);

OA22x2_ASAP7_75t_L g123 ( 
.A1(n_25),
.A2(n_30),
.B1(n_46),
.B2(n_51),
.Y(n_123)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_29),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_30),
.A2(n_46),
.B(n_51),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_31)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_32),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_33),
.Y(n_135)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_34),
.Y(n_159)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_50),
.A2(n_131),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_96),
.B2(n_122),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B1(n_89),
.B2(n_90),
.Y(n_55)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_56),
.Y(n_127)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_63),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_64),
.A2(n_78),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_64),
.A2(n_78),
.B1(n_130),
.B2(n_154),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_64),
.B(n_78),
.Y(n_241)
);

NAND2x1_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_78),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_71),
.B1(n_73),
.B2(n_76),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_75),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

AOI22x1_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_85),
.B2(n_87),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_82),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_96),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_123),
.C(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_96),
.A2(n_122),
.B1(n_126),
.B2(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_120),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_97),
.B(n_186),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_109),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g215 ( 
.A1(n_98),
.A2(n_109),
.B1(n_216),
.B2(n_221),
.Y(n_215)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_110),
.B1(n_120),
.B2(n_144),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_99),
.A2(n_144),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_99),
.B(n_217),
.Y(n_229)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_102),
.B1(n_104),
.B2(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_112),
.B1(n_114),
.B2(n_117),
.Y(n_111)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_103),
.Y(n_239)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_103),
.Y(n_279)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_110),
.B(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_123),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_124),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_123),
.B(n_226),
.C(n_240),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_123),
.A2(n_124),
.B1(n_240),
.B2(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_123),
.A2(n_124),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_123),
.B(n_201),
.C(n_356),
.Y(n_373)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_129),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.C(n_160),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_137),
.Y(n_390)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_142),
.A2(n_143),
.B(n_153),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_152),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_153),
.A2(n_342),
.B1(n_343),
.B2(n_346),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_153),
.Y(n_346)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_159),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_160),
.B(n_389),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B(n_189),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_161),
.B(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_183),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_162),
.A2(n_183),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_162),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_162),
.A2(n_189),
.B1(n_224),
.B2(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_171),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_168),
.Y(n_309)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_170),
.Y(n_237)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_170),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_171),
.B(n_236),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_172),
.A2(n_204),
.B1(n_210),
.B2(n_211),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_172),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_173),
.A2(n_236),
.B1(n_275),
.B2(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_173),
.A2(n_232),
.B1(n_236),
.B2(n_275),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_179),
.Y(n_182)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_179),
.Y(n_294)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_183),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_185),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_387),
.B(n_392),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI211xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_283),
.B(n_381),
.C(n_386),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_253),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_196),
.A2(n_253),
.B(n_382),
.C(n_385),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_242),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_197),
.B(n_242),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_222),
.C(n_225),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_198),
.B(n_222),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_200),
.A2(n_201),
.B1(n_228),
.B2(n_302),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_200),
.B(n_302),
.C(n_323),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_200),
.A2(n_201),
.B1(n_356),
.B2(n_357),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_214),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_203),
.A2(n_214),
.B1(n_215),
.B2(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_231),
.B(n_234),
.Y(n_230)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_209),
.Y(n_292)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_214),
.A2(n_215),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_214),
.A2(n_215),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_215),
.B(n_274),
.C(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_215),
.B(n_338),
.C(n_340),
.Y(n_351)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_259),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_228),
.A2(n_302),
.B1(n_303),
.B2(n_310),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_228),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_228),
.A2(n_230),
.B1(n_302),
.B2(n_372),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_230),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_240),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_252),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_248),
.B(n_250),
.C(n_252),
.Y(n_391)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_254),
.B(n_256),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_261),
.C(n_263),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_263),
.B(n_379),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_264),
.B(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_273),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_265),
.A2(n_273),
.B1(n_274),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_273),
.A2(n_274),
.B1(n_314),
.B2(n_315),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_274),
.B(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_365),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_350),
.B(n_364),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_335),
.B(n_349),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_320),
.B(n_334),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_312),
.B(n_319),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_299),
.B(n_311),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_296),
.B(n_298),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_295),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_300),
.B1(n_344),
.B2(n_345),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_344),
.C(n_346),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_310),
.Y(n_318)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_322),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_333),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_331),
.B2(n_332),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_332),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_348),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_348),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_340),
.B1(n_341),
.B2(n_347),
.Y(n_336)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_337),
.Y(n_347)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_345),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_352),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_358),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_360),
.C(n_361),
.Y(n_374)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_356),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NOR2x1_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_375),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_374),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_374),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_368),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_373),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_373),
.C(n_377),
.Y(n_376)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_375),
.A2(n_383),
.B(n_384),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_378),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_388),
.B(n_391),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx12f_ASAP7_75t_L g397 ( 
.A(n_394),
.Y(n_397)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);


endmodule