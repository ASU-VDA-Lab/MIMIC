module fake_aes_10983_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
AND2x4_ASAP7_75t_L g3 ( .A(n_1), .B(n_2), .Y(n_3) );
BUFx4f_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
BUFx2_ASAP7_75t_SL g5 ( .A(n_3), .Y(n_5) );
NAND2x1p5_ASAP7_75t_L g6 ( .A(n_3), .B(n_0), .Y(n_6) );
NOR2xp67_ASAP7_75t_L g7 ( .A(n_5), .B(n_3), .Y(n_7) );
AOI22xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_6), .B1(n_3), .B2(n_4), .Y(n_8) );
AOI322xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_0), .A3(n_1), .B1(n_2), .B2(n_4), .C1(n_6), .C2(n_3), .Y(n_9) );
AOI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_6), .B1(n_4), .B2(n_2), .Y(n_10) );
AOI222xp33_ASAP7_75t_SL g11 ( .A1(n_10), .A2(n_0), .B1(n_1), .B2(n_4), .C1(n_2), .C2(n_9), .Y(n_11) );
endmodule