module fake_jpeg_3234_n_87 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_87);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_87;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_23),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_25),
.C(n_22),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_27),
.B(n_1),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_30),
.B1(n_29),
.B2(n_27),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_0),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_51),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_41),
.B1(n_37),
.B2(n_27),
.Y(n_55)
);

AND2x6_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_49),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_0),
.Y(n_59)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_38),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_27),
.B1(n_2),
.B2(n_3),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_58),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_38),
.B1(n_2),
.B2(n_3),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_60),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_7),
.C(n_8),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_6),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_13),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_53),
.B(n_59),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_68),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_12),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_18),
.Y(n_73)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_73),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_72),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_75),
.Y(n_82)
);

OAI21x1_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_62),
.B(n_76),
.Y(n_83)
);

AOI322xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_76),
.A3(n_77),
.B1(n_65),
.B2(n_78),
.C1(n_79),
.C2(n_17),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_15),
.Y(n_87)
);


endmodule