module fake_jpeg_19275_n_257 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_10),
.B(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_33),
.B(n_25),
.Y(n_56)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_23),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_25),
.B1(n_21),
.B2(n_17),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_40),
.B1(n_39),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_21),
.B1(n_25),
.B2(n_27),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_43),
.A2(n_22),
.B1(n_20),
.B2(n_16),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_38),
.Y(n_44)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_53),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_56),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_23),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_59),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_19),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_53),
.A2(n_40),
.B(n_39),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_38),
.C(n_35),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_64),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_35),
.C(n_34),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_66),
.B(n_31),
.Y(n_105)
);

AOI32xp33_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_35),
.A3(n_34),
.B1(n_19),
.B2(n_32),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_74),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_25),
.B1(n_39),
.B2(n_34),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_80),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_79),
.Y(n_91)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_34),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_51),
.Y(n_83)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_22),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_54),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_20),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_83),
.A2(n_104),
.B(n_71),
.Y(n_130)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_77),
.B1(n_44),
.B2(n_78),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_89),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_32),
.C(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_61),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_79),
.B(n_66),
.C(n_60),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_46),
.B1(n_49),
.B2(n_22),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_116),
.B1(n_126),
.B2(n_133),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_110),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_88),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_115),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_46),
.B1(n_81),
.B2(n_49),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_87),
.A2(n_65),
.B(n_76),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_130),
.B(n_84),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_88),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_64),
.B1(n_82),
.B2(n_44),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_84),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_30),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_70),
.B1(n_75),
.B2(n_74),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_72),
.B1(n_69),
.B2(n_28),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_130),
.B1(n_96),
.B2(n_86),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_103),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_106),
.B(n_71),
.C(n_30),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_28),
.C(n_26),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_26),
.B1(n_24),
.B2(n_2),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_100),
.Y(n_138)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_100),
.Y(n_139)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_106),
.B1(n_91),
.B2(n_107),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_143),
.B(n_150),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_91),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_84),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_148),
.A2(n_160),
.B(n_133),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g150 ( 
.A(n_112),
.B(n_89),
.C(n_84),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_101),
.B1(n_98),
.B2(n_94),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_120),
.B1(n_118),
.B2(n_121),
.Y(n_161)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_102),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_103),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_116),
.C(n_126),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_165),
.C(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_120),
.C(n_121),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_148),
.B(n_141),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_24),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_172),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_18),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_18),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_181),
.A2(n_141),
.B1(n_157),
.B2(n_156),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_3),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_155),
.C(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_169),
.Y(n_205)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_193),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_134),
.Y(n_191)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_191),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_196),
.B(n_198),
.Y(n_208)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_183),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_154),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_162),
.A2(n_153),
.B1(n_152),
.B2(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_200),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_164),
.Y(n_200)
);

XOR2x2_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_160),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_165),
.B1(n_180),
.B2(n_177),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_167),
.B(n_145),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_202),
.A2(n_166),
.B1(n_153),
.B2(n_145),
.Y(n_213)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_205),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_197),
.B(n_152),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_209),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_201),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_213),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_192),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_188),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_215),
.A2(n_189),
.B1(n_193),
.B2(n_186),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_220),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_210),
.B(n_207),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_225),
.C(n_5),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_182),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_188),
.C(n_184),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_173),
.C(n_172),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_185),
.B1(n_176),
.B2(n_171),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_227),
.B1(n_209),
.B2(n_204),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_208),
.B(n_198),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_232),
.C(n_219),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_206),
.B(n_211),
.C(n_208),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_234),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_231),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_223),
.A2(n_184),
.B(n_6),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_5),
.C(n_6),
.Y(n_233)
);

OAI321xp33_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_236),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_241)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_225),
.B(n_6),
.CI(n_7),
.CON(n_236),
.SN(n_236)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_243),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_222),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_242),
.Y(n_247)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_218),
.B1(n_8),
.B2(n_9),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_7),
.C(n_9),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_237),
.A2(n_229),
.B(n_238),
.Y(n_244)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_233),
.C(n_11),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_247),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_252),
.A2(n_248),
.B(n_251),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_254),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_255),
.A2(n_253),
.B(n_12),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g257 ( 
.A(n_256),
.Y(n_257)
);


endmodule