module fake_jpeg_4880_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_47),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_54),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_32),
.Y(n_91)
);

AO22x1_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_19),
.B1(n_23),
.B2(n_21),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_19),
.B(n_27),
.C(n_24),
.Y(n_100)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_52),
.B(n_71),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_25),
.B1(n_30),
.B2(n_26),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_53),
.A2(n_19),
.B1(n_22),
.B2(n_17),
.Y(n_103)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_57),
.Y(n_101)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_60),
.Y(n_86)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_42),
.A2(n_30),
.B1(n_25),
.B2(n_26),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_33),
.B1(n_37),
.B2(n_31),
.Y(n_83)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_30),
.B1(n_25),
.B2(n_33),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_33),
.B1(n_31),
.B2(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_72),
.B(n_79),
.Y(n_109)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_82),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_76),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_30),
.B1(n_25),
.B2(n_37),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_81),
.B1(n_89),
.B2(n_95),
.Y(n_124)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVxp67_ASAP7_75t_SL g107 ( 
.A(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_31),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_84),
.B1(n_97),
.B2(n_61),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_91),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_45),
.B1(n_16),
.B2(n_34),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_93),
.Y(n_115)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_32),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_79),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_16),
.B1(n_34),
.B2(n_28),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_34),
.B1(n_28),
.B2(n_19),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_24),
.B1(n_19),
.B2(n_29),
.Y(n_97)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_19),
.B(n_29),
.C(n_17),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_104),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_47),
.B(n_65),
.Y(n_123)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_122),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_111),
.B1(n_113),
.B2(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_67),
.B1(n_48),
.B2(n_71),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_94),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_77),
.B(n_48),
.C(n_67),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_118),
.C(n_117),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_69),
.B(n_52),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_73),
.B(n_80),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_69),
.C(n_41),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_47),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_121),
.Y(n_134)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_123),
.A2(n_127),
.B1(n_99),
.B2(n_78),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_47),
.B(n_62),
.C(n_68),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_65),
.B1(n_41),
.B2(n_24),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_24),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_84),
.A2(n_65),
.B1(n_20),
.B2(n_29),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_104),
.B1(n_80),
.B2(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_139),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_140),
.A2(n_162),
.B1(n_125),
.B2(n_132),
.Y(n_171)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_141),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_155),
.B1(n_164),
.B2(n_90),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_29),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_81),
.B1(n_89),
.B2(n_100),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_127),
.B1(n_105),
.B2(n_129),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_148),
.Y(n_167)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_156),
.B(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_86),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_153),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_76),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_163),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_109),
.B(n_94),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_154),
.A2(n_113),
.B(n_131),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_74),
.B1(n_93),
.B2(n_92),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_85),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_118),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_158),
.C(n_124),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_101),
.C(n_76),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_111),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_105),
.Y(n_184)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_161),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_124),
.A2(n_82),
.B1(n_88),
.B2(n_98),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_114),
.B(n_76),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_17),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_178),
.C(n_179),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_185),
.B(n_154),
.Y(n_205)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_156),
.A2(n_128),
.B1(n_106),
.B2(n_113),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_174),
.A2(n_182),
.B1(n_186),
.B2(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_184),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_123),
.C(n_110),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_110),
.C(n_130),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_180),
.A2(n_135),
.B(n_161),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_125),
.B(n_119),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_127),
.B1(n_119),
.B2(n_133),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_114),
.C(n_126),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_199),
.C(n_22),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_188),
.B(n_192),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_178),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_137),
.B(n_20),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_136),
.A2(n_98),
.B1(n_90),
.B2(n_20),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_194),
.B(n_134),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_160),
.B1(n_161),
.B2(n_146),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_20),
.C(n_29),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_22),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_211),
.Y(n_241)
);

XOR2x2_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_164),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_204),
.B(n_186),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_205),
.B(n_217),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_138),
.B(n_150),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_206),
.A2(n_212),
.B1(n_218),
.B2(n_190),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_209),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_222),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_194),
.A2(n_159),
.B(n_148),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_141),
.B1(n_135),
.B2(n_165),
.Y(n_212)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_161),
.B(n_20),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_229),
.B1(n_190),
.B2(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_146),
.Y(n_220)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_181),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_20),
.B1(n_22),
.B2(n_17),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_225),
.B1(n_198),
.B2(n_197),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_168),
.A2(n_22),
.B(n_17),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_198),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_22),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_228),
.C(n_223),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_188),
.A2(n_17),
.B(n_2),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_220),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_233),
.C(n_247),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_232),
.B(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_187),
.C(n_179),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_242),
.B1(n_243),
.B2(n_253),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_214),
.A2(n_174),
.B1(n_180),
.B2(n_167),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_235),
.A2(n_237),
.B(n_217),
.Y(n_273)
);

AOI22x1_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_171),
.B1(n_182),
.B2(n_199),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_206),
.B(n_211),
.Y(n_267)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_246),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_192),
.B1(n_172),
.B2(n_170),
.Y(n_243)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_202),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_177),
.C(n_196),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_226),
.B1(n_218),
.B2(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_9),
.Y(n_251)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_201),
.B(n_1),
.C(n_2),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_225),
.C(n_202),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_208),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_221),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_229),
.B1(n_215),
.B2(n_207),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_210),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_213),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_245),
.B(n_203),
.Y(n_257)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_272),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_260),
.B(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_203),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_264),
.B(n_4),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_205),
.C(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_274),
.C(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_248),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_268),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_241),
.B(n_252),
.Y(n_285)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_224),
.B(n_247),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_219),
.C(n_216),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_242),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_239),
.B1(n_236),
.B2(n_244),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_279),
.A2(n_281),
.B1(n_273),
.B2(n_270),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_259),
.A2(n_235),
.B1(n_232),
.B2(n_236),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_285),
.B(n_274),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_293),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_241),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_227),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_11),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_272),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_11),
.Y(n_292)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_297),
.C(n_293),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_262),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_300),
.Y(n_309)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_278),
.B(n_258),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_304),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_269),
.B1(n_268),
.B2(n_266),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_276),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_256),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_282),
.B(n_256),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_269),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_296),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_310),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_315),
.B(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_306),
.B(n_290),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_312),
.A2(n_313),
.B(n_318),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_297),
.A2(n_284),
.B1(n_283),
.B2(n_285),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_5),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_288),
.C(n_289),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_5),
.C(n_7),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_301),
.B(n_264),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_303),
.B(n_12),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_311),
.A2(n_303),
.B1(n_12),
.B2(n_10),
.Y(n_320)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_321),
.A2(n_328),
.B(n_15),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_327),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_12),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_309),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_314),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_330),
.B(n_328),
.C(n_320),
.Y(n_336)
);

AOI21x1_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_314),
.B(n_10),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_323),
.B(n_15),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_333),
.B(n_7),
.Y(n_337)
);

AOI21x1_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_338),
.B(n_334),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_332),
.B(n_329),
.Y(n_340)
);

NOR4xp25_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_7),
.C(n_8),
.D(n_327),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_341),
.A2(n_8),
.B(n_333),
.Y(n_342)
);


endmodule