module fake_jpeg_24820_n_232 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_232);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_8),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_18),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_41),
.C(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_27),
.Y(n_48)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_1),
.CON(n_41),
.SN(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_10),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_51),
.Y(n_64)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_52),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_55),
.B1(n_26),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_24),
.B1(n_32),
.B2(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_21),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_54),
.A2(n_37),
.B1(n_41),
.B2(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_74),
.B1(n_78),
.B2(n_83),
.Y(n_100)
);

OR2x4_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_18),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_63),
.A2(n_67),
.B(n_81),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_65),
.B(n_70),
.Y(n_89)
);

NAND2x1_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_18),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_77),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_80),
.B1(n_21),
.B2(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_45),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_25),
.B1(n_36),
.B2(n_42),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_80)
);

NAND2x1p5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_46),
.B(n_17),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_19),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_22),
.B1(n_32),
.B2(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_49),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_49),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_1),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_97),
.B(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_87),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_103),
.B1(n_61),
.B2(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_105),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_2),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_50),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_64),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_28),
.Y(n_99)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_104),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_62),
.A2(n_60),
.B1(n_59),
.B2(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_65),
.B(n_20),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_23),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_75),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_64),
.A2(n_27),
.B1(n_49),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_105),
.B1(n_95),
.B2(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_30),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_111),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_106),
.B(n_64),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_115),
.B(n_125),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_73),
.B(n_67),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_97),
.B1(n_103),
.B2(n_88),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_131),
.B1(n_125),
.B2(n_134),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_117),
.A2(n_108),
.A3(n_100),
.B1(n_104),
.B2(n_99),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_84),
.C(n_23),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_72),
.B1(n_68),
.B2(n_77),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_134),
.B1(n_76),
.B2(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_129),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_61),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_87),
.B(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_128),
.B(n_133),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_69),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_66),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_135),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_86),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_14),
.C(n_15),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_88),
.B(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_143),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_119),
.Y(n_162)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_100),
.A3(n_89),
.B1(n_93),
.B2(n_66),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_150),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_126),
.B(n_89),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_141),
.B(n_152),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_145),
.B1(n_154),
.B2(n_114),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_146),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_76),
.B1(n_101),
.B2(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_113),
.Y(n_171)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_118),
.C(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_110),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_102),
.B1(n_92),
.B2(n_84),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_120),
.C(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_132),
.B(n_115),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_156),
.B(n_143),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_162),
.B(n_175),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_124),
.B1(n_115),
.B2(n_119),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_173),
.B1(n_142),
.B2(n_154),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_120),
.Y(n_166)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

OAI32xp33_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_156),
.A3(n_138),
.B1(n_149),
.B2(n_140),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_172),
.Y(n_192)
);

NAND4xp25_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_114),
.C(n_153),
.D(n_157),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_145),
.CI(n_139),
.CON(n_182),
.SN(n_182)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_174),
.B1(n_175),
.B2(n_165),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_165),
.B(n_172),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_155),
.B(n_158),
.C(n_149),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_112),
.B1(n_122),
.B2(n_118),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_185),
.B(n_191),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_160),
.B(n_161),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_180),
.A2(n_183),
.B1(n_187),
.B2(n_189),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_141),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_164),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_184),
.C(n_171),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_167),
.A2(n_136),
.B(n_151),
.C(n_146),
.D(n_150),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_12),
.B(n_15),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_170),
.A2(n_75),
.B1(n_27),
.B2(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_159),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_198),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_197),
.B(n_201),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_179),
.A2(n_162),
.B(n_164),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_203),
.B1(n_192),
.B2(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_186),
.B(n_23),
.Y(n_211)
);

OAI31xp33_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_159),
.A3(n_166),
.B(n_169),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_208),
.C(n_210),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_193),
.A2(n_180),
.B1(n_178),
.B2(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_190),
.C(n_199),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_190),
.B(n_185),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_209),
.A2(n_210),
.B(n_212),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_195),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_11),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_217),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_216),
.B(n_7),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_12),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_12),
.B(n_6),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_23),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_208),
.B(n_6),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_223),
.C(n_7),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_7),
.B(n_10),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_224),
.A2(n_13),
.B(n_14),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_220),
.B1(n_219),
.B2(n_10),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_226),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_SL g229 ( 
.A1(n_227),
.A2(n_228),
.B(n_13),
.C(n_23),
.Y(n_229)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_221),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_3),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_230),
.B(n_3),
.Y(n_232)
);


endmodule