module real_jpeg_6876_n_9 (n_5, n_4, n_8, n_0, n_43, n_1, n_2, n_45, n_6, n_44, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_43;
input n_1;
input n_2;
input n_45;
input n_6;
input n_44;
input n_7;
input n_3;

output n_9;

wire n_17;
wire n_37;
wire n_21;
wire n_35;
wire n_33;
wire n_38;
wire n_29;
wire n_10;
wire n_31;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

NAND3xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_7),
.C(n_12),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_4),
.A2(n_21),
.B(n_43),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_21),
.C(n_45),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_6),
.A2(n_8),
.B(n_21),
.Y(n_20)
);

NAND3xp33_ASAP7_75t_L g39 ( 
.A(n_6),
.B(n_8),
.C(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_19),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_15),
.Y(n_10)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B(n_18),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_24),
.B(n_39),
.Y(n_19)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_29),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_37),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B(n_30),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.C(n_38),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_44),
.Y(n_29)
);


endmodule