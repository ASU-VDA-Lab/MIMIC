module fake_jpeg_29527_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_2),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_0),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_19),
.C(n_42),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_0),
.B(n_1),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_56),
.C(n_60),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_65),
.A2(n_62),
.B1(n_48),
.B2(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_75),
.B1(n_54),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_48),
.B1(n_57),
.B2(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_58),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_51),
.Y(n_79)
);

OR2x2_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_51),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_51),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_1),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_84),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_91),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_93),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_45),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_97),
.Y(n_101)
);

OAI21x1_ASAP7_75t_R g95 ( 
.A1(n_74),
.A2(n_20),
.B(n_41),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_8),
.Y(n_113)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NOR2x1p5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_2),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_80),
.C(n_78),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_103),
.C(n_110),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_3),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_106),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_21),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_111),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_105),
.B(n_27),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_7),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_17),
.C(n_18),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_113),
.A2(n_14),
.B(n_15),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_127),
.B1(n_24),
.B2(n_30),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_124),
.B(n_125),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_105),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_104),
.B(n_29),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_130),
.A2(n_116),
.B(n_34),
.C(n_35),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_31),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_136),
.B(n_137),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_134),
.A2(n_118),
.B(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_133),
.C(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_139),
.B(n_123),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_129),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_131),
.Y(n_143)
);

OAI21x1_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_140),
.B(n_131),
.Y(n_144)
);

NAND4xp25_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_135),
.C(n_104),
.D(n_38),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_33),
.Y(n_146)
);


endmodule