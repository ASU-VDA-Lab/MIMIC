module fake_jpeg_651_n_52 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_52);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_52;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_12),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_11),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_21),
.Y(n_27)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_2),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_14),
.B(n_1),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_25),
.B(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_22),
.A2(n_13),
.B1(n_3),
.B2(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_6),
.B1(n_23),
.B2(n_19),
.Y(n_33)
);

AND2x6_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_20),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_34),
.C(n_35),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_36),
.A2(n_23),
.B(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_40),
.B(n_30),
.C(n_38),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_34),
.C(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_41),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

AOI21x1_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_45),
.B(n_43),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_50),
.B(n_48),
.Y(n_51)
);

INVxp33_ASAP7_75t_SL g52 ( 
.A(n_51),
.Y(n_52)
);


endmodule