module fake_jpeg_1626_n_453 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_453);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_453;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_45),
.Y(n_97)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_47),
.Y(n_111)
);

CKINVDCx9p33_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_55),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_52),
.Y(n_133)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_27),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_54),
.B(n_60),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_27),
.B(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_57),
.Y(n_127)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_59),
.Y(n_143)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_15),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_62),
.Y(n_118)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_22),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_0),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_84),
.Y(n_89)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx11_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_85),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_86),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_21),
.B1(n_40),
.B2(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_107),
.B1(n_113),
.B2(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_32),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_94),
.B(n_104),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_79),
.A2(n_38),
.B1(n_30),
.B2(n_41),
.Y(n_96)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_96),
.A2(n_131),
.B1(n_1),
.B2(n_4),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_58),
.B(n_38),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_21),
.B1(n_40),
.B2(n_34),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_38),
.B1(n_34),
.B2(n_40),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_117),
.B1(n_142),
.B2(n_5),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_70),
.A2(n_29),
.B1(n_28),
.B2(n_24),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_49),
.A2(n_41),
.B1(n_30),
.B2(n_24),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_130),
.B1(n_19),
.B2(n_52),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_71),
.A2(n_29),
.B1(n_20),
.B2(n_24),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_59),
.A2(n_28),
.B1(n_20),
.B2(n_44),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_139),
.B1(n_141),
.B2(n_75),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_50),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_138),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_81),
.A2(n_39),
.B1(n_33),
.B2(n_32),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_63),
.A2(n_69),
.B1(n_39),
.B2(n_31),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_46),
.A2(n_44),
.B(n_39),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_6),
.C(n_8),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_83),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_80),
.A2(n_44),
.B1(n_33),
.B2(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_75),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_1),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_65),
.A2(n_31),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_91),
.B(n_1),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_147),
.B(n_158),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_148),
.B(n_137),
.C(n_120),
.Y(n_218)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_154),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_155),
.B(n_184),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_96),
.A2(n_52),
.B1(n_19),
.B2(n_3),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_156),
.A2(n_161),
.B1(n_172),
.B2(n_183),
.Y(n_206)
);

INVx13_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_157),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_135),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_106),
.Y(n_159)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_112),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_19),
.B1(n_2),
.B2(n_4),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx5_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_117),
.A2(n_101),
.B1(n_128),
.B2(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_163),
.A2(n_92),
.B1(n_105),
.B2(n_122),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_164),
.B(n_169),
.Y(n_230)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_167),
.A2(n_188),
.B1(n_195),
.B2(n_196),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_170),
.B(n_199),
.Y(n_202)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_173),
.A2(n_133),
.B(n_124),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_6),
.C(n_8),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_176),
.C(n_185),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_118),
.B(n_8),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_179),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_9),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_190),
.Y(n_200)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_110),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_109),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_181),
.B(n_186),
.Y(n_231)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_182),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_90),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_89),
.B(n_11),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_101),
.A2(n_11),
.B1(n_12),
.B2(n_140),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_197),
.B1(n_95),
.B2(n_105),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_130),
.A2(n_12),
.B1(n_97),
.B2(n_143),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_104),
.B(n_127),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_133),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_97),
.A2(n_114),
.B1(n_108),
.B2(n_89),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_108),
.A2(n_104),
.B1(n_129),
.B2(n_115),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_198),
.B(n_144),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_123),
.B(n_132),
.Y(n_199)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_174),
.B(n_134),
.CI(n_93),
.CON(n_208),
.SN(n_208)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_218),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_170),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_168),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_213),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_133),
.B(n_134),
.C(n_93),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_215),
.A2(n_195),
.B(n_165),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_132),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_152),
.A2(n_115),
.B1(n_129),
.B2(n_92),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_225),
.B1(n_236),
.B2(n_240),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_136),
.C(n_120),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_222),
.B(n_245),
.C(n_150),
.Y(n_266)
);

OAI211xp5_ASAP7_75t_L g271 ( 
.A1(n_226),
.A2(n_149),
.B(n_157),
.C(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_155),
.B(n_137),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_237),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_162),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_146),
.A2(n_122),
.B1(n_144),
.B2(n_192),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_176),
.B(n_144),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_175),
.B(n_144),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_167),
.B1(n_180),
.B2(n_185),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_161),
.A2(n_185),
.B1(n_167),
.B2(n_180),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_166),
.B1(n_177),
.B2(n_186),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_191),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_159),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_184),
.B(n_190),
.C(n_164),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_252),
.Y(n_308)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_207),
.B(n_159),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_257),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_260),
.B(n_286),
.Y(n_320)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g297 ( 
.A(n_261),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_203),
.A2(n_167),
.B1(n_154),
.B2(n_189),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_262),
.A2(n_221),
.B1(n_209),
.B2(n_232),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_264),
.A2(n_271),
.B(n_280),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_145),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_276),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_223),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_207),
.A2(n_171),
.B(n_179),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_267),
.A2(n_275),
.B(n_208),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_213),
.B(n_194),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_268),
.B(n_272),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_277),
.B1(n_281),
.B2(n_220),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_198),
.C(n_193),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_274),
.C(n_283),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_201),
.B(n_219),
.Y(n_272)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_273),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_203),
.B(n_210),
.C(n_224),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_207),
.A2(n_215),
.B(n_230),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_224),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_206),
.B1(n_205),
.B2(n_212),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_278),
.Y(n_324)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_211),
.B(n_202),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_206),
.A2(n_211),
.B1(n_200),
.B2(n_229),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_217),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_210),
.B(n_200),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_217),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_289),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_238),
.Y(n_286)
);

INVx5_ASAP7_75t_SL g287 ( 
.A(n_204),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_204),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_241),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_288),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_227),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_303),
.B1(n_307),
.B2(n_319),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_291),
.B(n_292),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_248),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_259),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_298),
.B(n_309),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_289),
.B(n_241),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_299),
.B(n_301),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_246),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_236),
.B1(n_240),
.B2(n_247),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_226),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_314),
.C(n_321),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_247),
.B1(n_208),
.B2(n_225),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_255),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_310),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_255),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_312),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_316),
.A2(n_317),
.B1(n_308),
.B2(n_293),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_263),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_221),
.Y(n_318)
);

OAI21xp33_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_261),
.B(n_250),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_253),
.A2(n_209),
.B1(n_223),
.B2(n_228),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_286),
.Y(n_321)
);

OAI32xp33_ASAP7_75t_L g322 ( 
.A1(n_276),
.A2(n_228),
.A3(n_242),
.B1(n_260),
.B2(n_265),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_322),
.A2(n_300),
.B(n_319),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_253),
.A2(n_279),
.B1(n_275),
.B2(n_262),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_323),
.A2(n_290),
.B1(n_303),
.B2(n_307),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_328),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_306),
.A2(n_264),
.B(n_280),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_329),
.A2(n_339),
.B(n_343),
.Y(n_363)
);

NOR4xp25_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_326),
.C(n_258),
.D(n_311),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_SL g380 ( 
.A(n_330),
.B(n_346),
.C(n_331),
.Y(n_380)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_266),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_341),
.C(n_342),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_258),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_338),
.Y(n_364)
);

OAI32xp33_ASAP7_75t_L g336 ( 
.A1(n_296),
.A2(n_251),
.A3(n_249),
.B1(n_256),
.B2(n_252),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_267),
.B(n_256),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_345),
.B1(n_353),
.B2(n_297),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_270),
.C(n_269),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_282),
.C(n_285),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_310),
.A2(n_249),
.B(n_287),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_305),
.B(n_326),
.C(n_320),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_347),
.C(n_349),
.Y(n_375)
);

A2O1A1O1Ixp25_ASAP7_75t_L g346 ( 
.A1(n_296),
.A2(n_287),
.B(n_284),
.C(n_257),
.D(n_273),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_320),
.B(n_323),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_300),
.A2(n_292),
.B(n_312),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_291),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_298),
.B(n_315),
.C(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_308),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_355),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_300),
.B(n_324),
.C(n_295),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_352),
.B(n_313),
.Y(n_368)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_334),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_377),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_325),
.Y(n_362)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_344),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_338),
.B(n_304),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_366),
.B(n_368),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_313),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_369),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_333),
.B(n_313),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_335),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_297),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_371),
.A2(n_373),
.B1(n_376),
.B2(n_380),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_372),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_350),
.A2(n_297),
.B1(n_355),
.B2(n_345),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_328),
.A2(n_297),
.B1(n_354),
.B2(n_329),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_356),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_379),
.B(n_348),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_360),
.B(n_341),
.C(n_342),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_382),
.B(n_393),
.C(n_375),
.Y(n_402)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_358),
.A2(n_352),
.B1(n_347),
.B2(n_354),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_387),
.A2(n_397),
.B1(n_367),
.B2(n_361),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_389),
.C(n_393),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_364),
.B(n_366),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_400),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_395),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_339),
.C(n_343),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_367),
.B(n_332),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_373),
.A2(n_336),
.B1(n_351),
.B2(n_346),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g398 ( 
.A(n_359),
.B(n_379),
.CI(n_377),
.CON(n_398),
.SN(n_398)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_383),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_370),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_404),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_392),
.B(n_386),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_407),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_386),
.A2(n_361),
.B1(n_371),
.B2(n_365),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_368),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_363),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_408),
.B(n_410),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_363),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_382),
.B(n_374),
.C(n_378),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_411),
.B(n_413),
.C(n_414),
.Y(n_426)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_394),
.Y(n_412)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_412),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_374),
.C(n_378),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_380),
.Y(n_414)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_415),
.Y(n_429)
);

AOI21x1_ASAP7_75t_SL g422 ( 
.A1(n_416),
.A2(n_398),
.B(n_394),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_389),
.B(n_383),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_417),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_409),
.A2(n_385),
.B(n_398),
.Y(n_419)
);

INVxp33_ASAP7_75t_L g432 ( 
.A(n_419),
.Y(n_432)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_422),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_401),
.A2(n_399),
.B(n_397),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_423),
.A2(n_399),
.B1(n_396),
.B2(n_417),
.Y(n_433)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_411),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_427),
.B(n_407),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_426),
.B(n_413),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_435),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_428),
.B(n_402),
.C(n_406),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_431),
.B(n_433),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_434),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_406),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_418),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_438),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_421),
.B(n_415),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_432),
.A2(n_419),
.B(n_422),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_440),
.A2(n_432),
.B(n_429),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_436),
.A2(n_418),
.B1(n_423),
.B2(n_420),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_440),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_439),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_L g448 ( 
.A(n_447),
.B(n_442),
.C(n_441),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_448),
.B(n_444),
.C(n_430),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_449),
.B(n_435),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_451),
.A2(n_431),
.B1(n_429),
.B2(n_428),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_452),
.B(n_425),
.Y(n_453)
);


endmodule