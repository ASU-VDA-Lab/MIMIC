module fake_jpeg_17400_n_202 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_13),
.Y(n_21)
);

AOI21xp33_ASAP7_75t_L g22 ( 
.A1(n_8),
.A2(n_1),
.B(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_1),
.A2(n_2),
.B(n_13),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_9),
.B(n_4),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_19),
.A2(n_22),
.B1(n_34),
.B2(n_18),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_23),
.B1(n_27),
.B2(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_45),
.Y(n_62)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_6),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_52),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_25),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_35),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_54),
.Y(n_65)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_11),
.Y(n_52)
);

CKINVDCx9p33_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_6),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_57),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_22),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_15),
.B(n_7),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_16),
.A2(n_35),
.B(n_23),
.C(n_31),
.Y(n_59)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_30),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_68),
.B(n_69),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_30),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_72),
.B(n_81),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_75),
.A2(n_61),
.B(n_90),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_74),
.B1(n_76),
.B2(n_62),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_17),
.Y(n_80)
);

INVx2_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_38),
.B(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_56),
.B(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_64),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_24),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_80),
.A2(n_50),
.B(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_45),
.B1(n_58),
.B2(n_49),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_48),
.B1(n_51),
.B2(n_24),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_73),
.A2(n_48),
.B(n_51),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_99),
.C(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_97),
.B(n_110),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_73),
.C(n_70),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_73),
.B(n_74),
.C(n_86),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_75),
.A2(n_82),
.B1(n_63),
.B2(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_88),
.B1(n_87),
.B2(n_85),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_85),
.B1(n_60),
.B2(n_87),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_60),
.A2(n_64),
.B1(n_91),
.B2(n_66),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_89),
.C(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_67),
.C(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_119),
.B1(n_120),
.B2(n_93),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_114),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_80),
.B1(n_14),
.B2(n_19),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_46),
.C(n_68),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_99),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_125),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_111),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_103),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_129),
.B(n_141),
.Y(n_149)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_136),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_133),
.B1(n_126),
.B2(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_139),
.B(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_98),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_93),
.B(n_117),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_104),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_94),
.B1(n_95),
.B2(n_103),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_127),
.B1(n_137),
.B2(n_140),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_164),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_93),
.B(n_118),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_150),
.A2(n_161),
.B(n_163),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_154),
.B(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_104),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_144),
.B(n_129),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_162),
.A2(n_145),
.B(n_133),
.C(n_127),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_165),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_153),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_171),
.C(n_174),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_169),
.A2(n_164),
.B1(n_154),
.B2(n_163),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_128),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_156),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_142),
.C(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_134),
.C(n_138),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_176),
.B(n_177),
.C(n_159),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_136),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_179),
.Y(n_190)
);

AO21x1_ASAP7_75t_L g179 ( 
.A1(n_170),
.A2(n_150),
.B(n_146),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_172),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_156),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_186),
.B(n_185),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_183),
.A2(n_169),
.B1(n_155),
.B2(n_152),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_171),
.C(n_174),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_159),
.C(n_176),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_189),
.C(n_169),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_172),
.C(n_177),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_180),
.B(n_184),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_193),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_194),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_181),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_197),
.A3(n_190),
.B1(n_166),
.B2(n_169),
.C1(n_188),
.C2(n_196),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_201),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_196),
.C(n_195),
.Y(n_201)
);


endmodule