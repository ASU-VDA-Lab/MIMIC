module real_aes_7813_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g450 ( .A(n_0), .Y(n_450) );
INVx1_ASAP7_75t_L g500 ( .A(n_1), .Y(n_500) );
INVx1_ASAP7_75t_L g193 ( .A(n_2), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_3), .A2(n_37), .B1(n_165), .B2(n_509), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g204 ( .A1(n_4), .A2(n_122), .B(n_205), .Y(n_204) );
AOI22xp5_ASAP7_75t_SL g457 ( .A1(n_5), .A2(n_448), .B1(n_458), .B2(n_746), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_6), .B(n_152), .Y(n_492) );
AND2x6_ASAP7_75t_L g127 ( .A(n_7), .B(n_128), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_8), .A2(n_173), .B(n_174), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_9), .B(n_38), .Y(n_451) );
INVx1_ASAP7_75t_L g754 ( .A(n_9), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_10), .B(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g210 ( .A(n_11), .Y(n_210) );
INVx1_ASAP7_75t_L g148 ( .A(n_12), .Y(n_148) );
INVx1_ASAP7_75t_L g496 ( .A(n_13), .Y(n_496) );
INVx1_ASAP7_75t_L g181 ( .A(n_14), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_15), .B(n_196), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_16), .B(n_144), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_17), .A2(n_41), .B1(n_742), .B2(n_743), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_17), .Y(n_743) );
AO32x2_ASAP7_75t_L g506 ( .A1(n_18), .A2(n_143), .A3(n_152), .B1(n_478), .B2(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_19), .B(n_165), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_20), .B(n_138), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_21), .B(n_144), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_22), .A2(n_50), .B1(n_165), .B2(n_509), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_23), .B(n_122), .Y(n_121) );
AOI22xp33_ASAP7_75t_SL g545 ( .A1(n_24), .A2(n_78), .B1(n_165), .B2(n_196), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_25), .B(n_165), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_26), .B(n_203), .Y(n_231) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_27), .A2(n_178), .B(n_180), .C(n_182), .Y(n_177) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_28), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_29), .B(n_156), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_30), .B(n_163), .Y(n_194) );
INVx1_ASAP7_75t_L g220 ( .A(n_31), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_32), .B(n_156), .Y(n_522) );
INVx2_ASAP7_75t_L g125 ( .A(n_33), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_34), .B(n_165), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_35), .B(n_156), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g129 ( .A1(n_36), .A2(n_127), .B(n_130), .C(n_133), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_38), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g218 ( .A(n_39), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_40), .B(n_163), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_41), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g737 ( .A1(n_42), .A2(n_738), .B1(n_739), .B2(n_745), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_42), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_43), .B(n_165), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_44), .A2(n_89), .B1(n_141), .B2(n_509), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_45), .B(n_165), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_46), .B(n_165), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g221 ( .A(n_47), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_48), .B(n_476), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_49), .B(n_122), .Y(n_166) );
AOI22xp33_ASAP7_75t_SL g557 ( .A1(n_51), .A2(n_61), .B1(n_165), .B2(n_196), .Y(n_557) );
AOI22xp33_ASAP7_75t_SL g104 ( .A1(n_52), .A2(n_105), .B1(n_749), .B2(n_759), .Y(n_104) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_53), .A2(n_130), .B1(n_196), .B2(n_217), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_54), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_55), .B(n_165), .Y(n_477) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_56), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_57), .B(n_165), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_58), .A2(n_208), .B(n_209), .C(n_211), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_59), .Y(n_258) );
INVx1_ASAP7_75t_L g206 ( .A(n_60), .Y(n_206) );
INVx1_ASAP7_75t_L g128 ( .A(n_62), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_63), .B(n_165), .Y(n_501) );
INVx1_ASAP7_75t_L g147 ( .A(n_64), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_65), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_66), .A2(n_75), .B1(n_443), .B2(n_444), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g443 ( .A(n_66), .Y(n_443) );
AO32x2_ASAP7_75t_L g542 ( .A1(n_66), .A2(n_152), .A3(n_155), .B1(n_478), .B2(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g474 ( .A(n_67), .Y(n_474) );
INVx1_ASAP7_75t_L g517 ( .A(n_68), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_SL g228 ( .A1(n_69), .A2(n_138), .B(n_211), .C(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_L g230 ( .A(n_70), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_71), .B(n_196), .Y(n_518) );
INVx1_ASAP7_75t_L g758 ( .A(n_72), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_73), .Y(n_223) );
INVx1_ASAP7_75t_L g251 ( .A(n_74), .Y(n_251) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_75), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_76), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g439 ( .A1(n_77), .A2(n_91), .B1(n_440), .B2(n_441), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_77), .Y(n_440) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_79), .A2(n_127), .B(n_130), .C(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_80), .B(n_509), .Y(n_531) );
OAI22xp5_ASAP7_75t_SL g739 ( .A1(n_81), .A2(n_740), .B1(n_741), .B2(n_744), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_81), .Y(n_744) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_82), .B(n_196), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_83), .B(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g145 ( .A(n_84), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_85), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_86), .B(n_196), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_87), .A2(n_127), .B(n_130), .C(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g447 ( .A(n_88), .B(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g461 ( .A(n_88), .Y(n_461) );
NAND3xp33_ASAP7_75t_SL g755 ( .A(n_88), .B(n_450), .C(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_90), .A2(n_103), .B1(n_196), .B2(n_197), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_91), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_92), .B(n_156), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_93), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g158 ( .A1(n_94), .A2(n_127), .B(n_130), .C(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_95), .Y(n_168) );
INVx1_ASAP7_75t_L g227 ( .A(n_96), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_97), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_98), .B(n_135), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_99), .B(n_196), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_100), .B(n_152), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_101), .A2(n_122), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_102), .B(n_758), .Y(n_757) );
AOI22x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B1(n_455), .B2(n_457), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g456 ( .A(n_107), .Y(n_456) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_445), .B(n_452), .Y(n_110) );
XOR2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_442), .Y(n_111) );
OAI22xp5_ASAP7_75t_SL g112 ( .A1(n_113), .A2(n_114), .B1(n_438), .B2(n_439), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g459 ( .A1(n_114), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
AND2x2_ASAP7_75t_SL g114 ( .A(n_115), .B(n_407), .Y(n_114) );
NOR3xp33_ASAP7_75t_L g115 ( .A(n_116), .B(n_300), .C(n_373), .Y(n_115) );
OAI211xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_185), .B(n_232), .C(n_284), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_153), .Y(n_118) );
AND2x2_ASAP7_75t_L g248 ( .A(n_119), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g267 ( .A(n_119), .Y(n_267) );
INVx2_ASAP7_75t_L g282 ( .A(n_119), .Y(n_282) );
INVx1_ASAP7_75t_L g312 ( .A(n_119), .Y(n_312) );
AND2x2_ASAP7_75t_L g362 ( .A(n_119), .B(n_283), .Y(n_362) );
AOI32xp33_ASAP7_75t_L g389 ( .A1(n_119), .A2(n_317), .A3(n_390), .B1(n_392), .B2(n_393), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_119), .B(n_238), .Y(n_395) );
AND2x2_ASAP7_75t_L g422 ( .A(n_119), .B(n_265), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_119), .B(n_431), .Y(n_430) );
OR2x6_ASAP7_75t_L g119 ( .A(n_120), .B(n_149), .Y(n_119) );
AOI21xp5_ASAP7_75t_SL g120 ( .A1(n_121), .A2(n_129), .B(n_142), .Y(n_120) );
BUFx2_ASAP7_75t_L g173 ( .A(n_122), .Y(n_173) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_127), .Y(n_122) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_123), .B(n_127), .Y(n_190) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_126), .Y(n_123) );
INVx1_ASAP7_75t_L g476 ( .A(n_124), .Y(n_476) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g131 ( .A(n_125), .Y(n_131) );
INVx1_ASAP7_75t_L g197 ( .A(n_125), .Y(n_197) );
INVx1_ASAP7_75t_L g132 ( .A(n_126), .Y(n_132) );
INVx3_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
INVx1_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_126), .Y(n_163) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_126), .Y(n_179) );
INVx4_ASAP7_75t_SL g183 ( .A(n_127), .Y(n_183) );
BUFx3_ASAP7_75t_L g478 ( .A(n_127), .Y(n_478) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_127), .A2(n_485), .B(n_488), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_127), .A2(n_495), .B(n_499), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_127), .A2(n_516), .B(n_519), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_127), .A2(n_525), .B(n_529), .Y(n_524) );
INVx5_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx3_ASAP7_75t_L g141 ( .A(n_131), .Y(n_141) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_131), .Y(n_165) );
INVx1_ASAP7_75t_L g509 ( .A(n_131), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_137), .B(n_139), .Y(n_133) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_135), .A2(n_193), .B(n_194), .C(n_195), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_135), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_135), .A2(n_486), .B(n_487), .Y(n_485) );
INVx2_ASAP7_75t_L g491 ( .A(n_135), .Y(n_491) );
O2A1O1Ixp5_ASAP7_75t_SL g516 ( .A1(n_135), .A2(n_211), .B(n_517), .C(n_518), .Y(n_516) );
INVx5_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_136), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_136), .B(n_230), .Y(n_229) );
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_136), .A2(n_163), .B1(n_544), .B2(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g528 ( .A(n_138), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_139), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
INVx1_ASAP7_75t_L g256 ( .A(n_142), .Y(n_256) );
OA21x2_ASAP7_75t_L g468 ( .A1(n_142), .A2(n_469), .B(n_479), .Y(n_468) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_142), .A2(n_494), .B(n_502), .Y(n_493) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AO21x2_ASAP7_75t_L g187 ( .A1(n_143), .A2(n_188), .B(n_198), .Y(n_187) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_143), .A2(n_215), .B(n_222), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_143), .B(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_145), .B(n_146), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
NOR2xp33_ASAP7_75t_SL g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx3_ASAP7_75t_L g203 ( .A(n_151), .Y(n_203) );
AO21x1_ASAP7_75t_L g554 ( .A1(n_151), .A2(n_555), .B(n_558), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g579 ( .A(n_151), .B(n_478), .C(n_555), .Y(n_579) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_152), .A2(n_225), .B(n_231), .Y(n_224) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_152), .A2(n_484), .B(n_492), .Y(n_483) );
AND2x2_ASAP7_75t_L g311 ( .A(n_153), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g333 ( .A(n_153), .Y(n_333) );
AND2x2_ASAP7_75t_L g418 ( .A(n_153), .B(n_248), .Y(n_418) );
AND2x2_ASAP7_75t_L g421 ( .A(n_153), .B(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g153 ( .A(n_154), .B(n_170), .Y(n_153) );
INVx2_ASAP7_75t_L g240 ( .A(n_154), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_154), .B(n_265), .Y(n_271) );
AND2x2_ASAP7_75t_L g281 ( .A(n_154), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g317 ( .A(n_154), .Y(n_317) );
AO21x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_167), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_156), .A2(n_172), .B(n_184), .Y(n_171) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_156), .A2(n_515), .B(n_522), .Y(n_514) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_156), .A2(n_524), .B(n_532), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_158), .B(n_166), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_164), .Y(n_159) );
INVx4_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g208 ( .A(n_163), .Y(n_208) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_163), .A2(n_491), .B1(n_508), .B2(n_510), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_163), .A2(n_491), .B1(n_556), .B2(n_557), .Y(n_555) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx3_ASAP7_75t_L g211 ( .A(n_165), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_169), .B(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_169), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g259 ( .A(n_170), .B(n_240), .Y(n_259) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g241 ( .A(n_171), .Y(n_241) );
AND2x2_ASAP7_75t_L g283 ( .A(n_171), .B(n_265), .Y(n_283) );
AND2x2_ASAP7_75t_L g352 ( .A(n_171), .B(n_249), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .C(n_183), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_176), .A2(n_183), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_176), .A2(n_183), .B(n_227), .C(n_228), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_178), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g498 ( .A(n_178), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_178), .A2(n_520), .B(n_521), .Y(n_519) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g217 ( .A1(n_179), .A2(n_218), .B1(n_219), .B2(n_220), .Y(n_217) );
INVx2_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
OAI22xp33_ASAP7_75t_L g215 ( .A1(n_183), .A2(n_190), .B1(n_216), .B2(n_221), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_200), .Y(n_185) );
OR2x2_ASAP7_75t_L g246 ( .A(n_186), .B(n_214), .Y(n_246) );
INVx1_ASAP7_75t_L g325 ( .A(n_186), .Y(n_325) );
AND2x2_ASAP7_75t_L g339 ( .A(n_186), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_186), .B(n_213), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_186), .B(n_337), .Y(n_391) );
AND2x2_ASAP7_75t_L g399 ( .A(n_186), .B(n_400), .Y(n_399) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx3_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
AND2x2_ASAP7_75t_L g306 ( .A(n_187), .B(n_214), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_190), .A2(n_251), .B(n_252), .Y(n_250) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_195), .A2(n_496), .B(n_497), .C(n_498), .Y(n_495) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_200), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g433 ( .A(n_200), .Y(n_433) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_213), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_201), .B(n_277), .Y(n_299) );
OR2x2_ASAP7_75t_L g328 ( .A(n_201), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g360 ( .A(n_201), .B(n_340), .Y(n_360) );
INVx1_ASAP7_75t_SL g380 ( .A(n_201), .Y(n_380) );
AND2x2_ASAP7_75t_L g384 ( .A(n_201), .B(n_245), .Y(n_384) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_SL g237 ( .A(n_202), .B(n_213), .Y(n_237) );
AND2x2_ASAP7_75t_L g244 ( .A(n_202), .B(n_224), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_202), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g287 ( .A(n_202), .B(n_269), .Y(n_287) );
INVx1_ASAP7_75t_SL g294 ( .A(n_202), .Y(n_294) );
BUFx2_ASAP7_75t_L g305 ( .A(n_202), .Y(n_305) );
AND2x2_ASAP7_75t_L g321 ( .A(n_202), .B(n_236), .Y(n_321) );
AND2x2_ASAP7_75t_L g336 ( .A(n_202), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g400 ( .A(n_202), .B(n_214), .Y(n_400) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_212), .Y(n_202) );
O2A1O1Ixp5_ASAP7_75t_L g473 ( .A1(n_208), .A2(n_474), .B(n_475), .C(n_477), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_208), .A2(n_530), .B(n_531), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_213), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g324 ( .A(n_213), .B(n_325), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_213), .A2(n_342), .B1(n_345), .B2(n_348), .C(n_353), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_213), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
INVx3_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
BUFx2_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
AND2x2_ASAP7_75t_L g293 ( .A(n_224), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g310 ( .A(n_224), .Y(n_310) );
OR2x2_ASAP7_75t_L g329 ( .A(n_224), .B(n_269), .Y(n_329) );
INVx3_ASAP7_75t_L g337 ( .A(n_224), .Y(n_337) );
AND2x2_ASAP7_75t_L g340 ( .A(n_224), .B(n_269), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_238), .B1(n_242), .B2(n_247), .C(n_260), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_235), .B(n_309), .Y(n_434) );
OR2x2_ASAP7_75t_L g437 ( .A(n_235), .B(n_268), .Y(n_437) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
OAI221xp5_ASAP7_75t_SL g260 ( .A1(n_236), .A2(n_261), .B1(n_268), .B2(n_270), .C(n_273), .Y(n_260) );
AND2x2_ASAP7_75t_L g277 ( .A(n_236), .B(n_269), .Y(n_277) );
AND2x2_ASAP7_75t_L g285 ( .A(n_236), .B(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_236), .B(n_293), .Y(n_292) );
NAND2x1_ASAP7_75t_L g335 ( .A(n_236), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g387 ( .A(n_236), .B(n_329), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_238), .A2(n_347), .B1(n_376), .B2(n_378), .Y(n_375) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI322xp5_ASAP7_75t_L g284 ( .A1(n_239), .A2(n_248), .A3(n_285), .B1(n_288), .B2(n_291), .C1(n_295), .C2(n_298), .Y(n_284) );
OR2x2_ASAP7_75t_L g296 ( .A(n_239), .B(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_240), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g275 ( .A(n_240), .B(n_249), .Y(n_275) );
INVx1_ASAP7_75t_L g290 ( .A(n_240), .Y(n_290) );
AND2x2_ASAP7_75t_L g356 ( .A(n_240), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g266 ( .A(n_241), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g357 ( .A(n_241), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_241), .B(n_265), .Y(n_431) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_245), .B(n_380), .Y(n_379) );
INVx3_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g331 ( .A(n_246), .B(n_278), .Y(n_331) );
OR2x2_ASAP7_75t_L g428 ( .A(n_246), .B(n_279), .Y(n_428) );
INVx1_ASAP7_75t_L g409 ( .A(n_247), .Y(n_409) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_259), .Y(n_247) );
INVx4_ASAP7_75t_L g297 ( .A(n_248), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_248), .B(n_316), .Y(n_322) );
INVx2_ASAP7_75t_L g265 ( .A(n_249), .Y(n_265) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_256), .B(n_257), .Y(n_249) );
INVx1_ASAP7_75t_L g347 ( .A(n_259), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_259), .B(n_319), .Y(n_388) );
AOI21xp33_ASAP7_75t_L g334 ( .A1(n_261), .A2(n_335), .B(n_338), .Y(n_334) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g319 ( .A(n_265), .Y(n_319) );
INVx1_ASAP7_75t_L g346 ( .A(n_265), .Y(n_346) );
INVx1_ASAP7_75t_L g272 ( .A(n_266), .Y(n_272) );
AND2x2_ASAP7_75t_L g274 ( .A(n_266), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g370 ( .A(n_267), .B(n_356), .Y(n_370) );
AND2x2_ASAP7_75t_L g392 ( .A(n_267), .B(n_352), .Y(n_392) );
BUFx2_ASAP7_75t_L g344 ( .A(n_269), .Y(n_344) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
AOI32xp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_276), .A3(n_277), .B1(n_278), .B2(n_280), .Y(n_273) );
INVx1_ASAP7_75t_L g354 ( .A(n_274), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_274), .A2(n_402), .B1(n_403), .B2(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_277), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_277), .B(n_336), .Y(n_377) );
AND2x2_ASAP7_75t_L g424 ( .A(n_277), .B(n_309), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_278), .B(n_325), .Y(n_372) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g425 ( .A(n_280), .Y(n_425) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
INVx1_ASAP7_75t_L g350 ( .A(n_281), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_283), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g397 ( .A(n_283), .B(n_317), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_283), .B(n_312), .Y(n_404) );
INVx1_ASAP7_75t_SL g386 ( .A(n_285), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_286), .B(n_337), .Y(n_364) );
NOR4xp25_ASAP7_75t_L g410 ( .A(n_286), .B(n_309), .C(n_411), .D(n_414), .Y(n_410) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_287), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVxp67_ASAP7_75t_L g367 ( .A(n_290), .Y(n_367) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OAI21xp33_ASAP7_75t_L g417 ( .A1(n_293), .A2(n_384), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g309 ( .A(n_294), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g358 ( .A(n_297), .Y(n_358) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND4xp25_ASAP7_75t_SL g300 ( .A(n_301), .B(n_326), .C(n_341), .D(n_361), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_307), .B(n_311), .C(n_313), .Y(n_301) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g393 ( .A(n_306), .B(n_336), .Y(n_393) );
AND2x2_ASAP7_75t_L g402 ( .A(n_306), .B(n_380), .Y(n_402) );
INVx3_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_309), .B(n_344), .Y(n_406) );
AND2x2_ASAP7_75t_L g318 ( .A(n_312), .B(n_319), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_320), .B1(n_322), .B2(n_323), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
AND2x2_ASAP7_75t_L g416 ( .A(n_316), .B(n_362), .Y(n_416) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_318), .B(n_367), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_319), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_330), .B(n_332), .C(n_334), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_327), .A2(n_362), .B1(n_363), .B2(n_365), .C(n_368), .Y(n_361) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_335), .A2(n_420), .B1(n_423), .B2(n_425), .C(n_426), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_336), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_344), .B(n_413), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g374 ( .A(n_346), .Y(n_374) );
INVx1_ASAP7_75t_SL g348 ( .A(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_349), .A2(n_369), .B1(n_371), .B2(n_372), .Y(n_368) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AOI21xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B(n_359), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_358), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_369), .A2(n_395), .B1(n_433), .B2(n_434), .C(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
OAI211xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B(n_381), .C(n_401), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_385), .C(n_394), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
A2O1A1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g413 ( .A(n_391), .Y(n_413) );
OAI21xp5_ASAP7_75t_SL g435 ( .A1(n_392), .A2(n_418), .B(n_436), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_398), .Y(n_394) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVxp67_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g427 ( .A1(n_404), .A2(n_428), .B(n_429), .Y(n_427) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_419), .C(n_432), .Y(n_407) );
OAI211xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_415), .C(n_417), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
CKINVDCx14_ASAP7_75t_R g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
NOR2x2_ASAP7_75t_L g748 ( .A(n_448), .B(n_461), .Y(n_748) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_452), .B(n_456), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
XNOR2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_737), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR3x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_665), .C(n_714), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_580), .C(n_608), .D(n_638), .E(n_652), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_503), .B1(n_533), .B2(n_538), .C(n_547), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_480), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_467), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g560 ( .A(n_468), .Y(n_560) );
AND2x2_ASAP7_75t_L g568 ( .A(n_468), .B(n_483), .Y(n_568) );
AND2x2_ASAP7_75t_L g591 ( .A(n_468), .B(n_482), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_468), .B(n_493), .Y(n_606) );
OR2x2_ASAP7_75t_L g615 ( .A(n_468), .B(n_554), .Y(n_615) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_468), .Y(n_618) );
AND2x2_ASAP7_75t_L g726 ( .A(n_468), .B(n_554), .Y(n_726) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_473), .B(n_478), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_475), .A2(n_491), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_480), .B(n_618), .Y(n_674) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
OAI311xp33_ASAP7_75t_L g616 ( .A1(n_481), .A2(n_617), .A3(n_618), .B1(n_619), .C1(n_634), .Y(n_616) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .Y(n_481) );
AND2x2_ASAP7_75t_L g577 ( .A(n_482), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g584 ( .A(n_482), .Y(n_584) );
AND2x2_ASAP7_75t_L g705 ( .A(n_482), .B(n_537), .Y(n_705) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_483), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g561 ( .A(n_483), .B(n_493), .Y(n_561) );
AND2x2_ASAP7_75t_L g613 ( .A(n_483), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g627 ( .A(n_483), .B(n_560), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_491), .Y(n_488) );
INVx2_ASAP7_75t_L g537 ( .A(n_493), .Y(n_537) );
AND2x2_ASAP7_75t_L g576 ( .A(n_493), .B(n_560), .Y(n_576) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_511), .Y(n_503) );
OR2x2_ASAP7_75t_L g671 ( .A(n_504), .B(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_504), .B(n_677), .Y(n_688) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_505), .B(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g546 ( .A(n_506), .Y(n_546) );
AND2x2_ASAP7_75t_L g612 ( .A(n_506), .B(n_542), .Y(n_612) );
AND2x2_ASAP7_75t_L g623 ( .A(n_506), .B(n_523), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_506), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_511), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_511), .B(n_573), .Y(n_617) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g604 ( .A(n_512), .B(n_563), .Y(n_604) );
OR2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_523), .Y(n_512) );
INVx2_ASAP7_75t_L g540 ( .A(n_513), .Y(n_540) );
AND2x2_ASAP7_75t_L g631 ( .A(n_513), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g550 ( .A(n_514), .Y(n_550) );
OR2x2_ASAP7_75t_L g648 ( .A(n_514), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_514), .Y(n_711) );
AND2x2_ASAP7_75t_L g551 ( .A(n_523), .B(n_546), .Y(n_551) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
AND2x2_ASAP7_75t_L g592 ( .A(n_523), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g633 ( .A(n_523), .Y(n_633) );
INVx1_ASAP7_75t_L g649 ( .A(n_523), .Y(n_649) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_523), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .Y(n_525) );
INVxp67_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_535), .B(n_637), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_535), .A2(n_622), .B1(n_671), .B2(n_681), .Y(n_680) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
OAI211xp5_ASAP7_75t_SL g714 ( .A1(n_536), .A2(n_715), .B(n_717), .C(n_735), .Y(n_714) );
INVx2_ASAP7_75t_L g567 ( .A(n_537), .Y(n_567) );
AND2x2_ASAP7_75t_L g625 ( .A(n_537), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g636 ( .A(n_537), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_538), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
AND2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_573), .Y(n_609) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g641 ( .A(n_540), .B(n_632), .Y(n_641) );
AND2x2_ASAP7_75t_L g660 ( .A(n_540), .B(n_574), .Y(n_660) );
AND2x4_ASAP7_75t_L g596 ( .A(n_541), .B(n_570), .Y(n_596) );
AND2x2_ASAP7_75t_L g734 ( .A(n_541), .B(n_710), .Y(n_734) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_542), .Y(n_563) );
INVx1_ASAP7_75t_L g574 ( .A(n_542), .Y(n_574) );
INVx1_ASAP7_75t_L g673 ( .A(n_542), .Y(n_673) );
OR2x2_ASAP7_75t_L g564 ( .A(n_546), .B(n_550), .Y(n_564) );
AND2x2_ASAP7_75t_L g573 ( .A(n_546), .B(n_574), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g593 ( .A(n_546), .B(n_594), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_552), .B1(n_562), .B2(n_565), .C(n_569), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_549), .A2(n_570), .B(n_572), .C(n_575), .Y(n_569) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx1_ASAP7_75t_L g594 ( .A(n_550), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_550), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_SL g677 ( .A(n_550), .B(n_571), .Y(n_677) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_550), .Y(n_684) );
AND2x2_ASAP7_75t_L g602 ( .A(n_551), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g639 ( .A(n_551), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_561), .Y(n_552) );
INVx2_ASAP7_75t_L g630 ( .A(n_553), .Y(n_630) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_553), .A2(n_563), .B1(n_680), .B2(n_682), .C1(n_683), .C2(n_685), .Y(n_679) );
AND2x2_ASAP7_75t_L g736 ( .A(n_553), .B(n_705), .Y(n_736) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_560), .Y(n_553) );
INVx1_ASAP7_75t_L g626 ( .A(n_554), .Y(n_626) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g578 ( .A(n_559), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g664 ( .A(n_561), .B(n_598), .Y(n_664) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_562), .A2(n_676), .B(n_678), .Y(n_675) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx2_ASAP7_75t_L g603 ( .A(n_563), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_563), .B(n_570), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_563), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
INVx3_ASAP7_75t_L g629 ( .A(n_567), .Y(n_629) );
OR2x2_ASAP7_75t_L g681 ( .A(n_567), .B(n_603), .Y(n_681) );
AND2x2_ASAP7_75t_L g597 ( .A(n_568), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g635 ( .A(n_568), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_568), .B(n_629), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_568), .B(n_625), .Y(n_651) );
AND2x2_ASAP7_75t_L g655 ( .A(n_568), .B(n_637), .Y(n_655) );
INVxp67_ASAP7_75t_L g587 ( .A(n_570), .Y(n_587) );
BUFx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_572), .A2(n_645), .B1(n_650), .B2(n_651), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_572), .B(n_677), .Y(n_707) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g693 ( .A(n_573), .B(n_684), .Y(n_693) );
AND2x2_ASAP7_75t_L g722 ( .A(n_573), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g727 ( .A(n_573), .B(n_677), .Y(n_727) );
INVx1_ASAP7_75t_L g640 ( .A(n_574), .Y(n_640) );
BUFx2_ASAP7_75t_L g646 ( .A(n_574), .Y(n_646) );
INVx1_ASAP7_75t_L g731 ( .A(n_575), .Y(n_731) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g582 ( .A(n_576), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g607 ( .A(n_577), .Y(n_607) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_578), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g590 ( .A(n_578), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g599 ( .A(n_578), .Y(n_599) );
INVx3_ASAP7_75t_L g637 ( .A(n_578), .Y(n_637) );
OR2x2_ASAP7_75t_L g703 ( .A(n_578), .B(n_704), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_585), .B(n_588), .C(n_600), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g717 ( .A1(n_581), .A2(n_718), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_717) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_595), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_591), .B(n_629), .Y(n_643) );
AND2x2_ASAP7_75t_L g685 ( .A(n_591), .B(n_625), .Y(n_685) );
INVx1_ASAP7_75t_SL g698 ( .A(n_592), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_592), .B(n_646), .Y(n_701) );
INVx1_ASAP7_75t_L g719 ( .A(n_593), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_597), .A2(n_687), .B1(n_689), .B2(n_693), .C(n_694), .Y(n_686) );
AND2x2_ASAP7_75t_L g713 ( .A(n_598), .B(n_705), .Y(n_713) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g697 ( .A(n_599), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g600 ( .A1(n_601), .A2(n_604), .B(n_605), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g668 ( .A(n_603), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g654 ( .A(n_604), .Y(n_654) );
INVx1_ASAP7_75t_L g682 ( .A(n_605), .Y(n_682) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_613), .C(n_616), .Y(n_608) );
OAI31xp33_ASAP7_75t_L g735 ( .A1(n_609), .A2(n_647), .A3(n_734), .B(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g709 ( .A(n_612), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_SL g730 ( .A(n_612), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_614), .B(n_629), .Y(n_657) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g732 ( .A(n_615), .B(n_629), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_624), .B1(n_628), .B2(n_631), .Y(n_619) );
NAND2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_623), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g659 ( .A(n_623), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g662 ( .A(n_623), .B(n_646), .Y(n_662) );
AND2x2_ASAP7_75t_L g716 ( .A(n_623), .B(n_711), .Y(n_716) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g691 ( .A(n_627), .Y(n_691) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .Y(n_628) );
OAI32xp33_ASAP7_75t_L g694 ( .A1(n_629), .A2(n_663), .A3(n_695), .B1(n_697), .B2(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g669 ( .A(n_632), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_632), .B(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g692 ( .A(n_636), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B(n_642), .C(n_644), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_640), .B(n_677), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_641), .A2(n_653), .B1(n_654), .B2(n_655), .C(n_656), .Y(n_652) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g653 ( .A(n_651), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_661), .B2(n_663), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND4xp25_ASAP7_75t_SL g718 ( .A(n_661), .B(n_719), .C(n_720), .D(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g663 ( .A(n_664), .Y(n_663) );
NAND4xp25_ASAP7_75t_SL g665 ( .A(n_666), .B(n_679), .C(n_686), .D(n_699), .Y(n_665) );
O2A1O1Ixp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B(n_674), .C(n_675), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_SL g696 ( .A(n_672), .Y(n_696) );
INVx2_ASAP7_75t_L g720 ( .A(n_677), .Y(n_720) );
OR2x2_ASAP7_75t_L g729 ( .A(n_684), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_706), .Y(n_699) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g725 ( .A(n_705), .B(n_726), .Y(n_725) );
AOI21xp33_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_708), .B(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx3_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx5_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx9p33_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_752), .Y(n_760) );
OR2x4_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
endmodule