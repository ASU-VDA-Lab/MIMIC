module fake_jpeg_17803_n_329 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_21),
.Y(n_49)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_21),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_53),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_40),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_29),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_17),
.Y(n_86)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_88),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_38),
.B1(n_19),
.B2(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_72),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_19),
.B1(n_42),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_85),
.B1(n_82),
.B2(n_57),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_89),
.Y(n_100)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_19),
.B1(n_28),
.B2(n_24),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_37),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_24),
.B1(n_22),
.B2(n_32),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_43),
.B1(n_41),
.B2(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_37),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_27),
.B1(n_20),
.B2(n_18),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_76),
.B1(n_78),
.B2(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_99),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_60),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_69),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_51),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_117),
.B(n_33),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_50),
.B1(n_52),
.B2(n_63),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_76),
.B1(n_78),
.B2(n_43),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_58),
.C(n_43),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_113),
.C(n_104),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_70),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_121),
.B(n_101),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_95),
.A2(n_73),
.B1(n_84),
.B2(n_82),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_128),
.B1(n_131),
.B2(n_136),
.Y(n_151)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_143),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_134),
.C(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_140),
.C(n_132),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_89),
.Y(n_127)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_67),
.C(n_62),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_17),
.B1(n_25),
.B2(n_29),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_62),
.B1(n_13),
.B2(n_14),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_97),
.B1(n_100),
.B2(n_115),
.Y(n_159)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_114),
.B(n_0),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_99),
.B(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_97),
.B(n_86),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_34),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_125),
.A2(n_116),
.B1(n_117),
.B2(n_107),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_152),
.B(n_157),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_146),
.B(n_96),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_154),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_116),
.B1(n_117),
.B2(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_111),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_166),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_159),
.B(n_175),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_160),
.A2(n_162),
.B(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_119),
.B(n_106),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_163),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_129),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_93),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_174),
.C(n_131),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_109),
.B(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_103),
.Y(n_170)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_31),
.B(n_23),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_171),
.B(n_173),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_118),
.B1(n_98),
.B2(n_31),
.Y(n_172)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_33),
.B(n_34),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_34),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_177),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

INVx13_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_179),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_199),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_185),
.C(n_191),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_144),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_148),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_186),
.A2(n_177),
.B(n_157),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_149),
.B(n_153),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_192),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_121),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_135),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_194),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_142),
.C(n_139),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_174),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_160),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_203),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_157),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_209),
.A2(n_31),
.B1(n_30),
.B2(n_26),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_222),
.Y(n_242)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_213),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_230),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g243 ( 
.A1(n_216),
.A2(n_205),
.B(n_187),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_154),
.Y(n_218)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_124),
.B1(n_173),
.B2(n_142),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_219),
.A2(n_229),
.B1(n_193),
.B2(n_194),
.Y(n_235)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_225),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_139),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_227),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_232),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_183),
.A2(n_130),
.B1(n_129),
.B2(n_67),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_130),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_62),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_198),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_186),
.B1(n_200),
.B2(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_208),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_252),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_212),
.A2(n_227),
.B1(n_220),
.B2(n_226),
.Y(n_240)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_240),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_187),
.B1(n_204),
.B2(n_178),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_231),
.B(n_214),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_250),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

XNOR2x1_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_188),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g252 ( 
.A(n_209),
.B(n_185),
.CI(n_188),
.CON(n_252),
.SN(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_218),
.A2(n_182),
.B1(n_31),
.B2(n_30),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_219),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_213),
.A2(n_182),
.B1(n_2),
.B2(n_1),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_216),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_242),
.A2(n_224),
.B(n_211),
.Y(n_258)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_237),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_264),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_233),
.C(n_230),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_269),
.C(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_236),
.B(n_223),
.C(n_221),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_211),
.C(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_241),
.B(n_238),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_271),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_215),
.C(n_67),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_255),
.Y(n_282)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_268),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_234),
.Y(n_275)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_257),
.A2(n_251),
.B1(n_244),
.B2(n_239),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_249),
.Y(n_278)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_278),
.Y(n_294)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_243),
.B(n_248),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_259),
.A2(n_246),
.B1(n_254),
.B2(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_9),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_284),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_L g286 ( 
.A1(n_261),
.A2(n_30),
.A3(n_26),
.B1(n_23),
.B2(n_16),
.C1(n_6),
.C2(n_7),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g299 ( 
.A(n_286),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_10),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_287),
.B(n_13),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_298),
.C(n_299),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_283),
.A2(n_256),
.B(n_269),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_295),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_262),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_298),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_267),
.B(n_266),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_281),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_262),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_277),
.B(n_274),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_304),
.B(n_306),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_273),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_280),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_285),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_307),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_290),
.B1(n_292),
.B2(n_276),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_30),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_308),
.A2(n_310),
.B1(n_26),
.B2(n_23),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_26),
.B1(n_23),
.B2(n_16),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_315),
.C(n_302),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_309),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_16),
.C(n_5),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_319),
.B1(n_321),
.B2(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_R g319 ( 
.A(n_317),
.B(n_312),
.C(n_311),
.Y(n_319)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_320),
.A2(n_13),
.B(n_5),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_323),
.B(n_8),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_325),
.A2(n_12),
.B1(n_8),
.B2(n_9),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_10),
.C(n_12),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_2),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_2),
.B(n_323),
.Y(n_329)
);


endmodule