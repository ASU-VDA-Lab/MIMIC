module fake_jpeg_2320_n_569 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_569);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_569;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVxp33_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_57),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_30),
.B(n_8),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_58),
.B(n_75),
.Y(n_131)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_35),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_84),
.Y(n_113)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_66),
.Y(n_115)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_8),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_77),
.Y(n_165)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_80),
.Y(n_175)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_36),
.B(n_37),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_89),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_22),
.B(n_8),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_87),
.Y(n_163)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_37),
.B(n_9),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_7),
.B(n_1),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_91),
.C(n_22),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_28),
.B(n_7),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_93),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_95),
.Y(n_173)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_96),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_44),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_23),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_28),
.Y(n_98)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_28),
.Y(n_100)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_100),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_101),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_103),
.Y(n_176)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_40),
.Y(n_107)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_54),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_40),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_112),
.B(n_48),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_52),
.B1(n_18),
.B2(n_53),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_114),
.A2(n_116),
.B1(n_130),
.B2(n_145),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_45),
.B1(n_40),
.B2(n_48),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_74),
.A2(n_18),
.B1(n_53),
.B2(n_51),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_48),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_134),
.B(n_135),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_98),
.B(n_48),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_39),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_136),
.B(n_148),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_141),
.B(n_144),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_78),
.B(n_46),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_80),
.A2(n_33),
.B1(n_38),
.B2(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_68),
.B(n_39),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_46),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_153),
.B(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_73),
.B(n_48),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_77),
.A2(n_45),
.B1(n_23),
.B2(n_34),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_63),
.B1(n_41),
.B2(n_29),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_43),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_56),
.B(n_29),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_43),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_166),
.B(n_40),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_67),
.A2(n_45),
.B1(n_48),
.B2(n_40),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_169),
.A2(n_63),
.B1(n_96),
.B2(n_92),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_111),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_179),
.B(n_231),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_180),
.A2(n_186),
.B1(n_211),
.B2(n_221),
.Y(n_266)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g299 ( 
.A(n_181),
.Y(n_299)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_176),
.Y(n_182)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_182),
.Y(n_263)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_125),
.Y(n_183)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_183),
.Y(n_296)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_184),
.Y(n_245)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_161),
.A2(n_95),
.B1(n_102),
.B2(n_101),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_146),
.Y(n_187)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_187),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_113),
.A2(n_76),
.B1(n_79),
.B2(n_86),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_188),
.A2(n_229),
.B(n_12),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_189),
.A2(n_225),
.B1(n_230),
.B2(n_240),
.Y(n_287)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_120),
.Y(n_191)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_193),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_114),
.A2(n_41),
.B1(n_99),
.B2(n_82),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_194),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_303)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_195),
.Y(n_272)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_196),
.Y(n_290)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

OA22x2_ASAP7_75t_SL g200 ( 
.A1(n_134),
.A2(n_54),
.B1(n_109),
.B2(n_59),
.Y(n_200)
);

OA22x2_ASAP7_75t_SL g286 ( 
.A1(n_200),
.A2(n_47),
.B1(n_4),
.B2(n_5),
.Y(n_286)
);

AOI21xp33_ASAP7_75t_L g258 ( 
.A1(n_202),
.A2(n_238),
.B(n_239),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_203),
.Y(n_253)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_204),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_110),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_205),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_126),
.A2(n_25),
.B1(n_53),
.B2(n_51),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_126),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_208),
.B(n_212),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_126),
.A2(n_31),
.B1(n_51),
.B2(n_25),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_209),
.Y(n_283)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_117),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_138),
.A2(n_25),
.B1(n_32),
.B2(n_31),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g212 ( 
.A(n_143),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_150),
.B(n_87),
.C(n_31),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_214),
.B(n_223),
.C(n_196),
.Y(n_268)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_152),
.Y(n_217)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_123),
.Y(n_218)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_218),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_220),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_168),
.A2(n_32),
.B1(n_94),
.B2(n_47),
.Y(n_221)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

INVx11_ASAP7_75t_SL g278 ( 
.A(n_222),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_159),
.Y(n_223)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_223),
.Y(n_281)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_158),
.Y(n_224)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_224),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_115),
.A2(n_32),
.B1(n_40),
.B2(n_94),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_110),
.Y(n_228)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g229 ( 
.A(n_154),
.B(n_0),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_123),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_116),
.A2(n_38),
.B1(n_33),
.B2(n_47),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_137),
.B1(n_165),
.B2(n_178),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_140),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_242),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_236),
.Y(n_274)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_121),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_124),
.Y(n_239)
);

INVx4_ASAP7_75t_SL g240 ( 
.A(n_172),
.Y(n_240)
);

AND2x4_ASAP7_75t_L g241 ( 
.A(n_127),
.B(n_38),
.Y(n_241)
);

OR2x4_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_54),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_132),
.B(n_0),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_158),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_243),
.A2(n_4),
.B1(n_12),
.B2(n_14),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_244),
.A2(n_254),
.B1(n_255),
.B2(n_261),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_193),
.A2(n_131),
.B1(n_163),
.B2(n_170),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_247),
.A2(n_187),
.B(n_210),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_207),
.A2(n_175),
.B1(n_165),
.B2(n_139),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_175),
.B1(n_151),
.B2(n_157),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_177),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_260),
.B(n_277),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_186),
.A2(n_177),
.B1(n_170),
.B2(n_169),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_173),
.B1(n_133),
.B2(n_47),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_262),
.A2(n_271),
.B1(n_294),
.B2(n_244),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_268),
.B(n_277),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_229),
.A2(n_174),
.B(n_54),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_270),
.A2(n_276),
.B(n_300),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_180),
.A2(n_173),
.B1(n_133),
.B2(n_47),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_208),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_202),
.B(n_33),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_216),
.A2(n_174),
.B1(n_47),
.B2(n_50),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_279),
.A2(n_282),
.B1(n_289),
.B2(n_303),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_188),
.A2(n_242),
.B1(n_215),
.B2(n_201),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_214),
.B(n_0),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_284),
.B(n_288),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_235),
.B(n_1),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_212),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_15),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_2),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_200),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_241),
.A2(n_4),
.B1(n_6),
.B2(n_10),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_200),
.B(n_184),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_305),
.A2(n_321),
.B(n_324),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_306),
.B(n_308),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_246),
.A2(n_221),
.B1(n_241),
.B2(n_185),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_318),
.B1(n_319),
.B2(n_328),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_354),
.C(n_314),
.Y(n_385)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_311),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_312),
.B(n_322),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_278),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_254),
.A2(n_191),
.B1(n_236),
.B2(n_226),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_246),
.A2(n_182),
.B1(n_204),
.B2(n_195),
.Y(n_319)
);

AO21x2_ASAP7_75t_SL g320 ( 
.A1(n_286),
.A2(n_222),
.B(n_240),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_320),
.A2(n_252),
.B1(n_292),
.B2(n_314),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_270),
.A2(n_187),
.B(n_198),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_269),
.B(n_197),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_284),
.B(n_192),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_323),
.B(n_329),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_230),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_326),
.Y(n_361)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_327),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_262),
.A2(n_181),
.B1(n_218),
.B2(n_183),
.Y(n_328)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_295),
.Y(n_331)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_331),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_266),
.A2(n_224),
.B1(n_243),
.B2(n_205),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_332),
.A2(n_349),
.B1(n_292),
.B2(n_273),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_264),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_245),
.Y(n_334)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_334),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_190),
.Y(n_336)
);

INVxp33_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_228),
.Y(n_337)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_253),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_341),
.Y(n_357)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_245),
.Y(n_339)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_339),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_265),
.A2(n_17),
.B(n_15),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_344),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_257),
.B(n_15),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_272),
.Y(n_343)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_265),
.A2(n_16),
.B(n_283),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_268),
.B(n_16),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_346),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_290),
.B(n_247),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_289),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_347),
.B(n_353),
.Y(n_387)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_263),
.Y(n_348)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_348),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_290),
.A2(n_16),
.B1(n_283),
.B2(n_286),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_287),
.A2(n_16),
.B(n_302),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_329),
.Y(n_386)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_352),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_253),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_249),
.B(n_250),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_347),
.A2(n_255),
.B1(n_294),
.B2(n_274),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_363),
.A2(n_365),
.B1(n_369),
.B2(n_372),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_325),
.A2(n_302),
.B1(n_297),
.B2(n_273),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_364),
.A2(n_368),
.B(n_381),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_346),
.A2(n_297),
.B1(n_259),
.B2(n_301),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_310),
.A2(n_248),
.B1(n_301),
.B2(n_280),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_310),
.A2(n_248),
.B1(n_293),
.B2(n_251),
.Y(n_372)
);

OAI22xp33_ASAP7_75t_SL g373 ( 
.A1(n_320),
.A2(n_259),
.B1(n_296),
.B2(n_291),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_373),
.A2(n_320),
.B1(n_377),
.B2(n_328),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_308),
.A2(n_272),
.B1(n_275),
.B2(n_291),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_384),
.B1(n_318),
.B2(n_330),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_304),
.A2(n_256),
.B1(n_275),
.B2(n_296),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_379),
.A2(n_333),
.B1(n_334),
.B2(n_339),
.Y(n_405)
);

OAI22x1_ASAP7_75t_SL g384 ( 
.A1(n_320),
.A2(n_252),
.B1(n_305),
.B2(n_344),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_385),
.B(n_354),
.C(n_311),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_323),
.B(n_336),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_394),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_322),
.Y(n_391)
);

CKINVDCx14_ASAP7_75t_R g410 ( 
.A(n_391),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_342),
.B(n_309),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_337),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_396),
.B(n_331),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_397),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_338),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_400),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_394),
.B(n_385),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_403),
.C(n_413),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_389),
.B(n_342),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_375),
.B(n_345),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_402),
.B(n_362),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_405),
.A2(n_363),
.B1(n_369),
.B2(n_380),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_406),
.B(n_427),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_320),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_319),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_408),
.B(n_415),
.Y(n_442)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_411),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_417),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_355),
.B(n_321),
.C(n_324),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_393),
.A2(n_350),
.B1(n_329),
.B2(n_304),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_422),
.B1(n_386),
.B2(n_387),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_L g415 ( 
.A1(n_375),
.A2(n_315),
.B(n_312),
.Y(n_415)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_384),
.B(n_329),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_416),
.Y(n_439)
);

OAI21xp33_ASAP7_75t_L g417 ( 
.A1(n_360),
.A2(n_349),
.B(n_324),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_371),
.B(n_337),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_424),
.C(n_425),
.Y(n_444)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_361),
.Y(n_419)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_357),
.B(n_316),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_428),
.Y(n_435)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_393),
.A2(n_306),
.B1(n_307),
.B2(n_332),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_355),
.B(n_317),
.C(n_326),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_366),
.B(n_343),
.C(n_351),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_388),
.A2(n_313),
.B(n_340),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_426),
.A2(n_430),
.B(n_367),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_390),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_372),
.B(n_327),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_433),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_388),
.A2(n_348),
.B(n_352),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_366),
.B(n_371),
.C(n_360),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_378),
.C(n_383),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_368),
.B(n_378),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_441),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_398),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_416),
.A2(n_359),
.B1(n_365),
.B2(n_379),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_443),
.B(n_445),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_410),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_446),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_448),
.B(n_402),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_356),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_449),
.B(n_450),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_362),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_463),
.C(n_404),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_424),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_452),
.B(n_453),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_405),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_416),
.A2(n_359),
.B1(n_364),
.B2(n_367),
.Y(n_454)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_455),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_408),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_456),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_414),
.A2(n_376),
.B1(n_380),
.B2(n_382),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_460),
.A2(n_412),
.B(n_430),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_429),
.A2(n_376),
.B1(n_382),
.B2(n_358),
.Y(n_461)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_423),
.A2(n_392),
.B1(n_390),
.B2(n_395),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_423),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_404),
.B(n_395),
.C(n_392),
.Y(n_463)
);

XOR2x2_ASAP7_75t_L g466 ( 
.A(n_449),
.B(n_432),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_466),
.B(n_488),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_436),
.B(n_450),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_469),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_437),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_418),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_471),
.B(n_440),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_472),
.B(n_474),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_448),
.B(n_409),
.Y(n_474)
);

NAND3xp33_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_400),
.C(n_431),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_475),
.A2(n_439),
.B1(n_435),
.B2(n_447),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_413),
.C(n_431),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_479),
.C(n_481),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_425),
.C(n_409),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_433),
.C(n_422),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_483),
.A2(n_443),
.B1(n_459),
.B2(n_461),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_433),
.C(n_407),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_486),
.C(n_487),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_407),
.C(n_411),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_446),
.B(n_419),
.C(n_401),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_434),
.B(n_426),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_401),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_437),
.Y(n_511)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_491),
.Y(n_519)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_473),
.Y(n_495)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_495),
.Y(n_520)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_486),
.Y(n_496)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_468),
.B(n_464),
.C(n_447),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_498),
.B(n_499),
.Y(n_527)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_476),
.Y(n_499)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_484),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_501),
.A2(n_504),
.B1(n_508),
.B2(n_509),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_506),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_511),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_464),
.C(n_454),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_507),
.C(n_469),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_489),
.A2(n_460),
.B(n_459),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_482),
.B(n_437),
.C(n_459),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_467),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_510),
.B(n_483),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_482),
.B(n_455),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_512),
.B(n_481),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_515),
.B(n_518),
.Y(n_534)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_507),
.A2(n_465),
.B(n_487),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_516),
.A2(n_421),
.B1(n_514),
.B2(n_515),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_517),
.B(n_529),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_505),
.A2(n_480),
.B1(n_456),
.B2(n_462),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_521),
.A2(n_528),
.B1(n_493),
.B2(n_500),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_522),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_479),
.C(n_466),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_526),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_478),
.C(n_488),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_512),
.A2(n_438),
.B1(n_457),
.B2(n_428),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_498),
.B(n_472),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_527),
.B(n_492),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_531),
.B(n_519),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_513),
.A2(n_439),
.B1(n_503),
.B2(n_511),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_532),
.A2(n_540),
.B1(n_534),
.B2(n_536),
.Y(n_551)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_533),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_493),
.C(n_500),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_535),
.B(n_540),
.C(n_543),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_525),
.A2(n_438),
.B(n_457),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_536),
.A2(n_537),
.B(n_532),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_458),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_523),
.A2(n_494),
.B1(n_458),
.B2(n_474),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_538),
.B(n_542),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_494),
.C(n_427),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_518),
.B(n_516),
.C(n_526),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_516),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_551),
.Y(n_557)
);

NOR2x1_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_538),
.Y(n_547)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_547),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_549),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_539),
.B(n_514),
.C(n_529),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_520),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_553),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_545),
.B(n_535),
.C(n_541),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_559),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_544),
.C(n_546),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_554),
.B(n_549),
.Y(n_560)
);

AO21x1_ASAP7_75t_L g564 ( 
.A1(n_560),
.A2(n_561),
.B(n_551),
.Y(n_564)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_555),
.Y(n_561)
);

NAND2x1_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_556),
.Y(n_563)
);

AO21x1_ASAP7_75t_L g565 ( 
.A1(n_563),
.A2(n_564),
.B(n_557),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_565),
.B(n_558),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_566),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_550),
.C(n_547),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_550),
.Y(n_569)
);


endmodule