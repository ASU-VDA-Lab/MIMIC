module fake_jpeg_15730_n_315 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_33),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_43),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_31),
.B1(n_20),
.B2(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_60),
.B1(n_63),
.B2(n_19),
.Y(n_72)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_26),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_51),
.B(n_54),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_38),
.B(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_16),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_31),
.B1(n_20),
.B2(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_31),
.B1(n_33),
.B2(n_19),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_67),
.Y(n_99)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_43),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_19),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_68),
.A2(n_76),
.B1(n_79),
.B2(n_83),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_72),
.A2(n_102),
.B1(n_90),
.B2(n_82),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_40),
.B1(n_44),
.B2(n_39),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_74),
.A2(n_75),
.B1(n_57),
.B2(n_49),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_46),
.A2(n_42),
.B1(n_40),
.B2(n_43),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_95),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_26),
.B1(n_32),
.B2(n_22),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_88),
.B1(n_93),
.B2(n_97),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_48),
.B(n_0),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_33),
.B1(n_42),
.B2(n_16),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_47),
.B(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_85),
.B(n_28),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_29),
.B1(n_27),
.B2(n_32),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_100),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_48),
.A2(n_29),
.B1(n_40),
.B2(n_18),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_44),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_55),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_25),
.B1(n_18),
.B2(n_24),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_113),
.B(n_121),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_115),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_101),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_119),
.B1(n_96),
.B2(n_98),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_72),
.C(n_86),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_79),
.C(n_21),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_128),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_68),
.B(n_18),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_57),
.B1(n_44),
.B2(n_39),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_122),
.A2(n_91),
.B1(n_74),
.B2(n_94),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_68),
.B(n_21),
.CI(n_30),
.CON(n_123),
.SN(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_130),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_89),
.B(n_62),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_124),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_13),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_44),
.Y(n_130)
);

OAI22x1_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_104),
.B1(n_111),
.B2(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_132),
.A2(n_148),
.B1(n_113),
.B2(n_122),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_76),
.B(n_79),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_135),
.A2(n_141),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_137),
.B(n_155),
.Y(n_170)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_125),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_130),
.B(n_108),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_123),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_96),
.B1(n_98),
.B2(n_92),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_143),
.A2(n_145),
.B1(n_156),
.B2(n_128),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_107),
.B(n_87),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_157),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_74),
.B(n_21),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_74),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_115),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_158),
.B(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_114),
.B(n_71),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_44),
.B1(n_39),
.B2(n_25),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_30),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_30),
.B(n_1),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_110),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_162),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_169),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_164),
.A2(n_174),
.B1(n_178),
.B2(n_189),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_123),
.B(n_129),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_175),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_195),
.C(n_182),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_147),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_120),
.B(n_105),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_135),
.B(n_157),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_21),
.C(n_30),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_28),
.C(n_13),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_154),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_39),
.Y(n_186)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_132),
.A2(n_150),
.B1(n_131),
.B2(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_188),
.A2(n_191),
.B1(n_12),
.B2(n_14),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_136),
.A2(n_103),
.B1(n_125),
.B2(n_11),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_146),
.A2(n_11),
.B1(n_15),
.B2(n_14),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_194),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_125),
.Y(n_193)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_147),
.B(n_10),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_171),
.A2(n_133),
.B1(n_148),
.B2(n_134),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_196),
.A2(n_198),
.B1(n_204),
.B2(n_183),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_133),
.B1(n_134),
.B2(n_142),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_208),
.B(n_209),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_217),
.C(n_220),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_140),
.B1(n_158),
.B2(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_165),
.A2(n_153),
.B1(n_160),
.B2(n_12),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_0),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_165),
.B(n_1),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_210),
.A2(n_170),
.B(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_185),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_214),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_160),
.C(n_103),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_94),
.C(n_69),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_175),
.C(n_179),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_178),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_179),
.B(n_1),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_180),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_204),
.C(n_196),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_192),
.Y(n_224)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_224),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_197),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_226),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_227),
.B(n_228),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_219),
.B(n_172),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_242),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_235),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_236),
.A2(n_237),
.B1(n_202),
.B2(n_212),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_213),
.A2(n_164),
.B(n_191),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_241),
.Y(n_256)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_186),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_211),
.C(n_199),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_240),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_217),
.C(n_198),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_249),
.C(n_254),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_252),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_211),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_209),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_212),
.C(n_234),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_229),
.B(n_206),
.C(n_176),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_215),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_230),
.B(n_209),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_222),
.C(n_244),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_216),
.Y(n_262)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_262),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_272),
.B(n_273),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_243),
.B1(n_232),
.B2(n_240),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_208),
.B1(n_231),
.B2(n_236),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_275),
.C(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_247),
.B(n_226),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_231),
.B(n_224),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_253),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_261),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_288),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_253),
.C(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_281),
.C(n_285),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_241),
.B1(n_245),
.B2(n_270),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_280),
.A2(n_210),
.B1(n_2),
.B2(n_3),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_271),
.C(n_268),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_286),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_190),
.C(n_168),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_267),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_283),
.A2(n_168),
.B1(n_190),
.B2(n_210),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_296),
.B1(n_297),
.B2(n_10),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_2),
.Y(n_303)
);

OR2x2_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_8),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_2),
.B(n_3),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_8),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_69),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

AOI31xp33_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_281),
.A3(n_277),
.B(n_279),
.Y(n_299)
);

OAI22x1_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_302),
.B1(n_303),
.B2(n_304),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_1),
.C(n_2),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_295),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_6),
.B(n_7),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_289),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g310 ( 
.A(n_305),
.Y(n_310)
);

AOI21xp33_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_300),
.B(n_303),
.Y(n_309)
);

AOI321xp33_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_306),
.A3(n_308),
.B1(n_292),
.B2(n_293),
.C(n_13),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_311),
.B(n_7),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_310),
.C(n_14),
.Y(n_313)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_313),
.B(n_292),
.CI(n_10),
.CON(n_314),
.SN(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_307),
.Y(n_315)
);


endmodule