module fake_netlist_5_1158_n_2416 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_226, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2416);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2416;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_2323;
wire n_2203;
wire n_1243;
wire n_1016;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2249;
wire n_2180;
wire n_344;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_1070;
wire n_777;
wire n_422;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_283;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_1079;
wire n_457;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2339;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_2346;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_2400;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1928;
wire n_1848;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2282;
wire n_2002;
wire n_510;
wire n_2371;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1726;
wire n_665;
wire n_1584;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_791;
wire n_732;
wire n_1533;
wire n_1979;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2363;
wire n_916;
wire n_1081;
wire n_493;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_703;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_2375;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_1337;
wire n_420;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_2414;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2044;
wire n_1990;
wire n_2013;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_1),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_37),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_13),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_73),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_80),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_30),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_75),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_31),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_60),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_99),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_166),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_30),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_32),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_37),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_20),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_170),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_70),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_195),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g253 ( 
.A(n_15),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_155),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_181),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_79),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_189),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_58),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_19),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_105),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_190),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_7),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_109),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_6),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_51),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_192),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_17),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_148),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_36),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_111),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_88),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_66),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_32),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_176),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_122),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_88),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_143),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_70),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_18),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_210),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_114),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_27),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_102),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_156),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_215),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_41),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_56),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_97),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_121),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_89),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_59),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_199),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_175),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_232),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_219),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_19),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_12),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_207),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_177),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_49),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_130),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_194),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_126),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g309 ( 
.A(n_7),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_72),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_107),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_91),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_200),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_11),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_36),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_94),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_163),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_80),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_179),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_96),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_108),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_119),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_231),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_69),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_62),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_168),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_188),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_118),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_134),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_42),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_193),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_49),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_120),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_38),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_167),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_89),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_53),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_214),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_56),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_185),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_137),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_161),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_196),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_90),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_1),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_68),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_213),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_145),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_151),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_95),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_123),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_50),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_160),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_136),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_153),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_55),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_184),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_94),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_50),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_165),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_191),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_142),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_46),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_203),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_201),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_112),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_131),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_162),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_85),
.Y(n_369)
);

INVx2_ASAP7_75t_SL g370 ( 
.A(n_125),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_33),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_221),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_72),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_204),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_67),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_228),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_227),
.Y(n_377)
);

BUFx2_ASAP7_75t_SL g378 ( 
.A(n_73),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_22),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_86),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_31),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_25),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_93),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_86),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_67),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_171),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_182),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_85),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_68),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_35),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_97),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_217),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_229),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_38),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_140),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_0),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_183),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_60),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_139),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_225),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_144),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_39),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_216),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_45),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_41),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_150),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_169),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_146),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_39),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_71),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_100),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_79),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_14),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_81),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_82),
.Y(n_415)
);

BUFx10_ASAP7_75t_L g416 ( 
.A(n_132),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_222),
.Y(n_417)
);

BUFx10_ASAP7_75t_L g418 ( 
.A(n_54),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_4),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_17),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_3),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_2),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_157),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_84),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_103),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_54),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_22),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_40),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_53),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_128),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_45),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_25),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_75),
.Y(n_434)
);

BUFx10_ASAP7_75t_L g435 ( 
.A(n_104),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_26),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_226),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_99),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_62),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_63),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_57),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_48),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_173),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_174),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_35),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_78),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_5),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_113),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_133),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_66),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_28),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_106),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_211),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_21),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_149),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_34),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_91),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_255),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_243),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_286),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_252),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_254),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_256),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_379),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_263),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_379),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_296),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_367),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_379),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_271),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_273),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_260),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_277),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_253),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_260),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_266),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_253),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_260),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_260),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_278),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_283),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_287),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_260),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_374),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_260),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_419),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_288),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_289),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_298),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_258),
.B(n_0),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_308),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_302),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_291),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_308),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_305),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_338),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_436),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_338),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_291),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_436),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_436),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_311),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_436),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_313),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_317),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_321),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_245),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_327),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_328),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_245),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_329),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_331),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_245),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_261),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_350),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_258),
.B(n_2),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_306),
.B(n_326),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_261),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_335),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_261),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_341),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_280),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_375),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_375),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_342),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_293),
.B(n_4),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_267),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_343),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_350),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_348),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_280),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_349),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_351),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_353),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_354),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_234),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_355),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_267),
.Y(n_547)
);

INVxp67_ASAP7_75t_SL g548 ( 
.A(n_280),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_267),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_272),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_361),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_272),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_362),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_272),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_266),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_364),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_365),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_366),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_368),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_404),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_404),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_376),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_334),
.B(n_5),
.Y(n_563)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_386),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_316),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_316),
.Y(n_566)
);

NOR2xp67_ASAP7_75t_L g567 ( 
.A(n_334),
.B(n_6),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_378),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_387),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_399),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_316),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_403),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_433),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_345),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_345),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_406),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_266),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_345),
.Y(n_578)
);

NOR2xp67_ASAP7_75t_L g579 ( 
.A(n_334),
.B(n_8),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_408),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_346),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_479),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_525),
.B(n_535),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_482),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_482),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_459),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_461),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_499),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_465),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_485),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_460),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_458),
.B(n_293),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_462),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_485),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_465),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_531),
.B(n_347),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_463),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_465),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_486),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_466),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_526),
.B(n_284),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_548),
.B(n_377),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_490),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_469),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_540),
.B(n_377),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_477),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_492),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_520),
.B(n_417),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_492),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_495),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_478),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_495),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_505),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_540),
.B(n_347),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_474),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_491),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_540),
.B(n_377),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_505),
.B(n_395),
.Y(n_622)
);

AND2x2_ASAP7_75t_SL g623 ( 
.A(n_498),
.B(n_357),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_508),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_480),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_508),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_502),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_487),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_509),
.B(n_370),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_488),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_483),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_483),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

OA21x2_ASAP7_75t_L g634 ( 
.A1(n_483),
.A2(n_352),
.B(n_346),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_489),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_511),
.B(n_395),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_511),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_513),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_513),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_521),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_555),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_555),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_555),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_577),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_577),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_458),
.B(n_370),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_577),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_494),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_464),
.B(n_401),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_524),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_496),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_504),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_560),
.B(n_433),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_497),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_464),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_467),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_467),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_468),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_468),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_500),
.Y(n_660)
);

BUFx6f_ASAP7_75t_SL g661 ( 
.A(n_470),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_395),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_503),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_470),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_510),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_472),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_472),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

INVx2_ASAP7_75t_SL g669 ( 
.A(n_563),
.Y(n_669)
);

AND2x6_ASAP7_75t_L g670 ( 
.A(n_473),
.B(n_400),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_473),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_512),
.Y(n_672)
);

INVx1_ASAP7_75t_SL g673 ( 
.A(n_538),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_475),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_475),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_476),
.B(n_567),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_R g677 ( 
.A(n_514),
.B(n_426),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_528),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_666),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_634),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_666),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_666),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_656),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_656),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_604),
.B(n_515),
.Y(n_685)
);

OR2x2_ASAP7_75t_SL g686 ( 
.A(n_585),
.B(n_560),
.Y(n_686)
);

OR2x2_ASAP7_75t_SL g687 ( 
.A(n_585),
.B(n_532),
.Y(n_687)
);

OR2x2_ASAP7_75t_SL g688 ( 
.A(n_598),
.B(n_533),
.Y(n_688)
);

INVx6_ASAP7_75t_L g689 ( 
.A(n_636),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_636),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_669),
.B(n_517),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_591),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_673),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_604),
.B(n_518),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_601),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_669),
.B(n_537),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_609),
.B(n_357),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_670),
.Y(n_699)
);

INVx6_ASAP7_75t_L g700 ( 
.A(n_636),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_670),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_673),
.B(n_539),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_601),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_634),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_609),
.B(n_357),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_609),
.B(n_443),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_591),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_634),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_657),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_650),
.B(n_538),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_669),
.B(n_543),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_591),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_623),
.B(n_546),
.Y(n_713)
);

INVx4_ASAP7_75t_SL g714 ( 
.A(n_670),
.Y(n_714)
);

OR2x6_ASAP7_75t_L g715 ( 
.A(n_650),
.B(n_378),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_636),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_621),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_621),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_634),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_677),
.B(n_551),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_634),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_657),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_591),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_623),
.B(n_556),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_658),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_612),
.Y(n_726)
);

AO21x2_ASAP7_75t_L g727 ( 
.A1(n_676),
.A2(n_649),
.B(n_646),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_605),
.B(n_516),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_658),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_659),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_621),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_622),
.B(n_662),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_622),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_659),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_667),
.Y(n_735)
);

AND2x6_ASAP7_75t_L g736 ( 
.A(n_605),
.B(n_443),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_677),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_622),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_667),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_671),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_653),
.B(n_563),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_597),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_671),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_623),
.B(n_443),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_605),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_593),
.B(n_557),
.Y(n_746)
);

INVx5_ASAP7_75t_L g747 ( 
.A(n_670),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_676),
.B(n_558),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_662),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_597),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_590),
.Y(n_751)
);

OR2x2_ASAP7_75t_L g752 ( 
.A(n_598),
.B(n_561),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_618),
.B(n_570),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_655),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_662),
.B(n_400),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_618),
.B(n_297),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_655),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_655),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_595),
.B(n_572),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_588),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_597),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_584),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_597),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_606),
.Y(n_764)
);

INVxp33_ASAP7_75t_L g765 ( 
.A(n_590),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_582),
.B(n_519),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_580),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_603),
.B(n_530),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_608),
.B(n_534),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_606),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_582),
.B(n_519),
.Y(n_771)
);

NOR2xp67_ASAP7_75t_L g772 ( 
.A(n_610),
.B(n_568),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_664),
.B(n_471),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_664),
.B(n_400),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_664),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_674),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_594),
.B(n_297),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_615),
.A2(n_493),
.B(n_545),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_594),
.B(n_522),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_606),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_674),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_627),
.B(n_567),
.Y(n_782)
);

NAND2x1p5_ASAP7_75t_L g783 ( 
.A(n_674),
.B(n_284),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_644),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_675),
.B(n_476),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_646),
.B(n_573),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_625),
.B(n_541),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_632),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_583),
.B(n_522),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_670),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_640),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_583),
.B(n_523),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_644),
.Y(n_793)
);

AND2x2_ASAP7_75t_SL g794 ( 
.A(n_649),
.B(n_247),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_675),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_589),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_632),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_675),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_586),
.B(n_523),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_619),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_586),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_587),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_629),
.B(n_400),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_587),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_620),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_592),
.B(n_401),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_592),
.B(n_527),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_628),
.A2(n_542),
.B1(n_553),
.B2(n_544),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_L g810 ( 
.A(n_670),
.B(n_400),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_652),
.B(n_507),
.Y(n_811)
);

BUFx4f_ASAP7_75t_L g812 ( 
.A(n_670),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_596),
.Y(n_813)
);

AND2x2_ASAP7_75t_SL g814 ( 
.A(n_652),
.B(n_247),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_596),
.B(n_527),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_600),
.B(n_529),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_632),
.Y(n_817)
);

NOR2x1p5_ASAP7_75t_L g818 ( 
.A(n_630),
.B(n_275),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_644),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_668),
.B(n_507),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_647),
.Y(n_821)
);

BUFx4f_ASAP7_75t_L g822 ( 
.A(n_670),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_632),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_600),
.B(n_319),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_647),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_647),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_635),
.B(n_648),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_602),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_632),
.Y(n_829)
);

BUFx6f_ASAP7_75t_L g830 ( 
.A(n_632),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_602),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_629),
.B(n_400),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_651),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_632),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_607),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_607),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_611),
.B(n_529),
.Y(n_837)
);

NAND3xp33_ASAP7_75t_L g838 ( 
.A(n_654),
.B(n_481),
.C(n_484),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_611),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_613),
.B(n_319),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_724),
.A2(n_562),
.B1(n_564),
.B2(n_559),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_722),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_685),
.B(n_660),
.Y(n_843)
);

INVx2_ASAP7_75t_SL g844 ( 
.A(n_694),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_SL g845 ( 
.A(n_726),
.B(n_663),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_762),
.A2(n_576),
.B1(n_569),
.B2(n_661),
.Y(n_846)
);

INVx2_ASAP7_75t_SL g847 ( 
.A(n_694),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_713),
.B(n_762),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_680),
.A2(n_670),
.B(n_614),
.Y(n_849)
);

O2A1O1Ixp5_ASAP7_75t_L g850 ( 
.A1(n_680),
.A2(n_614),
.B(n_616),
.C(n_613),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_744),
.A2(n_661),
.B1(n_672),
.B2(n_665),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_732),
.B(n_616),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_744),
.A2(n_579),
.B(n_259),
.C(n_262),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_794),
.A2(n_352),
.B1(n_383),
.B2(n_346),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_741),
.A2(n_661),
.B1(n_437),
.B2(n_444),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_710),
.Y(n_856)
);

AND2x6_ASAP7_75t_SL g857 ( 
.A(n_787),
.B(n_234),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_717),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_710),
.B(n_745),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_722),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_711),
.B(n_437),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_691),
.B(n_501),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_717),
.Y(n_863)
);

AND2x6_ASAP7_75t_SL g864 ( 
.A(n_746),
.B(n_238),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_833),
.B(n_668),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_697),
.B(n_745),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_690),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_732),
.B(n_431),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_732),
.B(n_448),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_725),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_733),
.B(n_617),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_804),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_733),
.B(n_617),
.Y(n_873)
);

AND2x6_ASAP7_75t_SL g874 ( 
.A(n_759),
.B(n_767),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_738),
.B(n_624),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_748),
.B(n_661),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_738),
.B(n_624),
.Y(n_877)
);

INVx8_ASAP7_75t_L g878 ( 
.A(n_782),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_719),
.B(n_449),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_719),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_731),
.B(n_275),
.Y(n_881)
);

BUFx6f_ASAP7_75t_SL g882 ( 
.A(n_833),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_749),
.B(n_626),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_690),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_725),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_716),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_818),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_695),
.B(n_369),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_834),
.A2(n_731),
.B(n_708),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_749),
.B(n_626),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_756),
.B(n_633),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_728),
.B(n_678),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_729),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_756),
.B(n_633),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_716),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_756),
.A2(n_579),
.B(n_259),
.C(n_262),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_752),
.B(n_369),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_728),
.B(n_309),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_752),
.B(n_391),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_741),
.A2(n_455),
.B1(n_453),
.B2(n_269),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_704),
.A2(n_643),
.B(n_631),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_743),
.B(n_637),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_743),
.B(n_637),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_704),
.A2(n_643),
.B(n_631),
.Y(n_904)
);

AND2x6_ASAP7_75t_SL g905 ( 
.A(n_715),
.B(n_238),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_794),
.B(n_638),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_741),
.A2(n_269),
.B1(n_299),
.B2(n_250),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_786),
.B(n_391),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_718),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_729),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_777),
.B(n_638),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_786),
.B(n_410),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_753),
.B(n_410),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_741),
.A2(n_736),
.B1(n_783),
.B2(n_698),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_811),
.Y(n_915)
);

AOI22xp5_ASAP7_75t_L g916 ( 
.A1(n_736),
.A2(n_299),
.B1(n_303),
.B2(n_250),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_777),
.B(n_639),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_777),
.B(n_639),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_SL g919 ( 
.A1(n_814),
.A2(n_318),
.B1(n_384),
.B2(n_282),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_719),
.B(n_303),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_708),
.A2(n_643),
.B(n_631),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_730),
.B(n_322),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_730),
.B(n_322),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_736),
.A2(n_383),
.B1(n_352),
.B2(n_235),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_739),
.B(n_323),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_811),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_719),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_736),
.A2(n_383),
.B1(n_235),
.B2(n_236),
.Y(n_928)
);

INVxp33_ASAP7_75t_L g929 ( 
.A(n_820),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_792),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_739),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_719),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_737),
.B(n_340),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_804),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_683),
.B(n_323),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_684),
.B(n_333),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_801),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_801),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_737),
.B(n_340),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_709),
.B(n_333),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_792),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_734),
.A2(n_372),
.B(n_392),
.C(n_360),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_783),
.B(n_360),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_735),
.B(n_372),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_726),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_740),
.B(n_392),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_681),
.B(n_682),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_679),
.B(n_393),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_792),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_815),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_815),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_815),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_816),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_838),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_679),
.B(n_393),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_816),
.Y(n_956)
);

INVx8_ASAP7_75t_L g957 ( 
.A(n_782),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_783),
.B(n_721),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_721),
.B(n_397),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_812),
.B(n_397),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_689),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_736),
.B(n_407),
.Y(n_962)
);

NAND3xp33_ASAP7_75t_SL g963 ( 
.A(n_778),
.B(n_442),
.C(n_421),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_812),
.B(n_822),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_736),
.B(n_781),
.Y(n_965)
);

AND2x6_ASAP7_75t_SL g966 ( 
.A(n_715),
.B(n_240),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_820),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_702),
.B(n_421),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_802),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_773),
.B(n_233),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_781),
.B(n_407),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_688),
.B(n_237),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_802),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_715),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_816),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_772),
.B(n_309),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_828),
.B(n_411),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_751),
.B(n_236),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_715),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_805),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_805),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_698),
.A2(n_411),
.B1(n_452),
.B2(n_424),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_698),
.A2(n_452),
.B1(n_424),
.B2(n_416),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_831),
.B(n_642),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_698),
.A2(n_416),
.B1(n_435),
.B2(n_340),
.Y(n_985)
);

NOR3xp33_ASAP7_75t_SL g986 ( 
.A(n_760),
.B(n_244),
.C(n_239),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_785),
.A2(n_643),
.B(n_631),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_688),
.B(n_246),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_835),
.B(n_642),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_836),
.B(n_642),
.Y(n_990)
);

NAND2x1_ASAP7_75t_L g991 ( 
.A(n_689),
.B(n_641),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_812),
.B(n_642),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_813),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_813),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_822),
.B(n_642),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_839),
.B(n_642),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_727),
.B(n_642),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_686),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_766),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_L g1000 ( 
.A(n_698),
.B(n_248),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_822),
.B(n_340),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_727),
.B(n_641),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_727),
.B(n_645),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_814),
.B(n_782),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_692),
.B(n_645),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_766),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_692),
.B(n_536),
.Y(n_1007)
);

AND2x6_ASAP7_75t_SL g1008 ( 
.A(n_782),
.B(n_240),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_771),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_720),
.B(n_249),
.Y(n_1010)
);

OR2x2_ASAP7_75t_L g1011 ( 
.A(n_687),
.B(n_314),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_771),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_692),
.B(n_536),
.Y(n_1013)
);

AOI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_698),
.A2(n_416),
.B1(n_435),
.B2(n_454),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_927),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_927),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_866),
.B(n_824),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_856),
.B(n_926),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_848),
.A2(n_706),
.B1(n_705),
.B2(n_700),
.Y(n_1019)
);

INVx1_ASAP7_75t_SL g1020 ( 
.A(n_934),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_945),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_930),
.B(n_705),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_842),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_927),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_842),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_963),
.B(n_796),
.C(n_760),
.Y(n_1026)
);

AND3x1_ASAP7_75t_L g1027 ( 
.A(n_986),
.B(n_769),
.C(n_809),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_848),
.A2(n_700),
.B1(n_689),
.B2(n_705),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_905),
.Y(n_1029)
);

NOR3xp33_ASAP7_75t_SL g1030 ( 
.A(n_972),
.B(n_800),
.C(n_796),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_882),
.Y(n_1031)
);

AOI22xp33_ASAP7_75t_L g1032 ( 
.A1(n_888),
.A2(n_706),
.B1(n_705),
.B2(n_700),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_927),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_915),
.B(n_687),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_932),
.Y(n_1035)
);

AND2x2_ASAP7_75t_SL g1036 ( 
.A(n_854),
.B(n_810),
.Y(n_1036)
);

INVx5_ASAP7_75t_L g1037 ( 
.A(n_932),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_860),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_932),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_872),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_866),
.A2(n_700),
.B1(n_689),
.B2(n_705),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_932),
.Y(n_1042)
);

BUFx4f_ASAP7_75t_SL g1043 ( 
.A(n_844),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_892),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_847),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_845),
.B(n_800),
.Y(n_1046)
);

BUFx10_ASAP7_75t_L g1047 ( 
.A(n_882),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_860),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_913),
.B(n_840),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_SL g1050 ( 
.A(n_972),
.B(n_806),
.C(n_257),
.Y(n_1050)
);

AND2x4_ASAP7_75t_L g1051 ( 
.A(n_941),
.B(n_705),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_929),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_870),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_859),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_870),
.Y(n_1055)
);

AND3x1_ASAP7_75t_SL g1056 ( 
.A(n_909),
.B(n_242),
.C(n_241),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_888),
.A2(n_706),
.B1(n_755),
.B2(n_750),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_961),
.Y(n_1058)
);

NAND2x1_ASAP7_75t_L g1059 ( 
.A(n_961),
.B(n_699),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_964),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_885),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_SL g1062 ( 
.A(n_1004),
.B(n_827),
.Y(n_1062)
);

INVx6_ASAP7_75t_L g1063 ( 
.A(n_881),
.Y(n_1063)
);

NOR2x1_ASAP7_75t_L g1064 ( 
.A(n_933),
.B(n_768),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_908),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_885),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_893),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_893),
.Y(n_1068)
);

INVx6_ASAP7_75t_L g1069 ( 
.A(n_881),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_880),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_967),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_913),
.A2(n_761),
.B(n_750),
.C(n_807),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_910),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_851),
.B(n_765),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_L g1075 ( 
.A(n_843),
.B(n_791),
.C(n_806),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_910),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_931),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_L g1078 ( 
.A(n_843),
.B(n_425),
.C(n_314),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_862),
.B(n_686),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_931),
.Y(n_1080)
);

BUFx4f_ASAP7_75t_L g1081 ( 
.A(n_878),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_999),
.B(n_789),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_937),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_SL g1084 ( 
.A(n_865),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_968),
.A2(n_706),
.B1(n_755),
.B2(n_750),
.Y(n_1085)
);

OR2x2_ASAP7_75t_SL g1086 ( 
.A(n_1011),
.B(n_241),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_937),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_970),
.B(n_706),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_970),
.B(n_706),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_862),
.B(n_761),
.Y(n_1090)
);

OR2x2_ASAP7_75t_L g1091 ( 
.A(n_908),
.B(n_912),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_976),
.B(n_699),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_938),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_993),
.B(n_761),
.Y(n_1094)
);

HB1xp67_ASAP7_75t_L g1095 ( 
.A(n_865),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_841),
.Y(n_1096)
);

HB1xp67_ASAP7_75t_L g1097 ( 
.A(n_865),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_878),
.B(n_699),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_878),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_938),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_949),
.B(n_789),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_994),
.B(n_799),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_969),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_861),
.B(n_701),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_964),
.B(n_701),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_969),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_973),
.B(n_799),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_973),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_954),
.B(n_701),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_980),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_957),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_980),
.B(n_808),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_SL g1113 ( 
.A(n_974),
.B(n_790),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_950),
.B(n_951),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_981),
.B(n_808),
.Y(n_1115)
);

AND2x4_ASAP7_75t_L g1116 ( 
.A(n_952),
.B(n_837),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_981),
.B(n_837),
.Y(n_1117)
);

INVx3_ASAP7_75t_L g1118 ( 
.A(n_991),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_846),
.B(n_790),
.Y(n_1119)
);

NOR3xp33_ASAP7_75t_SL g1120 ( 
.A(n_988),
.B(n_265),
.C(n_251),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_978),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_850),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_968),
.A2(n_755),
.B1(n_779),
.B2(n_757),
.Y(n_1123)
);

INVx4_ASAP7_75t_L g1124 ( 
.A(n_957),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_SL g1125 ( 
.A(n_988),
.B(n_270),
.C(n_268),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_953),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1006),
.B(n_758),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_956),
.B(n_714),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_852),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_966),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1009),
.B(n_779),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_975),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_965),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_998),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_867),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1012),
.B(n_758),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_897),
.B(n_790),
.Y(n_1137)
);

BUFx12f_ASAP7_75t_L g1138 ( 
.A(n_1008),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_957),
.Y(n_1139)
);

NOR3xp33_ASAP7_75t_SL g1140 ( 
.A(n_912),
.B(n_276),
.C(n_274),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_884),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_874),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_886),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_895),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_992),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1007),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1013),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_891),
.B(n_754),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_894),
.B(n_775),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1005),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_SL g1151 ( 
.A(n_897),
.B(n_281),
.C(n_279),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_858),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_863),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_857),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_906),
.B(n_911),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_979),
.B(n_714),
.Y(n_1156)
);

NAND2xp33_ASAP7_75t_SL g1157 ( 
.A(n_887),
.B(n_242),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_871),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_978),
.Y(n_1159)
);

BUFx2_ASAP7_75t_L g1160 ( 
.A(n_978),
.Y(n_1160)
);

NOR3xp33_ASAP7_75t_SL g1161 ( 
.A(n_899),
.B(n_292),
.C(n_290),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_947),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_873),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_899),
.B(n_294),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_898),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_L g1166 ( 
.A(n_914),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_875),
.Y(n_1167)
);

BUFx2_ASAP7_75t_L g1168 ( 
.A(n_958),
.Y(n_1168)
);

AND2x2_ASAP7_75t_SL g1169 ( 
.A(n_854),
.B(n_810),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_948),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_984),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_917),
.B(n_776),
.Y(n_1172)
);

INVxp67_ASAP7_75t_SL g1173 ( 
.A(n_920),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_877),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_868),
.B(n_714),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_883),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_918),
.B(n_795),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_902),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_992),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_890),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_903),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_959),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_989),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1002),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1003),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_876),
.B(n_798),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_955),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_990),
.Y(n_1188)
);

BUFx5_ASAP7_75t_L g1189 ( 
.A(n_995),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_876),
.B(n_779),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_996),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_922),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_997),
.Y(n_1193)
);

BUFx2_ASAP7_75t_SL g1194 ( 
.A(n_995),
.Y(n_1194)
);

INVx3_ASAP7_75t_L g1195 ( 
.A(n_962),
.Y(n_1195)
);

BUFx8_ASAP7_75t_L g1196 ( 
.A(n_864),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_923),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_925),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_SL g1199 ( 
.A(n_919),
.B(n_300),
.C(n_295),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_907),
.Y(n_1200)
);

AND2x4_ASAP7_75t_L g1201 ( 
.A(n_868),
.B(n_714),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_924),
.B(n_707),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_924),
.B(n_707),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_889),
.B(n_712),
.Y(n_1204)
);

INVx4_ASAP7_75t_L g1205 ( 
.A(n_920),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_1000),
.B(n_301),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1010),
.B(n_307),
.Y(n_1207)
);

AO22x1_ASAP7_75t_L g1208 ( 
.A1(n_1010),
.A2(n_755),
.B1(n_264),
.B2(n_409),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_900),
.B(n_693),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_939),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_SL g1211 ( 
.A(n_1037),
.B(n_960),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1091),
.B(n_869),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1207),
.A2(n_855),
.B1(n_869),
.B2(n_943),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1066),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1049),
.B(n_935),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1066),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1048),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1048),
.Y(n_1218)
);

INVx2_ASAP7_75t_SL g1219 ( 
.A(n_1018),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1137),
.A2(n_879),
.B(n_849),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1122),
.A2(n_904),
.B(n_901),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1124),
.B(n_943),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1017),
.B(n_1174),
.Y(n_1223)
);

CKINVDCx8_ASAP7_75t_R g1224 ( 
.A(n_1021),
.Y(n_1224)
);

INVxp67_ASAP7_75t_SL g1225 ( 
.A(n_1070),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1180),
.B(n_936),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1037),
.A2(n_1039),
.B(n_1035),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1054),
.B(n_985),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1091),
.A2(n_928),
.B(n_853),
.C(n_896),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1124),
.B(n_1001),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1122),
.A2(n_921),
.B(n_879),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1037),
.A2(n_1001),
.B(n_960),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_SL g1233 ( 
.A1(n_1205),
.A2(n_944),
.B(n_940),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_1021),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_1044),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1139),
.B(n_797),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1099),
.Y(n_1237)
);

OA22x2_ASAP7_75t_L g1238 ( 
.A1(n_1065),
.A2(n_1014),
.B1(n_428),
.B2(n_425),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_1047),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1181),
.B(n_946),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1184),
.B(n_977),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1042),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1166),
.B(n_928),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1184),
.B(n_971),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1042),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1155),
.A2(n_987),
.B(n_916),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1185),
.B(n_983),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1037),
.A2(n_747),
.B(n_788),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1204),
.A2(n_817),
.B(n_797),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_L g1250 ( 
.A1(n_1164),
.A2(n_942),
.B(n_797),
.C(n_817),
.Y(n_1250)
);

NOR2xp33_ASAP7_75t_L g1251 ( 
.A(n_1054),
.B(n_982),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1040),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1105),
.A2(n_1195),
.B(n_1193),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1053),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1185),
.B(n_693),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1105),
.A2(n_1195),
.B(n_1193),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1035),
.A2(n_823),
.B(n_788),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1166),
.B(n_1145),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1100),
.Y(n_1259)
);

NAND2x1p5_ASAP7_75t_L g1260 ( 
.A(n_1139),
.B(n_817),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1128),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1037),
.A2(n_747),
.B(n_788),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1105),
.A2(n_770),
.B(n_764),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1195),
.A2(n_770),
.B(n_764),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1193),
.A2(n_780),
.B(n_703),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1061),
.A2(n_780),
.B(n_703),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1039),
.A2(n_747),
.B(n_788),
.Y(n_1267)
);

BUFx10_ASAP7_75t_L g1268 ( 
.A(n_1175),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1039),
.A2(n_1035),
.B(n_1088),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1173),
.A2(n_723),
.B(n_712),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1166),
.A2(n_1205),
.B1(n_1090),
.B2(n_1019),
.Y(n_1271)
);

O2A1O1Ixp5_ASAP7_75t_L g1272 ( 
.A1(n_1089),
.A2(n_398),
.B(n_264),
.C(n_285),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1061),
.A2(n_696),
.B(n_723),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1165),
.B(n_309),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1039),
.A2(n_747),
.B(n_788),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1061),
.A2(n_696),
.B(n_742),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1103),
.A2(n_763),
.B(n_742),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1158),
.B(n_763),
.Y(n_1278)
);

OAI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1072),
.A2(n_793),
.B(n_784),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1042),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1042),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1158),
.B(n_755),
.Y(n_1282)
);

OA22x2_ASAP7_75t_L g1283 ( 
.A1(n_1210),
.A2(n_428),
.B1(n_285),
.B2(n_413),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1039),
.A2(n_747),
.B(n_823),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1163),
.B(n_755),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1044),
.B(n_1079),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1103),
.A2(n_1055),
.B(n_1053),
.Y(n_1287)
);

OAI22x1_ASAP7_75t_L g1288 ( 
.A1(n_1200),
.A2(n_312),
.B1(n_451),
.B2(n_414),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1163),
.B(n_784),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1103),
.A2(n_819),
.B(n_793),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1205),
.A2(n_304),
.A3(n_457),
.B(n_450),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1082),
.B(n_309),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1167),
.B(n_819),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1042),
.A2(n_829),
.B(n_823),
.Y(n_1294)
);

NAND2x1p5_ASAP7_75t_L g1295 ( 
.A(n_1139),
.B(n_1124),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1055),
.A2(n_825),
.B(n_821),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1202),
.A2(n_825),
.B(n_821),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1099),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1067),
.A2(n_826),
.B(n_549),
.Y(n_1299)
);

BUFx12f_ASAP7_75t_L g1300 ( 
.A(n_1047),
.Y(n_1300)
);

INVx4_ASAP7_75t_L g1301 ( 
.A(n_1139),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1092),
.A2(n_1182),
.B(n_1190),
.Y(n_1302)
);

OAI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1028),
.A2(n_823),
.B1(n_830),
.B2(n_829),
.Y(n_1303)
);

AOI211x1_ASAP7_75t_L g1304 ( 
.A1(n_1199),
.A2(n_447),
.B(n_415),
.C(n_413),
.Y(n_1304)
);

NAND2x1_ASAP7_75t_L g1305 ( 
.A(n_1015),
.B(n_823),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1167),
.B(n_826),
.Y(n_1306)
);

INVx2_ASAP7_75t_SL g1307 ( 
.A(n_1018),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1067),
.A2(n_1073),
.B(n_1068),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1036),
.A2(n_1169),
.B(n_1129),
.C(n_1182),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1068),
.A2(n_549),
.B(n_547),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1020),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1186),
.A2(n_550),
.B(n_547),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1082),
.B(n_418),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1078),
.B(n_418),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1073),
.A2(n_552),
.B(n_550),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_SL g1316 ( 
.A1(n_1080),
.A2(n_315),
.B(n_304),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1176),
.B(n_803),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1059),
.A2(n_830),
.B(n_829),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1139),
.B(n_552),
.Y(n_1319)
);

AOI21xp33_ASAP7_75t_L g1320 ( 
.A1(n_1034),
.A2(n_320),
.B(n_310),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1076),
.Y(n_1321)
);

AOI22xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1096),
.A2(n_429),
.B1(n_373),
.B2(n_324),
.Y(n_1322)
);

AOI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1059),
.A2(n_830),
.B(n_829),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1076),
.A2(n_565),
.B(n_554),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1176),
.B(n_1129),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1203),
.A2(n_832),
.B(n_803),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1077),
.A2(n_565),
.B(n_554),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1077),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1045),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1052),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1188),
.A2(n_571),
.B(n_566),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1188),
.A2(n_571),
.B(n_566),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1171),
.A2(n_1183),
.B(n_1094),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1172),
.A2(n_830),
.B(n_829),
.Y(n_1334)
);

INVx8_ASAP7_75t_L g1335 ( 
.A(n_1098),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1162),
.B(n_1192),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1128),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1168),
.A2(n_440),
.A3(n_359),
.B(n_371),
.Y(n_1338)
);

O2A1O1Ixp5_ASAP7_75t_L g1339 ( 
.A1(n_1119),
.A2(n_450),
.B(n_315),
.C(n_398),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1145),
.B(n_830),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1162),
.B(n_803),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1023),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1036),
.A2(n_832),
.B(n_803),
.Y(n_1343)
);

INVx5_ASAP7_75t_L g1344 ( 
.A(n_1098),
.Y(n_1344)
);

INVx4_ASAP7_75t_SL g1345 ( 
.A(n_1098),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1071),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1171),
.A2(n_575),
.B(n_574),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1080),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1060),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1178),
.B(n_803),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1183),
.A2(n_575),
.B(n_574),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1071),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1168),
.A2(n_440),
.A3(n_371),
.B(n_381),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1178),
.B(n_803),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1025),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1038),
.A2(n_581),
.B(n_578),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1083),
.A2(n_581),
.B(n_578),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1134),
.B(n_325),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1111),
.B(n_101),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1087),
.A2(n_415),
.B(n_381),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1170),
.B(n_832),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1197),
.B(n_1198),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1177),
.A2(n_832),
.B(n_409),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1169),
.A2(n_832),
.B(n_774),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1209),
.A2(n_832),
.B(n_774),
.Y(n_1365)
);

AND2x2_ASAP7_75t_SL g1366 ( 
.A(n_1200),
.B(n_359),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1041),
.A2(n_405),
.B1(n_339),
.B2(n_456),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1134),
.B(n_330),
.Y(n_1368)
);

NAND2x1_ASAP7_75t_L g1369 ( 
.A(n_1015),
.B(n_774),
.Y(n_1369)
);

INVx3_ASAP7_75t_SL g1370 ( 
.A(n_1031),
.Y(n_1370)
);

OAI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1109),
.A2(n_774),
.B(n_457),
.Y(n_1371)
);

AO21x1_ASAP7_75t_L g1372 ( 
.A1(n_1062),
.A2(n_388),
.B(n_432),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1197),
.B(n_332),
.Y(n_1373)
);

AOI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1093),
.A2(n_447),
.B(n_432),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1210),
.B(n_336),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1106),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1108),
.A2(n_388),
.B(n_774),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1032),
.A2(n_412),
.B1(n_446),
.B2(n_445),
.Y(n_1378)
);

NAND2x1_ASAP7_75t_L g1379 ( 
.A(n_1015),
.B(n_774),
.Y(n_1379)
);

NAND2x1_ASAP7_75t_L g1380 ( 
.A(n_1301),
.B(n_1060),
.Y(n_1380)
);

OR2x2_ASAP7_75t_L g1381 ( 
.A(n_1212),
.B(n_1107),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1217),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1234),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1212),
.B(n_1112),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1345),
.B(n_1111),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1213),
.A2(n_1069),
.B1(n_1063),
.B2(n_1081),
.Y(n_1386)
);

INVx1_ASAP7_75t_SL g1387 ( 
.A(n_1330),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1344),
.B(n_1060),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1253),
.A2(n_1110),
.B(n_1127),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1233),
.A2(n_1206),
.B(n_1117),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1257),
.A2(n_1104),
.B(n_1198),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1366),
.A2(n_1096),
.B1(n_1062),
.B2(n_1074),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1253),
.A2(n_1136),
.B(n_1115),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1345),
.B(n_1114),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1220),
.A2(n_1064),
.B(n_1151),
.C(n_1140),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1366),
.A2(n_1069),
.B1(n_1063),
.B2(n_1114),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1256),
.A2(n_1191),
.B(n_1149),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1345),
.B(n_1114),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1223),
.A2(n_1069),
.B1(n_1063),
.B2(n_1081),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1217),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1286),
.B(n_1034),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1375),
.B(n_1161),
.C(n_1125),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1218),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1234),
.Y(n_1404)
);

NAND2x1_ASAP7_75t_L g1405 ( 
.A(n_1301),
.B(n_1060),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1256),
.A2(n_1148),
.B(n_1152),
.Y(n_1406)
);

OAI21xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1243),
.A2(n_1057),
.B(n_1102),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1265),
.A2(n_1264),
.B(n_1287),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1215),
.B(n_1131),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1249),
.A2(n_1150),
.B(n_1209),
.Y(n_1410)
);

INVx4_ASAP7_75t_L g1411 ( 
.A(n_1335),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1309),
.B(n_1131),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1375),
.A2(n_1075),
.B1(n_1027),
.B2(n_1069),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1261),
.B(n_1101),
.Y(n_1414)
);

AO32x2_ASAP7_75t_L g1415 ( 
.A1(n_1271),
.A2(n_1144),
.A3(n_1135),
.B1(n_1056),
.B2(n_1086),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1265),
.A2(n_1264),
.B(n_1287),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1218),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1336),
.B(n_1150),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1249),
.A2(n_1147),
.B(n_1132),
.Y(n_1419)
);

AOI22x1_ASAP7_75t_L g1420 ( 
.A1(n_1302),
.A2(n_1194),
.B1(n_1145),
.B2(n_1179),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1254),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1362),
.B(n_1187),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1237),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1254),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1309),
.A2(n_1123),
.B(n_1085),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1308),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_L g1427 ( 
.A(n_1242),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1347),
.A2(n_1147),
.B(n_1146),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1347),
.A2(n_1146),
.B(n_1143),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1352),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1247),
.A2(n_1116),
.B(n_1101),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1296),
.A2(n_1152),
.B(n_1118),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1279),
.A2(n_1126),
.B(n_1143),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1229),
.A2(n_1116),
.B(n_1101),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1226),
.A2(n_1026),
.B(n_1187),
.C(n_1120),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1311),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1240),
.B(n_1116),
.Y(n_1437)
);

NOR2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1239),
.B(n_1031),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1333),
.A2(n_1208),
.B(n_1153),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1344),
.B(n_1060),
.Y(n_1440)
);

AND2x6_ASAP7_75t_L g1441 ( 
.A(n_1230),
.B(n_1145),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1296),
.A2(n_1152),
.B(n_1118),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_SL g1443 ( 
.A1(n_1258),
.A2(n_1243),
.B(n_1229),
.C(n_1340),
.Y(n_1443)
);

AO21x2_ASAP7_75t_L g1444 ( 
.A1(n_1372),
.A2(n_1153),
.B(n_1050),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1299),
.A2(n_1118),
.B(n_1024),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1228),
.A2(n_1063),
.B1(n_1144),
.B2(n_1157),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1299),
.A2(n_1024),
.B(n_1016),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1308),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1325),
.B(n_1145),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1333),
.A2(n_1351),
.B(n_1312),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1355),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1301),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1310),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1214),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1241),
.B(n_1135),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1246),
.A2(n_1113),
.B(n_1133),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1251),
.A2(n_1142),
.B1(n_1121),
.B2(n_1095),
.Y(n_1457)
);

AOI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1251),
.A2(n_1142),
.B1(n_1097),
.B2(n_1084),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1331),
.A2(n_1024),
.B(n_1016),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1331),
.A2(n_1033),
.B(n_1016),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1352),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1216),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1225),
.A2(n_1081),
.B1(n_1194),
.B2(n_1179),
.Y(n_1463)
);

CKINVDCx9p33_ASAP7_75t_R g1464 ( 
.A(n_1235),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1332),
.A2(n_1033),
.B(n_1058),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1258),
.B(n_1086),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1244),
.A2(n_1113),
.B(n_1133),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_1224),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1332),
.A2(n_1033),
.B(n_1058),
.Y(n_1469)
);

CKINVDCx14_ASAP7_75t_R g1470 ( 
.A(n_1311),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1351),
.A2(n_1058),
.B(n_1189),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1266),
.A2(n_1189),
.B(n_1133),
.Y(n_1472)
);

OAI222xp33_ASAP7_75t_L g1473 ( 
.A1(n_1238),
.A2(n_1154),
.B1(n_389),
.B2(n_390),
.C1(n_394),
.C2(n_430),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1320),
.B(n_1030),
.C(n_1157),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1230),
.A2(n_1179),
.B1(n_1144),
.B2(n_1133),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1314),
.A2(n_1160),
.B1(n_1141),
.B2(n_1159),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1292),
.B(n_1179),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1266),
.A2(n_1189),
.B(n_1133),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1373),
.B(n_1189),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1261),
.B(n_1098),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1259),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1289),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1290),
.A2(n_1189),
.B(n_1179),
.Y(n_1483)
);

NAND2x1p5_ASAP7_75t_L g1484 ( 
.A(n_1344),
.B(n_1141),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1290),
.A2(n_1189),
.B(n_1208),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1307),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1273),
.A2(n_1189),
.B(n_1141),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1238),
.A2(n_1160),
.B1(n_1141),
.B2(n_1084),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1273),
.A2(n_1276),
.B(n_1263),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1337),
.B(n_1156),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1288),
.A2(n_1313),
.B1(n_1219),
.B2(n_1378),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1293),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1346),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1276),
.A2(n_1141),
.B(n_1022),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1310),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1315),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1219),
.B(n_1201),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1315),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1263),
.A2(n_1022),
.B(n_1051),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1306),
.Y(n_1500)
);

INVx6_ASAP7_75t_L g1501 ( 
.A(n_1268),
.Y(n_1501)
);

OAI21xp33_ASAP7_75t_L g1502 ( 
.A1(n_1274),
.A2(n_1046),
.B(n_1154),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1277),
.A2(n_1022),
.B(n_1051),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1277),
.A2(n_1051),
.B(n_1175),
.Y(n_1504)
);

AO31x2_ASAP7_75t_L g1505 ( 
.A1(n_1303),
.A2(n_1201),
.A3(n_1175),
.B(n_10),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1231),
.A2(n_1201),
.B(n_1084),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1230),
.A2(n_1043),
.B1(n_1156),
.B2(n_1128),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1337),
.B(n_1156),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1231),
.A2(n_1047),
.B(n_116),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1329),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1367),
.A2(n_416),
.B1(n_435),
.B2(n_1130),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1344),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1255),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1324),
.A2(n_115),
.B(n_110),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1324),
.A2(n_1327),
.B(n_1221),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_SL g1516 ( 
.A1(n_1211),
.A2(n_117),
.B(n_230),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1359),
.B(n_124),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1322),
.B(n_1196),
.C(n_420),
.Y(n_1518)
);

O2A1O1Ixp33_ASAP7_75t_L g1519 ( 
.A1(n_1252),
.A2(n_1316),
.B(n_1358),
.C(n_1368),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1327),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1348),
.B(n_1342),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1376),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1348),
.A2(n_1029),
.B1(n_1130),
.B2(n_1138),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1278),
.B(n_337),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1321),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1328),
.B(n_344),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1359),
.B(n_129),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1221),
.A2(n_197),
.B(n_141),
.Y(n_1528)
);

INVx3_ASAP7_75t_L g1529 ( 
.A(n_1335),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1291),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1224),
.B(n_1029),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1356),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1370),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1356),
.A2(n_198),
.B(n_147),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1312),
.A2(n_435),
.B(n_202),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1272),
.A2(n_441),
.B(n_439),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1357),
.A2(n_186),
.B(n_152),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1357),
.A2(n_205),
.B(n_154),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1349),
.B(n_275),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1349),
.B(n_382),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1370),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_L g1542 ( 
.A1(n_1269),
.A2(n_208),
.B(n_224),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1360),
.A2(n_438),
.B(n_434),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1360),
.A2(n_180),
.B(n_223),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1359),
.B(n_356),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1237),
.B(n_1138),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1283),
.A2(n_382),
.B1(n_418),
.B2(n_1196),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1250),
.A2(n_427),
.B(n_423),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1349),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1298),
.B(n_138),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1349),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1298),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_1239),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1335),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1365),
.A2(n_178),
.B(n_220),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1300),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1291),
.Y(n_1557)
);

INVx2_ASAP7_75t_SL g1558 ( 
.A(n_1268),
.Y(n_1558)
);

NAND3xp33_ASAP7_75t_L g1559 ( 
.A(n_1304),
.B(n_1196),
.C(n_422),
.Y(n_1559)
);

INVxp67_ASAP7_75t_SL g1560 ( 
.A(n_1242),
.Y(n_1560)
);

BUFx4f_ASAP7_75t_SL g1561 ( 
.A(n_1300),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1319),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1297),
.A2(n_172),
.B(n_218),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1232),
.A2(n_158),
.B(n_159),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1400),
.Y(n_1565)
);

NAND2xp33_ASAP7_75t_SL g1566 ( 
.A(n_1517),
.B(n_1242),
.Y(n_1566)
);

OAI221xp5_ASAP7_75t_L g1567 ( 
.A1(n_1392),
.A2(n_1283),
.B1(n_1339),
.B2(n_1371),
.C(n_1361),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1401),
.B(n_1340),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1413),
.A2(n_1222),
.B1(n_1341),
.B2(n_1350),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1511),
.A2(n_1363),
.B1(n_1334),
.B2(n_1364),
.C(n_1343),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1402),
.A2(n_382),
.B1(n_418),
.B2(n_1222),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1409),
.B(n_1222),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1462),
.Y(n_1573)
);

AOI21xp33_ASAP7_75t_L g1574 ( 
.A1(n_1381),
.A2(n_1384),
.B(n_1519),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1394),
.Y(n_1575)
);

AO31x2_ASAP7_75t_L g1576 ( 
.A1(n_1530),
.A2(n_1317),
.A3(n_1354),
.B(n_1285),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1515),
.A2(n_1557),
.B(n_1416),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1381),
.A2(n_358),
.B1(n_363),
.B2(n_380),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1425),
.A2(n_1326),
.B(n_1282),
.C(n_1270),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1394),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1434),
.B(n_1295),
.Y(n_1581)
);

NOR2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1404),
.B(n_1374),
.Y(n_1582)
);

OAI222xp33_ASAP7_75t_L g1583 ( 
.A1(n_1466),
.A2(n_385),
.B1(n_396),
.B2(n_402),
.C1(n_1319),
.C2(n_1295),
.Y(n_1583)
);

OAI221xp5_ASAP7_75t_L g1584 ( 
.A1(n_1502),
.A2(n_1236),
.B1(n_1260),
.B2(n_1305),
.C(n_1369),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1418),
.B(n_1338),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1468),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_1468),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1474),
.A2(n_1319),
.B1(n_1268),
.B2(n_1281),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1400),
.Y(n_1589)
);

NAND2xp33_ASAP7_75t_SL g1590 ( 
.A(n_1552),
.B(n_1242),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1477),
.B(n_1539),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1477),
.B(n_1338),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1403),
.Y(n_1593)
);

INVx4_ASAP7_75t_L g1594 ( 
.A(n_1423),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1539),
.B(n_1338),
.Y(n_1595)
);

AOI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1384),
.A2(n_1280),
.B1(n_1281),
.B2(n_1245),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1423),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1473),
.A2(n_1547),
.B1(n_1536),
.B2(n_1548),
.C(n_1491),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1552),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1446),
.A2(n_1281),
.B1(n_1280),
.B2(n_1260),
.Y(n_1600)
);

OAI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1466),
.A2(n_1236),
.B1(n_1379),
.B2(n_1280),
.Y(n_1601)
);

CKINVDCx6p67_ASAP7_75t_R g1602 ( 
.A(n_1541),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1394),
.Y(n_1603)
);

AO221x1_ASAP7_75t_L g1604 ( 
.A1(n_1516),
.A2(n_1245),
.B1(n_1291),
.B2(n_1338),
.C(n_1353),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1427),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1385),
.B(n_1245),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1427),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1481),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1436),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1395),
.B(n_1245),
.C(n_1294),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1436),
.B(n_1353),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1454),
.Y(n_1612)
);

AOI21xp33_ASAP7_75t_L g1613 ( 
.A1(n_1431),
.A2(n_1377),
.B(n_1323),
.Y(n_1613)
);

INVx2_ASAP7_75t_SL g1614 ( 
.A(n_1387),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1385),
.B(n_1353),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1522),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1403),
.Y(n_1617)
);

NAND3xp33_ASAP7_75t_SL g1618 ( 
.A(n_1435),
.B(n_1458),
.C(n_1476),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1518),
.A2(n_1318),
.B1(n_1353),
.B2(n_1227),
.C(n_1291),
.Y(n_1619)
);

BUFx4f_ASAP7_75t_SL g1620 ( 
.A(n_1541),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1521),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1510),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1540),
.B(n_8),
.Y(n_1623)
);

AO21x2_ASAP7_75t_L g1624 ( 
.A1(n_1439),
.A2(n_1377),
.B(n_1284),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1451),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1385),
.B(n_1398),
.Y(n_1626)
);

AOI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1470),
.A2(n_1275),
.B1(n_1267),
.B2(n_1262),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1559),
.A2(n_1412),
.B1(n_1437),
.B2(n_1488),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1383),
.Y(n_1629)
);

INVx5_ASAP7_75t_L g1630 ( 
.A(n_1427),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1430),
.B(n_1461),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1497),
.B(n_1486),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1421),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1525),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1457),
.A2(n_1248),
.B1(n_10),
.B2(n_11),
.Y(n_1635)
);

NAND2x1_ASAP7_75t_L g1636 ( 
.A(n_1512),
.B(n_212),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1396),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_1637)
);

INVx3_ASAP7_75t_L g1638 ( 
.A(n_1398),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1515),
.A2(n_209),
.B(n_164),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1540),
.B(n_14),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1493),
.Y(n_1641)
);

AND2x2_ASAP7_75t_SL g1642 ( 
.A(n_1517),
.B(n_15),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1412),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1517),
.A2(n_16),
.B1(n_21),
.B2(n_23),
.Y(n_1644)
);

BUFx3_ASAP7_75t_L g1645 ( 
.A(n_1493),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1449),
.B(n_23),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1421),
.Y(n_1647)
);

AOI21xp33_ASAP7_75t_L g1648 ( 
.A1(n_1479),
.A2(n_24),
.B(n_26),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1382),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1407),
.A2(n_24),
.B(n_27),
.Y(n_1650)
);

NAND2x1_ASAP7_75t_L g1651 ( 
.A(n_1512),
.B(n_28),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1439),
.A2(n_29),
.B(n_33),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1455),
.B(n_29),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1427),
.Y(n_1654)
);

O2A1O1Ixp33_ASAP7_75t_SL g1655 ( 
.A1(n_1380),
.A2(n_34),
.B(n_40),
.C(n_42),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1417),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1417),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1527),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1398),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1404),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1527),
.A2(n_1545),
.B1(n_1386),
.B2(n_1441),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1411),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1464),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1422),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_1664)
);

INVx2_ASAP7_75t_SL g1665 ( 
.A(n_1533),
.Y(n_1665)
);

AO32x2_ASAP7_75t_L g1666 ( 
.A1(n_1475),
.A2(n_48),
.A3(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1497),
.B(n_52),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_R g1668 ( 
.A(n_1527),
.B(n_98),
.Y(n_1668)
);

CKINVDCx6p67_ASAP7_75t_R g1669 ( 
.A(n_1550),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1424),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1444),
.A2(n_98),
.B1(n_58),
.B2(n_59),
.Y(n_1671)
);

NAND2xp33_ASAP7_75t_L g1672 ( 
.A(n_1441),
.B(n_57),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1449),
.B(n_61),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1443),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.C(n_65),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1524),
.B(n_64),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1482),
.B(n_65),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1441),
.A2(n_96),
.B1(n_74),
.B2(n_76),
.Y(n_1677)
);

AOI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1444),
.A2(n_1492),
.B1(n_1482),
.B2(n_1500),
.Y(n_1678)
);

A2O1A1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1391),
.A2(n_69),
.B(n_74),
.C(n_76),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1444),
.A2(n_95),
.B1(n_78),
.B2(n_81),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_R g1681 ( 
.A(n_1383),
.B(n_77),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1507),
.A2(n_77),
.B1(n_82),
.B2(n_83),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1526),
.A2(n_83),
.B1(n_84),
.B2(n_87),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1549),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1408),
.A2(n_87),
.B(n_90),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1463),
.A2(n_92),
.B1(n_93),
.B2(n_1411),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1549),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1492),
.B(n_92),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1551),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1414),
.B(n_1508),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1500),
.B(n_1513),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1456),
.A2(n_1467),
.B(n_1397),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1411),
.A2(n_1554),
.B1(n_1513),
.B2(n_1388),
.Y(n_1693)
);

AOI21xp33_ASAP7_75t_L g1694 ( 
.A1(n_1399),
.A2(n_1562),
.B(n_1420),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1414),
.A2(n_1531),
.B1(n_1523),
.B2(n_1550),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1554),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1426),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1554),
.B(n_1414),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1484),
.A2(n_1480),
.B(n_1550),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1433),
.A2(n_1562),
.B1(n_1441),
.B2(n_1535),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1433),
.A2(n_1441),
.B1(n_1535),
.B2(n_1516),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1397),
.A2(n_1393),
.B(n_1389),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1529),
.B(n_1480),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1448),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1546),
.Y(n_1705)
);

OAI221xp5_ASAP7_75t_L g1706 ( 
.A1(n_1564),
.A2(n_1420),
.B1(n_1553),
.B2(n_1556),
.C(n_1440),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_SL g1707 ( 
.A(n_1553),
.B(n_1556),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1448),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1429),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1429),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1551),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1433),
.A2(n_1441),
.B1(n_1535),
.B2(n_1480),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1560),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1508),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1561),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1427),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1388),
.A2(n_1440),
.B1(n_1484),
.B2(n_1501),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1388),
.A2(n_1440),
.B1(n_1543),
.B2(n_1490),
.C(n_1529),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1529),
.A2(n_1543),
.B1(n_1563),
.B2(n_1390),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1484),
.A2(n_1501),
.B1(n_1558),
.B2(n_1512),
.Y(n_1720)
);

INVxp67_ASAP7_75t_L g1721 ( 
.A(n_1438),
.Y(n_1721)
);

AOI22xp33_ASAP7_75t_L g1722 ( 
.A1(n_1543),
.A2(n_1563),
.B1(n_1390),
.B2(n_1558),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1429),
.Y(n_1723)
);

AO21x1_ASAP7_75t_SL g1724 ( 
.A1(n_1415),
.A2(n_1505),
.B(n_1555),
.Y(n_1724)
);

CKINVDCx5p33_ASAP7_75t_R g1725 ( 
.A(n_1501),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1415),
.Y(n_1726)
);

OAI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1501),
.A2(n_1380),
.B1(n_1405),
.B2(n_1452),
.Y(n_1727)
);

NAND3xp33_ASAP7_75t_SL g1728 ( 
.A(n_1405),
.B(n_1532),
.C(n_1415),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1415),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1390),
.A2(n_1410),
.B1(n_1542),
.B2(n_1544),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1452),
.B(n_1499),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1410),
.A2(n_1542),
.B1(n_1544),
.B2(n_1419),
.Y(n_1732)
);

CKINVDCx5p33_ASAP7_75t_R g1733 ( 
.A(n_1452),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1410),
.A2(n_1419),
.B1(n_1428),
.B2(n_1393),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1506),
.Y(n_1735)
);

INVx2_ASAP7_75t_SL g1736 ( 
.A(n_1506),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1415),
.B(n_1505),
.Y(n_1737)
);

OAI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1428),
.A2(n_1498),
.B1(n_1495),
.B2(n_1520),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1499),
.B(n_1503),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1505),
.B(n_1503),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1505),
.Y(n_1741)
);

AO31x2_ASAP7_75t_L g1742 ( 
.A1(n_1532),
.A2(n_1520),
.A3(n_1498),
.B(n_1496),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1504),
.B(n_1428),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1505),
.Y(n_1744)
);

AOI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1504),
.A2(n_1555),
.B1(n_1494),
.B2(n_1528),
.Y(n_1745)
);

CKINVDCx6p67_ASAP7_75t_R g1746 ( 
.A(n_1509),
.Y(n_1746)
);

INVx4_ASAP7_75t_L g1747 ( 
.A(n_1419),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1389),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1450),
.B(n_1494),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_L g1750 ( 
.A1(n_1453),
.A2(n_1496),
.B1(n_1450),
.B2(n_1528),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1534),
.A2(n_1538),
.B1(n_1537),
.B2(n_1514),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1483),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1509),
.B(n_1538),
.C(n_1537),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1534),
.A2(n_1514),
.B1(n_1450),
.B2(n_1478),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1485),
.A2(n_1406),
.B1(n_1471),
.B2(n_1442),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1487),
.Y(n_1756)
);

BUFx12f_ASAP7_75t_L g1757 ( 
.A(n_1471),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1487),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1432),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1432),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_SL g1761 ( 
.A1(n_1642),
.A2(n_1485),
.B1(n_1472),
.B2(n_1478),
.Y(n_1761)
);

INVx5_ASAP7_75t_L g1762 ( 
.A(n_1757),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1695),
.A2(n_1669),
.B1(n_1578),
.B2(n_1628),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1621),
.B(n_1472),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1578),
.A2(n_1442),
.B1(n_1469),
.B2(n_1465),
.Y(n_1765)
);

AOI22x1_ASAP7_75t_L g1766 ( 
.A1(n_1582),
.A2(n_1469),
.B1(n_1465),
.B2(n_1459),
.Y(n_1766)
);

AOI222xp33_ASAP7_75t_L g1767 ( 
.A1(n_1598),
.A2(n_1459),
.B1(n_1460),
.B2(n_1445),
.C1(n_1447),
.C2(n_1408),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1599),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1679),
.A2(n_1445),
.B(n_1460),
.Y(n_1769)
);

INVx3_ASAP7_75t_L g1770 ( 
.A(n_1626),
.Y(n_1770)
);

BUFx3_ASAP7_75t_L g1771 ( 
.A(n_1641),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1674),
.A2(n_1447),
.B1(n_1416),
.B2(n_1489),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1642),
.A2(n_1489),
.B1(n_1618),
.B2(n_1643),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1591),
.B(n_1646),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_L g1775 ( 
.A1(n_1644),
.A2(n_1658),
.B1(n_1571),
.B2(n_1643),
.C(n_1675),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1623),
.B(n_1640),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1683),
.A2(n_1644),
.B1(n_1658),
.B2(n_1680),
.Y(n_1777)
);

OAI222xp33_ASAP7_75t_L g1778 ( 
.A1(n_1671),
.A2(n_1680),
.B1(n_1677),
.B2(n_1683),
.C1(n_1664),
.C2(n_1637),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1592),
.B(n_1595),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1599),
.Y(n_1780)
);

OAI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1571),
.A2(n_1679),
.B1(n_1668),
.B2(n_1672),
.C(n_1671),
.Y(n_1781)
);

INVx8_ASAP7_75t_L g1782 ( 
.A(n_1630),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1714),
.B(n_1690),
.Y(n_1783)
);

INVx11_ASAP7_75t_L g1784 ( 
.A(n_1757),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1573),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1566),
.A2(n_1692),
.B(n_1699),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1668),
.A2(n_1628),
.B1(n_1650),
.B2(n_1635),
.C(n_1661),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1705),
.B(n_1622),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1690),
.B(n_1632),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1681),
.A2(n_1648),
.B1(n_1574),
.B2(n_1682),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1614),
.B(n_1586),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1634),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1681),
.A2(n_1568),
.B1(n_1567),
.B2(n_1653),
.Y(n_1793)
);

BUFx4f_ASAP7_75t_L g1794 ( 
.A(n_1602),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1611),
.B(n_1673),
.Y(n_1795)
);

INVx5_ASAP7_75t_L g1796 ( 
.A(n_1581),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1663),
.A2(n_1568),
.B1(n_1665),
.B2(n_1572),
.Y(n_1797)
);

OAI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1660),
.A2(n_1596),
.B1(n_1588),
.B2(n_1706),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1703),
.B(n_1609),
.Y(n_1799)
);

AOI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1721),
.A2(n_1566),
.B1(n_1590),
.B2(n_1587),
.Y(n_1800)
);

OAI211xp5_ASAP7_75t_SL g1801 ( 
.A1(n_1676),
.A2(n_1688),
.B(n_1619),
.C(n_1678),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1632),
.B(n_1667),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1608),
.Y(n_1803)
);

OAI222xp33_ASAP7_75t_L g1804 ( 
.A1(n_1686),
.A2(n_1581),
.B1(n_1691),
.B2(n_1741),
.C1(n_1569),
.C2(n_1737),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1631),
.B(n_1645),
.Y(n_1805)
);

OAI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1655),
.A2(n_1631),
.B(n_1678),
.C(n_1712),
.Y(n_1806)
);

AOI22xp33_ASAP7_75t_L g1807 ( 
.A1(n_1615),
.A2(n_1620),
.B1(n_1581),
.B2(n_1645),
.Y(n_1807)
);

OAI211xp5_ASAP7_75t_L g1808 ( 
.A1(n_1655),
.A2(n_1712),
.B(n_1700),
.C(n_1585),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1713),
.B(n_1575),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1652),
.A2(n_1620),
.B1(n_1666),
.B2(n_1604),
.Y(n_1810)
);

AND2x4_ASAP7_75t_L g1811 ( 
.A(n_1575),
.B(n_1580),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1583),
.A2(n_1744),
.B1(n_1570),
.B2(n_1694),
.C(n_1700),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1616),
.Y(n_1813)
);

OAI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1596),
.A2(n_1733),
.B1(n_1725),
.B2(n_1629),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1652),
.A2(n_1744),
.B1(n_1625),
.B2(n_1698),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1666),
.A2(n_1685),
.B1(n_1726),
.B2(n_1729),
.Y(n_1816)
);

AOI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1610),
.A2(n_1698),
.B1(n_1659),
.B2(n_1603),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_SL g1818 ( 
.A1(n_1666),
.A2(n_1720),
.B1(n_1693),
.B2(n_1740),
.Y(n_1818)
);

OAI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1651),
.A2(n_1666),
.B1(n_1597),
.B2(n_1594),
.Y(n_1819)
);

BUFx5_ASAP7_75t_L g1820 ( 
.A(n_1760),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1707),
.A2(n_1638),
.B1(n_1659),
.B2(n_1627),
.Y(n_1821)
);

INVxp67_ASAP7_75t_R g1822 ( 
.A(n_1639),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1638),
.A2(n_1670),
.B1(n_1656),
.B2(n_1657),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1606),
.B(n_1594),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1715),
.B(n_1597),
.Y(n_1825)
);

AOI211xp5_ASAP7_75t_SL g1826 ( 
.A1(n_1601),
.A2(n_1718),
.B(n_1717),
.C(n_1584),
.Y(n_1826)
);

OAI211xp5_ASAP7_75t_L g1827 ( 
.A1(n_1701),
.A2(n_1722),
.B(n_1719),
.C(n_1732),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1701),
.A2(n_1696),
.B1(n_1662),
.B2(n_1579),
.Y(n_1828)
);

AO31x2_ASAP7_75t_L g1829 ( 
.A1(n_1747),
.A2(n_1748),
.A3(n_1749),
.B(n_1743),
.Y(n_1829)
);

AOI322xp5_ASAP7_75t_L g1830 ( 
.A1(n_1649),
.A2(n_1728),
.A3(n_1689),
.B1(n_1687),
.B2(n_1684),
.C1(n_1711),
.C2(n_1636),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1579),
.A2(n_1613),
.B(n_1751),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1606),
.B(n_1662),
.Y(n_1832)
);

AOI21xp33_ASAP7_75t_L g1833 ( 
.A1(n_1722),
.A2(n_1719),
.B(n_1600),
.Y(n_1833)
);

AOI222xp33_ASAP7_75t_L g1834 ( 
.A1(n_1565),
.A2(n_1647),
.B1(n_1617),
.B2(n_1589),
.C1(n_1593),
.C2(n_1633),
.Y(n_1834)
);

OAI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1727),
.A2(n_1730),
.B(n_1745),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1696),
.A2(n_1730),
.B1(n_1732),
.B2(n_1630),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1724),
.A2(n_1565),
.B1(n_1647),
.B2(n_1589),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1716),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1630),
.A2(n_1654),
.B1(n_1607),
.B2(n_1605),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1731),
.A2(n_1739),
.B1(n_1746),
.B2(n_1736),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1630),
.A2(n_1754),
.B1(n_1593),
.B2(n_1633),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1742),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1617),
.B(n_1605),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1697),
.A2(n_1704),
.B1(n_1708),
.B2(n_1747),
.Y(n_1844)
);

BUFx12f_ASAP7_75t_L g1845 ( 
.A(n_1607),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1607),
.B(n_1654),
.Y(n_1846)
);

OAI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1753),
.A2(n_1702),
.B1(n_1750),
.B2(n_1755),
.C(n_1734),
.Y(n_1847)
);

BUFx12f_ASAP7_75t_L g1848 ( 
.A(n_1654),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1735),
.A2(n_1756),
.B1(n_1743),
.B2(n_1758),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1742),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1735),
.A2(n_1752),
.B1(n_1624),
.B2(n_1759),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1742),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1576),
.B(n_1742),
.Y(n_1853)
);

INVx4_ASAP7_75t_L g1854 ( 
.A(n_1624),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1734),
.A2(n_1752),
.B1(n_1759),
.B2(n_1738),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1709),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1576),
.B(n_1577),
.Y(n_1857)
);

OAI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1710),
.A2(n_1723),
.B1(n_1738),
.B2(n_1577),
.Y(n_1858)
);

AOI222xp33_ASAP7_75t_L g1859 ( 
.A1(n_1710),
.A2(n_1576),
.B1(n_1577),
.B2(n_1723),
.C1(n_1366),
.C2(n_1199),
.Y(n_1859)
);

OAI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1576),
.A2(n_1668),
.B1(n_1091),
.B2(n_1674),
.Y(n_1860)
);

BUFx3_ASAP7_75t_L g1861 ( 
.A(n_1641),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1629),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1683),
.A2(n_604),
.B1(n_1164),
.B2(n_685),
.C(n_1079),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1621),
.B(n_1568),
.Y(n_1864)
);

AOI222xp33_ASAP7_75t_L g1865 ( 
.A1(n_1598),
.A2(n_1366),
.B1(n_1199),
.B2(n_1164),
.C1(n_888),
.C2(n_604),
.Y(n_1865)
);

BUFx12f_ASAP7_75t_L g1866 ( 
.A(n_1715),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1611),
.B(n_1592),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1744),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1642),
.A2(n_1672),
.B1(n_1366),
.B2(n_673),
.Y(n_1870)
);

OAI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1668),
.A2(n_1091),
.B1(n_1674),
.B2(n_1213),
.Y(n_1871)
);

AOI22xp33_ASAP7_75t_L g1872 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1872)
);

OAI22xp5_ASAP7_75t_L g1873 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1629),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1703),
.B(n_1609),
.Y(n_1875)
);

AOI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1672),
.A2(n_1391),
.B(n_1220),
.Y(n_1876)
);

OAI211xp5_ASAP7_75t_L g1877 ( 
.A1(n_1644),
.A2(n_685),
.B(n_919),
.C(n_1079),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1705),
.B(n_843),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1611),
.B(n_1592),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1621),
.B(n_1568),
.Y(n_1881)
);

AOI221xp5_ASAP7_75t_L g1882 ( 
.A1(n_1683),
.A2(n_604),
.B1(n_1164),
.B2(n_685),
.C(n_1079),
.Y(n_1882)
);

AOI22xp5_ASAP7_75t_L g1883 ( 
.A1(n_1618),
.A2(n_843),
.B1(n_1207),
.B2(n_1096),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1884)
);

AOI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1672),
.A2(n_1391),
.B(n_1220),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1598),
.B(n_1212),
.Y(n_1887)
);

OAI22xp5_ASAP7_75t_L g1888 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1888)
);

OA21x2_ASAP7_75t_L g1889 ( 
.A1(n_1702),
.A2(n_1732),
.B(n_1692),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1672),
.A2(n_1391),
.B(n_1220),
.Y(n_1890)
);

NAND3xp33_ASAP7_75t_L g1891 ( 
.A(n_1598),
.B(n_1207),
.C(n_843),
.Y(n_1891)
);

AOI221xp5_ASAP7_75t_L g1892 ( 
.A1(n_1683),
.A2(n_604),
.B1(n_1164),
.B2(n_685),
.C(n_1079),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1621),
.B(n_1568),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1591),
.B(n_1646),
.Y(n_1894)
);

AOI221xp5_ASAP7_75t_L g1895 ( 
.A1(n_1683),
.A2(n_604),
.B1(n_1164),
.B2(n_685),
.C(n_1079),
.Y(n_1895)
);

AOI22xp33_ASAP7_75t_L g1896 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1591),
.B(n_1646),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1672),
.A2(n_1391),
.B(n_1220),
.Y(n_1899)
);

OAI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1598),
.A2(n_1618),
.B1(n_1199),
.B2(n_1642),
.Y(n_1901)
);

OAI221xp5_ASAP7_75t_L g1902 ( 
.A1(n_1598),
.A2(n_685),
.B1(n_843),
.B2(n_1207),
.C(n_1079),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1672),
.A2(n_1391),
.B(n_1220),
.Y(n_1903)
);

OAI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1598),
.A2(n_1207),
.B(n_685),
.Y(n_1904)
);

BUFx2_ASAP7_75t_L g1905 ( 
.A(n_1599),
.Y(n_1905)
);

AOI211xp5_ASAP7_75t_SL g1906 ( 
.A1(n_1672),
.A2(n_1674),
.B(n_1683),
.C(n_843),
.Y(n_1906)
);

BUFx3_ASAP7_75t_L g1907 ( 
.A(n_1641),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1598),
.A2(n_1618),
.B1(n_1199),
.B2(n_1642),
.Y(n_1908)
);

AOI22xp33_ASAP7_75t_L g1909 ( 
.A1(n_1598),
.A2(n_1618),
.B1(n_1199),
.B2(n_1642),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1591),
.B(n_1646),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1672),
.A2(n_1391),
.B(n_1220),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1621),
.B(n_1568),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1591),
.B(n_1646),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1683),
.A2(n_604),
.B1(n_1164),
.B2(n_685),
.C(n_1079),
.Y(n_1916)
);

AOI22xp33_ASAP7_75t_L g1917 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1629),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1598),
.A2(n_1618),
.B1(n_1199),
.B2(n_1642),
.Y(n_1919)
);

OAI22xp33_ASAP7_75t_L g1920 ( 
.A1(n_1668),
.A2(n_1091),
.B1(n_1674),
.B2(n_1213),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1674),
.A2(n_1091),
.B1(n_1164),
.B2(n_1079),
.Y(n_1921)
);

OAI22xp5_ASAP7_75t_L g1922 ( 
.A1(n_1695),
.A2(n_1392),
.B1(n_1091),
.B2(n_843),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1612),
.Y(n_1923)
);

OAI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1668),
.A2(n_1091),
.B1(n_1674),
.B2(n_1213),
.Y(n_1924)
);

AOI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1683),
.A2(n_604),
.B1(n_1164),
.B2(n_685),
.C(n_1079),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1591),
.B(n_1646),
.Y(n_1926)
);

BUFx2_ASAP7_75t_SL g1927 ( 
.A(n_1762),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1857),
.B(n_1829),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1850),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1852),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1820),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1842),
.Y(n_1932)
);

INVx4_ASAP7_75t_L g1933 ( 
.A(n_1782),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1820),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1829),
.B(n_1779),
.Y(n_1935)
);

BUFx3_ASAP7_75t_L g1936 ( 
.A(n_1762),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1869),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1879),
.B(n_1788),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1829),
.B(n_1889),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1868),
.B(n_1880),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1829),
.B(n_1795),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1791),
.B(n_1883),
.Y(n_1942)
);

AOI221xp5_ASAP7_75t_L g1943 ( 
.A1(n_1863),
.A2(n_1882),
.B1(n_1925),
.B2(n_1895),
.C(n_1916),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1889),
.B(n_1856),
.Y(n_1944)
);

OR2x2_ASAP7_75t_L g1945 ( 
.A(n_1869),
.B(n_1853),
.Y(n_1945)
);

AOI22xp5_ASAP7_75t_L g1946 ( 
.A1(n_1892),
.A2(n_1902),
.B1(n_1877),
.B2(n_1781),
.Y(n_1946)
);

OAI22xp5_ASAP7_75t_L g1947 ( 
.A1(n_1777),
.A2(n_1870),
.B1(n_1896),
.B2(n_1867),
.Y(n_1947)
);

INVx2_ASAP7_75t_SL g1948 ( 
.A(n_1762),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1762),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1796),
.B(n_1840),
.Y(n_1950)
);

OR2x2_ASAP7_75t_L g1951 ( 
.A(n_1855),
.B(n_1849),
.Y(n_1951)
);

INVxp67_ASAP7_75t_L g1952 ( 
.A(n_1785),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1835),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1818),
.B(n_1816),
.Y(n_1954)
);

BUFx2_ASAP7_75t_L g1955 ( 
.A(n_1796),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1818),
.B(n_1816),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1837),
.B(n_1851),
.Y(n_1957)
);

BUFx3_ASAP7_75t_L g1958 ( 
.A(n_1796),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1923),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1837),
.B(n_1796),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1854),
.B(n_1761),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1854),
.B(n_1761),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1831),
.B(n_1764),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1847),
.B(n_1858),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1864),
.B(n_1881),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1803),
.Y(n_1966)
);

AND2x4_ASAP7_75t_L g1967 ( 
.A(n_1786),
.B(n_1769),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1813),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1833),
.B(n_1810),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1792),
.Y(n_1970)
);

INVx3_ASAP7_75t_L g1971 ( 
.A(n_1784),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1766),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1843),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1810),
.B(n_1815),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1844),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1815),
.B(n_1827),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1767),
.B(n_1859),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1858),
.B(n_1805),
.Y(n_1978)
);

BUFx3_ASAP7_75t_L g1979 ( 
.A(n_1771),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1789),
.B(n_1802),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1893),
.B(n_1914),
.Y(n_1981)
);

NOR2xp67_ASAP7_75t_L g1982 ( 
.A(n_1806),
.B(n_1808),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1844),
.Y(n_1983)
);

INVx1_ASAP7_75t_SL g1984 ( 
.A(n_1809),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1836),
.B(n_1774),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1765),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1841),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1887),
.B(n_1823),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1828),
.Y(n_1989)
);

INVxp67_ASAP7_75t_R g1990 ( 
.A(n_1839),
.Y(n_1990)
);

OAI22xp33_ASAP7_75t_L g1991 ( 
.A1(n_1906),
.A2(n_1775),
.B1(n_1924),
.B2(n_1871),
.Y(n_1991)
);

INVx4_ASAP7_75t_L g1992 ( 
.A(n_1782),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1823),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1834),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1846),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1783),
.Y(n_1996)
);

AO21x2_ASAP7_75t_L g1997 ( 
.A1(n_1904),
.A2(n_1885),
.B(n_1890),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1801),
.Y(n_1998)
);

INVxp67_ASAP7_75t_L g1999 ( 
.A(n_1768),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1894),
.B(n_1897),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1801),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1911),
.B(n_1915),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1860),
.B(n_1793),
.Y(n_2003)
);

BUFx3_ASAP7_75t_L g2004 ( 
.A(n_1861),
.Y(n_2004)
);

HB1xp67_ASAP7_75t_L g2005 ( 
.A(n_1826),
.Y(n_2005)
);

HB1xp67_ASAP7_75t_L g2006 ( 
.A(n_1812),
.Y(n_2006)
);

AND2x6_ASAP7_75t_L g2007 ( 
.A(n_1811),
.B(n_1821),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1819),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1819),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1772),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1797),
.B(n_1905),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1772),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1926),
.B(n_1773),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1773),
.B(n_1822),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1860),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1776),
.B(n_1807),
.Y(n_2016)
);

INVx1_ASAP7_75t_SL g2017 ( 
.A(n_1996),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1930),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1959),
.Y(n_2019)
);

AOI22xp33_ASAP7_75t_SL g2020 ( 
.A1(n_1947),
.A2(n_1891),
.B1(n_1763),
.B2(n_1787),
.Y(n_2020)
);

HB1xp67_ASAP7_75t_L g2021 ( 
.A(n_1937),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1943),
.A2(n_1865),
.B1(n_1777),
.B2(n_1870),
.Y(n_2022)
);

AOI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_1943),
.A2(n_1924),
.B1(n_1920),
.B2(n_1871),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1959),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1959),
.Y(n_2025)
);

AOI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1947),
.A2(n_1920),
.B1(n_1888),
.B2(n_1884),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1935),
.B(n_1780),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1946),
.A2(n_1908),
.B1(n_1919),
.B2(n_1901),
.Y(n_2028)
);

NOR4xp25_ASAP7_75t_SL g2029 ( 
.A(n_1953),
.B(n_1838),
.C(n_1862),
.D(n_1874),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_R g2030 ( 
.A(n_1971),
.B(n_1918),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1935),
.B(n_1830),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1965),
.B(n_1793),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1991),
.A2(n_1909),
.B1(n_1921),
.B2(n_1917),
.Y(n_2033)
);

AOI22xp33_ASAP7_75t_L g2034 ( 
.A1(n_1991),
.A2(n_1872),
.B1(n_1921),
.B2(n_1917),
.Y(n_2034)
);

OAI222xp33_ASAP7_75t_L g2035 ( 
.A1(n_1946),
.A2(n_1922),
.B1(n_1912),
.B2(n_1900),
.C1(n_1898),
.C2(n_1873),
.Y(n_2035)
);

OAI31xp33_ASAP7_75t_SL g2036 ( 
.A1(n_1954),
.A2(n_1798),
.A3(n_1814),
.B(n_1778),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1931),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1935),
.B(n_1928),
.Y(n_2038)
);

INVxp67_ASAP7_75t_L g2039 ( 
.A(n_1980),
.Y(n_2039)
);

OR2x2_ASAP7_75t_L g2040 ( 
.A(n_1941),
.B(n_1907),
.Y(n_2040)
);

INVxp67_ASAP7_75t_L g2041 ( 
.A(n_1980),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1937),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1928),
.B(n_1963),
.Y(n_2043)
);

OAI22xp5_ASAP7_75t_L g2044 ( 
.A1(n_1982),
.A2(n_1886),
.B1(n_1910),
.B2(n_1896),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1928),
.B(n_1875),
.Y(n_2045)
);

AOI221xp5_ASAP7_75t_L g2046 ( 
.A1(n_1953),
.A2(n_1867),
.B1(n_1886),
.B2(n_1910),
.C(n_1878),
.Y(n_2046)
);

AO21x2_ASAP7_75t_L g2047 ( 
.A1(n_1972),
.A2(n_1913),
.B(n_1903),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1963),
.B(n_1799),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_SL g2049 ( 
.A1(n_2005),
.A2(n_1878),
.B(n_1872),
.C(n_1790),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1965),
.B(n_1790),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1963),
.B(n_1817),
.Y(n_2051)
);

OR2x2_ASAP7_75t_L g2052 ( 
.A(n_1941),
.B(n_1899),
.Y(n_2052)
);

OR2x2_ASAP7_75t_L g2053 ( 
.A(n_1940),
.B(n_1876),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1945),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1929),
.Y(n_2055)
);

BUFx3_ASAP7_75t_L g2056 ( 
.A(n_1936),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1936),
.Y(n_2057)
);

BUFx3_ASAP7_75t_L g2058 ( 
.A(n_1936),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1981),
.B(n_1800),
.Y(n_2059)
);

AOI33xp33_ASAP7_75t_L g2060 ( 
.A1(n_1954),
.A2(n_1778),
.A3(n_1824),
.B1(n_1832),
.B2(n_1804),
.B3(n_1794),
.Y(n_2060)
);

INVxp67_ASAP7_75t_SL g2061 ( 
.A(n_1952),
.Y(n_2061)
);

NOR3xp33_ASAP7_75t_SL g2062 ( 
.A(n_1998),
.B(n_1825),
.C(n_1804),
.Y(n_2062)
);

AND2x2_ASAP7_75t_L g2063 ( 
.A(n_1973),
.B(n_1961),
.Y(n_2063)
);

BUFx3_ASAP7_75t_L g2064 ( 
.A(n_1949),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1973),
.B(n_1770),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1970),
.Y(n_2066)
);

NAND4xp25_ASAP7_75t_L g2067 ( 
.A(n_1982),
.B(n_1824),
.C(n_1832),
.D(n_1794),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_1940),
.B(n_1782),
.Y(n_2068)
);

OAI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_2005),
.A2(n_1845),
.B(n_1848),
.Y(n_2069)
);

BUFx3_ASAP7_75t_L g2070 ( 
.A(n_1949),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1981),
.B(n_1866),
.Y(n_2071)
);

HB1xp67_ASAP7_75t_L g2072 ( 
.A(n_1945),
.Y(n_2072)
);

NAND3xp33_ASAP7_75t_L g2073 ( 
.A(n_1998),
.B(n_2001),
.C(n_2006),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1970),
.Y(n_2074)
);

NOR4xp25_ASAP7_75t_SL g2075 ( 
.A(n_2001),
.B(n_1955),
.C(n_2009),
.D(n_2008),
.Y(n_2075)
);

BUFx6f_ASAP7_75t_L g2076 ( 
.A(n_1949),
.Y(n_2076)
);

AOI22xp33_ASAP7_75t_SL g2077 ( 
.A1(n_2003),
.A2(n_1954),
.B1(n_1956),
.B2(n_2006),
.Y(n_2077)
);

AND2x4_ASAP7_75t_L g2078 ( 
.A(n_1958),
.B(n_1931),
.Y(n_2078)
);

AOI22xp33_ASAP7_75t_L g2079 ( 
.A1(n_2003),
.A2(n_1942),
.B1(n_1969),
.B2(n_1956),
.Y(n_2079)
);

AO21x2_ASAP7_75t_L g2080 ( 
.A1(n_1972),
.A2(n_1997),
.B(n_1977),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1970),
.Y(n_2081)
);

AOI222xp33_ASAP7_75t_L g2082 ( 
.A1(n_1956),
.A2(n_1969),
.B1(n_1988),
.B2(n_1974),
.C1(n_1976),
.C2(n_1977),
.Y(n_2082)
);

OAI221xp5_ASAP7_75t_L g2083 ( 
.A1(n_1988),
.A2(n_1964),
.B1(n_1938),
.B2(n_1977),
.C(n_1994),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1978),
.B(n_1984),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_1980),
.B(n_1996),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_1973),
.B(n_1961),
.Y(n_2086)
);

BUFx6f_ASAP7_75t_L g2087 ( 
.A(n_1958),
.Y(n_2087)
);

NOR2xp67_ASAP7_75t_L g2088 ( 
.A(n_1978),
.B(n_1934),
.Y(n_2088)
);

OAI33xp33_ASAP7_75t_L g2089 ( 
.A1(n_1964),
.A2(n_2008),
.A3(n_2009),
.B1(n_1952),
.B2(n_2010),
.B3(n_2012),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_1969),
.A2(n_1967),
.B1(n_1974),
.B2(n_1997),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2038),
.B(n_1939),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2038),
.B(n_1939),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2021),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2018),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2080),
.B(n_1939),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2055),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2080),
.B(n_1932),
.Y(n_2097)
);

AND2x4_ASAP7_75t_SL g2098 ( 
.A(n_2076),
.B(n_1950),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2043),
.B(n_1975),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_2043),
.B(n_1975),
.Y(n_2100)
);

AOI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2020),
.A2(n_1997),
.B1(n_1976),
.B2(n_1974),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2063),
.B(n_1961),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_R g2103 ( 
.A(n_2023),
.B(n_1967),
.Y(n_2103)
);

BUFx3_ASAP7_75t_L g2104 ( 
.A(n_2087),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2080),
.B(n_1932),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2084),
.B(n_1986),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2061),
.B(n_1983),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2063),
.B(n_1962),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2019),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2086),
.B(n_2027),
.Y(n_2110)
);

HB1xp67_ASAP7_75t_L g2111 ( 
.A(n_2042),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2019),
.Y(n_2112)
);

AND2x4_ASAP7_75t_SL g2113 ( 
.A(n_2076),
.B(n_1950),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2086),
.B(n_1962),
.Y(n_2114)
);

AOI22xp33_ASAP7_75t_L g2115 ( 
.A1(n_2022),
.A2(n_1997),
.B1(n_1976),
.B2(n_2015),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2054),
.B(n_1983),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2027),
.B(n_1962),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2037),
.B(n_1967),
.Y(n_2118)
);

AND2x2_ASAP7_75t_L g2119 ( 
.A(n_2037),
.B(n_1967),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2024),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2072),
.B(n_1944),
.Y(n_2121)
);

INVx2_ASAP7_75t_SL g2122 ( 
.A(n_2078),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2053),
.B(n_1944),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2053),
.B(n_1944),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2084),
.B(n_2031),
.Y(n_2125)
);

OR2x2_ASAP7_75t_L g2126 ( 
.A(n_2052),
.B(n_1986),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2088),
.B(n_1960),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2088),
.B(n_1960),
.Y(n_2128)
);

AND2x2_ASAP7_75t_L g2129 ( 
.A(n_2045),
.B(n_1960),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2045),
.B(n_2014),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2024),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2025),
.Y(n_2132)
);

INVxp67_ASAP7_75t_L g2133 ( 
.A(n_2073),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2025),
.Y(n_2134)
);

INVx3_ASAP7_75t_L g2135 ( 
.A(n_2078),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2031),
.B(n_2015),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2066),
.Y(n_2137)
);

AND2x2_ASAP7_75t_L g2138 ( 
.A(n_2090),
.B(n_2014),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2065),
.B(n_2014),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2039),
.B(n_2041),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2066),
.B(n_1957),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2052),
.B(n_1987),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2091),
.B(n_2048),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2112),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2112),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2120),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2091),
.B(n_2048),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_2123),
.B(n_2017),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2120),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2131),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2133),
.B(n_2051),
.Y(n_2151)
);

AND2x4_ASAP7_75t_L g2152 ( 
.A(n_2098),
.B(n_2056),
.Y(n_2152)
);

INVx2_ASAP7_75t_SL g2153 ( 
.A(n_2104),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2133),
.B(n_2051),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2131),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2132),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2091),
.B(n_2092),
.Y(n_2157)
);

OAI21xp33_ASAP7_75t_SL g2158 ( 
.A1(n_2101),
.A2(n_2082),
.B(n_2079),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_2136),
.B(n_2083),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2092),
.B(n_2085),
.Y(n_2160)
);

INVxp67_ASAP7_75t_SL g2161 ( 
.A(n_2093),
.Y(n_2161)
);

AOI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_2101),
.A2(n_2028),
.B(n_2036),
.Y(n_2162)
);

HB1xp67_ASAP7_75t_L g2163 ( 
.A(n_2093),
.Y(n_2163)
);

INVx2_ASAP7_75t_L g2164 ( 
.A(n_2094),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2092),
.B(n_2087),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2142),
.B(n_2050),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2142),
.B(n_1999),
.Y(n_2167)
);

INVx2_ASAP7_75t_SL g2168 ( 
.A(n_2104),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2132),
.Y(n_2169)
);

AND2x4_ASAP7_75t_L g2170 ( 
.A(n_2098),
.B(n_2056),
.Y(n_2170)
);

NAND2x1p5_ASAP7_75t_L g2171 ( 
.A(n_2104),
.B(n_1955),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2134),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2123),
.B(n_2040),
.Y(n_2173)
);

AOI222xp33_ASAP7_75t_L g2174 ( 
.A1(n_2115),
.A2(n_2044),
.B1(n_2035),
.B2(n_2033),
.C1(n_2046),
.C2(n_2034),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2094),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2102),
.B(n_2087),
.Y(n_2176)
);

OR2x2_ASAP7_75t_L g2177 ( 
.A(n_2124),
.B(n_2040),
.Y(n_2177)
);

OR2x2_ASAP7_75t_L g2178 ( 
.A(n_2124),
.B(n_2074),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2134),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2094),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_2104),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2109),
.Y(n_2182)
);

OR2x6_ASAP7_75t_L g2183 ( 
.A(n_2107),
.B(n_1927),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2109),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2109),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2107),
.B(n_1999),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_2116),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2111),
.Y(n_2188)
);

NAND2xp5_ASAP7_75t_SL g2189 ( 
.A(n_2115),
.B(n_2073),
.Y(n_2189)
);

INVxp67_ASAP7_75t_L g2190 ( 
.A(n_2125),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2125),
.B(n_2077),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2111),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2094),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2096),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_2126),
.B(n_2074),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2096),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2102),
.B(n_2087),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_2126),
.B(n_2081),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2176),
.B(n_2130),
.Y(n_2199)
);

AOI221xp5_ASAP7_75t_L g2200 ( 
.A1(n_2158),
.A2(n_2189),
.B1(n_2162),
.B2(n_2159),
.C(n_2151),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2144),
.Y(n_2201)
);

NOR3xp33_ASAP7_75t_L g2202 ( 
.A(n_2189),
.B(n_2049),
.C(n_2023),
.Y(n_2202)
);

BUFx2_ASAP7_75t_L g2203 ( 
.A(n_2152),
.Y(n_2203)
);

HB1xp67_ASAP7_75t_L g2204 ( 
.A(n_2163),
.Y(n_2204)
);

AND2x2_ASAP7_75t_L g2205 ( 
.A(n_2176),
.B(n_2130),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2154),
.B(n_2099),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2144),
.Y(n_2207)
);

NOR2xp67_ASAP7_75t_L g2208 ( 
.A(n_2152),
.B(n_2122),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2166),
.B(n_2136),
.Y(n_2209)
);

NAND2xp33_ASAP7_75t_SL g2210 ( 
.A(n_2191),
.B(n_2030),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2187),
.B(n_2141),
.Y(n_2211)
);

NAND4xp25_ASAP7_75t_L g2212 ( 
.A(n_2174),
.B(n_2026),
.C(n_2060),
.D(n_2032),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2156),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2156),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2197),
.B(n_2130),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2145),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2152),
.B(n_2026),
.Y(n_2217)
);

NOR2xp33_ASAP7_75t_L g2218 ( 
.A(n_2190),
.B(n_2071),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2146),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2149),
.Y(n_2220)
);

INVxp67_ASAP7_75t_L g2221 ( 
.A(n_2161),
.Y(n_2221)
);

OR2x2_ASAP7_75t_L g2222 ( 
.A(n_2173),
.B(n_2099),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2173),
.B(n_2100),
.Y(n_2223)
);

OR2x2_ASAP7_75t_L g2224 ( 
.A(n_2177),
.B(n_2100),
.Y(n_2224)
);

NOR2xp67_ASAP7_75t_L g2225 ( 
.A(n_2170),
.B(n_2122),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2167),
.B(n_2186),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_SL g2227 ( 
.A(n_2170),
.B(n_2138),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_SL g2228 ( 
.A(n_2170),
.B(n_2138),
.Y(n_2228)
);

AOI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_2183),
.A2(n_2029),
.B(n_2089),
.Y(n_2229)
);

AND2x2_ASAP7_75t_SL g2230 ( 
.A(n_2197),
.B(n_2103),
.Y(n_2230)
);

OAI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_2171),
.A2(n_2138),
.B(n_2062),
.Y(n_2231)
);

INVx5_ASAP7_75t_L g2232 ( 
.A(n_2183),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2160),
.B(n_2141),
.Y(n_2233)
);

INVxp67_ASAP7_75t_L g2234 ( 
.A(n_2188),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2150),
.Y(n_2235)
);

NAND3xp33_ASAP7_75t_SL g2236 ( 
.A(n_2171),
.B(n_2029),
.C(n_2075),
.Y(n_2236)
);

INVxp67_ASAP7_75t_SL g2237 ( 
.A(n_2164),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2160),
.B(n_2141),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2148),
.B(n_2139),
.Y(n_2239)
);

INVx4_ASAP7_75t_L g2240 ( 
.A(n_2183),
.Y(n_2240)
);

OR2x2_ASAP7_75t_L g2241 ( 
.A(n_2177),
.B(n_2148),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_2171),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2155),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2192),
.B(n_2139),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2143),
.B(n_2139),
.Y(n_2245)
);

OR2x2_ASAP7_75t_L g2246 ( 
.A(n_2178),
.B(n_2126),
.Y(n_2246)
);

INVx2_ASAP7_75t_L g2247 ( 
.A(n_2164),
.Y(n_2247)
);

A2O1A1Ixp33_ASAP7_75t_L g2248 ( 
.A1(n_2153),
.A2(n_2103),
.B(n_1951),
.C(n_1989),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_2143),
.B(n_2129),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2169),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2172),
.Y(n_2251)
);

OR2x2_ASAP7_75t_L g2252 ( 
.A(n_2178),
.B(n_2106),
.Y(n_2252)
);

NOR2x1p5_ASAP7_75t_L g2253 ( 
.A(n_2165),
.B(n_1971),
.Y(n_2253)
);

HB1xp67_ASAP7_75t_L g2254 ( 
.A(n_2182),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2230),
.B(n_2157),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_2202),
.B(n_2147),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2230),
.B(n_2203),
.Y(n_2257)
);

OAI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_2200),
.A2(n_1951),
.B1(n_2183),
.B2(n_1990),
.Y(n_2258)
);

OAI21xp5_ASAP7_75t_SL g2259 ( 
.A1(n_2202),
.A2(n_2067),
.B(n_2069),
.Y(n_2259)
);

INVx2_ASAP7_75t_SL g2260 ( 
.A(n_2253),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2254),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2254),
.Y(n_2262)
);

NOR2xp33_ASAP7_75t_SL g2263 ( 
.A(n_2240),
.B(n_2248),
.Y(n_2263)
);

AND2x2_ASAP7_75t_L g2264 ( 
.A(n_2199),
.B(n_2157),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2205),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2204),
.Y(n_2266)
);

INVxp33_ASAP7_75t_L g2267 ( 
.A(n_2231),
.Y(n_2267)
);

OAI221xp5_ASAP7_75t_SL g2268 ( 
.A1(n_2212),
.A2(n_2095),
.B1(n_2059),
.B2(n_2011),
.C(n_2103),
.Y(n_2268)
);

AOI221xp5_ASAP7_75t_L g2269 ( 
.A1(n_2229),
.A2(n_2095),
.B1(n_2116),
.B2(n_2179),
.C(n_2153),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_2215),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2210),
.A2(n_1990),
.B1(n_2098),
.B2(n_2113),
.Y(n_2271)
);

OAI21xp33_ASAP7_75t_L g2272 ( 
.A1(n_2248),
.A2(n_2013),
.B(n_2095),
.Y(n_2272)
);

NOR2xp33_ASAP7_75t_L g2273 ( 
.A(n_2218),
.B(n_2000),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2217),
.A2(n_2113),
.B1(n_2098),
.B2(n_1950),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_2232),
.B(n_2168),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2201),
.Y(n_2276)
);

AOI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_2227),
.A2(n_2228),
.B1(n_2236),
.B2(n_2217),
.Y(n_2277)
);

AOI322xp5_ASAP7_75t_L g2278 ( 
.A1(n_2227),
.A2(n_2102),
.A3(n_2108),
.B1(n_2114),
.B2(n_2165),
.C1(n_2117),
.C2(n_2127),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2247),
.Y(n_2279)
);

OAI222xp33_ASAP7_75t_L g2280 ( 
.A1(n_2228),
.A2(n_2181),
.B1(n_2168),
.B2(n_2128),
.C1(n_2127),
.C2(n_2068),
.Y(n_2280)
);

OAI22xp5_ASAP7_75t_L g2281 ( 
.A1(n_2232),
.A2(n_2113),
.B1(n_2011),
.B2(n_1989),
.Y(n_2281)
);

NOR2x1_ASAP7_75t_SL g2282 ( 
.A(n_2232),
.B(n_2181),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2204),
.Y(n_2283)
);

OAI221xp5_ASAP7_75t_L g2284 ( 
.A1(n_2240),
.A2(n_2106),
.B1(n_2068),
.B2(n_1994),
.C(n_2121),
.Y(n_2284)
);

AOI222xp33_ASAP7_75t_L g2285 ( 
.A1(n_2221),
.A2(n_2013),
.B1(n_2016),
.B2(n_1989),
.C1(n_1993),
.C2(n_2010),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2218),
.B(n_2147),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2209),
.B(n_2108),
.Y(n_2287)
);

INVx1_ASAP7_75t_SL g2288 ( 
.A(n_2241),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2207),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2213),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2214),
.Y(n_2291)
);

OAI322xp33_ASAP7_75t_L g2292 ( 
.A1(n_2221),
.A2(n_2097),
.A3(n_2105),
.B1(n_2106),
.B2(n_2184),
.C1(n_2185),
.C2(n_2121),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2208),
.B(n_2225),
.Y(n_2293)
);

NAND3xp33_ASAP7_75t_L g2294 ( 
.A(n_2234),
.B(n_2012),
.C(n_1993),
.Y(n_2294)
);

OAI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2232),
.A2(n_2113),
.B1(n_2127),
.B2(n_2128),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2216),
.Y(n_2296)
);

OA21x2_ASAP7_75t_SL g2297 ( 
.A1(n_2267),
.A2(n_2226),
.B(n_2239),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_2257),
.B(n_2255),
.Y(n_2298)
);

AOI221xp5_ASAP7_75t_L g2299 ( 
.A1(n_2267),
.A2(n_2234),
.B1(n_2251),
.B2(n_2250),
.C(n_2219),
.Y(n_2299)
);

OAI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_2277),
.A2(n_2242),
.B1(n_2206),
.B2(n_2244),
.C(n_2211),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2288),
.B(n_2249),
.Y(n_2301)
);

AOI221xp5_ASAP7_75t_L g2302 ( 
.A1(n_2268),
.A2(n_2220),
.B1(n_2235),
.B2(n_2243),
.C(n_2237),
.Y(n_2302)
);

INVx1_ASAP7_75t_SL g2303 ( 
.A(n_2257),
.Y(n_2303)
);

OAI22xp33_ASAP7_75t_SL g2304 ( 
.A1(n_2263),
.A2(n_2224),
.B1(n_2222),
.B2(n_2223),
.Y(n_2304)
);

A2O1A1Ixp33_ASAP7_75t_L g2305 ( 
.A1(n_2269),
.A2(n_2272),
.B(n_2259),
.C(n_2258),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2255),
.B(n_2245),
.Y(n_2306)
);

OAI21xp33_ASAP7_75t_SL g2307 ( 
.A1(n_2275),
.A2(n_2238),
.B(n_2233),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2262),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2262),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2271),
.A2(n_2128),
.B1(n_2252),
.B2(n_2114),
.Y(n_2310)
);

AOI221xp5_ASAP7_75t_L g2311 ( 
.A1(n_2292),
.A2(n_2237),
.B1(n_2247),
.B2(n_2246),
.C(n_2196),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2256),
.B(n_2108),
.Y(n_2312)
);

OAI21xp33_ASAP7_75t_L g2313 ( 
.A1(n_2278),
.A2(n_2013),
.B(n_1985),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2276),
.Y(n_2314)
);

INVxp67_ASAP7_75t_L g2315 ( 
.A(n_2266),
.Y(n_2315)
);

OAI221xp5_ASAP7_75t_L g2316 ( 
.A1(n_2260),
.A2(n_2122),
.B1(n_2097),
.B2(n_2105),
.C(n_2194),
.Y(n_2316)
);

OAI22xp5_ASAP7_75t_L g2317 ( 
.A1(n_2274),
.A2(n_2114),
.B1(n_2135),
.B2(n_2117),
.Y(n_2317)
);

OAI21xp33_ASAP7_75t_SL g2318 ( 
.A1(n_2275),
.A2(n_2129),
.B(n_2117),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2276),
.Y(n_2319)
);

AOI22xp5_ASAP7_75t_L g2320 ( 
.A1(n_2260),
.A2(n_1950),
.B1(n_2007),
.B2(n_1985),
.Y(n_2320)
);

OR2x2_ASAP7_75t_L g2321 ( 
.A(n_2286),
.B(n_2195),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_SL g2322 ( 
.A(n_2294),
.B(n_2087),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2291),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2291),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_2273),
.B(n_2129),
.Y(n_2325)
);

INVxp67_ASAP7_75t_L g2326 ( 
.A(n_2283),
.Y(n_2326)
);

INVxp67_ASAP7_75t_SL g2327 ( 
.A(n_2282),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2303),
.B(n_2285),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2314),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2298),
.B(n_2293),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2308),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2309),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2306),
.B(n_2293),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2319),
.Y(n_2334)
);

AOI32xp33_ASAP7_75t_L g2335 ( 
.A1(n_2297),
.A2(n_2281),
.A3(n_2295),
.B1(n_2261),
.B2(n_2270),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2315),
.B(n_2296),
.Y(n_2336)
);

NAND3xp33_ASAP7_75t_L g2337 ( 
.A(n_2305),
.B(n_2299),
.C(n_2302),
.Y(n_2337)
);

NOR3xp33_ASAP7_75t_SL g2338 ( 
.A(n_2307),
.B(n_2280),
.C(n_2284),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2323),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_2315),
.B(n_2265),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2327),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_2304),
.B(n_2265),
.Y(n_2342)
);

NOR4xp75_ASAP7_75t_L g2343 ( 
.A(n_2300),
.B(n_2282),
.C(n_2287),
.D(n_1971),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2326),
.B(n_2270),
.Y(n_2344)
);

NAND2xp33_ASAP7_75t_L g2345 ( 
.A(n_2301),
.B(n_2289),
.Y(n_2345)
);

INVx1_ASAP7_75t_SL g2346 ( 
.A(n_2322),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2324),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2327),
.B(n_2264),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2326),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2321),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2312),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2330),
.B(n_2264),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2348),
.B(n_2322),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2347),
.Y(n_2354)
);

NAND4xp75_ASAP7_75t_L g2355 ( 
.A(n_2338),
.B(n_2318),
.C(n_2311),
.D(n_2290),
.Y(n_2355)
);

CKINVDCx5p33_ASAP7_75t_R g2356 ( 
.A(n_2341),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2341),
.B(n_2313),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2347),
.Y(n_2358)
);

AOI211xp5_ASAP7_75t_L g2359 ( 
.A1(n_2337),
.A2(n_2310),
.B(n_2317),
.C(n_2316),
.Y(n_2359)
);

OAI221xp5_ASAP7_75t_L g2360 ( 
.A1(n_2335),
.A2(n_2320),
.B1(n_2325),
.B2(n_2279),
.C(n_1971),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2347),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2348),
.Y(n_2362)
);

NAND4xp25_ASAP7_75t_L g2363 ( 
.A(n_2328),
.B(n_2340),
.C(n_2344),
.D(n_2342),
.Y(n_2363)
);

NOR3xp33_ASAP7_75t_L g2364 ( 
.A(n_2349),
.B(n_2279),
.C(n_2016),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2330),
.B(n_2000),
.Y(n_2365)
);

OAI21xp33_ASAP7_75t_L g2366 ( 
.A1(n_2333),
.A2(n_2016),
.B(n_2097),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2362),
.B(n_2333),
.Y(n_2367)
);

OAI211xp5_ASAP7_75t_SL g2368 ( 
.A1(n_2359),
.A2(n_2345),
.B(n_2336),
.C(n_2350),
.Y(n_2368)
);

NAND2xp33_ASAP7_75t_R g2369 ( 
.A(n_2356),
.B(n_2350),
.Y(n_2369)
);

AOI221xp5_ASAP7_75t_SL g2370 ( 
.A1(n_2363),
.A2(n_2345),
.B1(n_2346),
.B2(n_2351),
.C(n_2331),
.Y(n_2370)
);

AOI211x1_ASAP7_75t_L g2371 ( 
.A1(n_2360),
.A2(n_2351),
.B(n_2331),
.C(n_2332),
.Y(n_2371)
);

AOI222xp33_ASAP7_75t_L g2372 ( 
.A1(n_2357),
.A2(n_2332),
.B1(n_2339),
.B2(n_2329),
.C1(n_2334),
.C2(n_2343),
.Y(n_2372)
);

AOI221xp5_ASAP7_75t_L g2373 ( 
.A1(n_2357),
.A2(n_2334),
.B1(n_2193),
.B2(n_2180),
.C(n_2175),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2355),
.A2(n_2135),
.B1(n_2105),
.B2(n_2195),
.Y(n_2374)
);

OAI211xp5_ASAP7_75t_SL g2375 ( 
.A1(n_2353),
.A2(n_2135),
.B(n_2193),
.C(n_2180),
.Y(n_2375)
);

A2O1A1Ixp33_ASAP7_75t_L g2376 ( 
.A1(n_2352),
.A2(n_2070),
.B(n_2056),
.C(n_2057),
.Y(n_2376)
);

AOI221xp5_ASAP7_75t_L g2377 ( 
.A1(n_2364),
.A2(n_2361),
.B1(n_2358),
.B2(n_2354),
.C(n_2366),
.Y(n_2377)
);

OAI22xp33_ASAP7_75t_L g2378 ( 
.A1(n_2365),
.A2(n_2087),
.B1(n_2076),
.B2(n_2135),
.Y(n_2378)
);

A2O1A1Ixp33_ASAP7_75t_L g2379 ( 
.A1(n_2359),
.A2(n_2070),
.B(n_2058),
.C(n_2057),
.Y(n_2379)
);

AND2x4_ASAP7_75t_L g2380 ( 
.A(n_2367),
.B(n_2379),
.Y(n_2380)
);

NOR2x1_ASAP7_75t_L g2381 ( 
.A(n_2368),
.B(n_2175),
.Y(n_2381)
);

AOI21xp33_ASAP7_75t_SL g2382 ( 
.A1(n_2372),
.A2(n_2198),
.B(n_1948),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_2374),
.A2(n_2369),
.B1(n_2370),
.B2(n_2377),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2376),
.B(n_2198),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2371),
.B(n_2373),
.Y(n_2385)
);

NAND2xp33_ASAP7_75t_SL g2386 ( 
.A(n_2375),
.B(n_2076),
.Y(n_2386)
);

NOR2xp33_ASAP7_75t_R g2387 ( 
.A(n_2378),
.B(n_1979),
.Y(n_2387)
);

AOI221xp5_ASAP7_75t_L g2388 ( 
.A1(n_2382),
.A2(n_2076),
.B1(n_1995),
.B2(n_2047),
.C(n_2118),
.Y(n_2388)
);

NOR4xp75_ASAP7_75t_L g2389 ( 
.A(n_2385),
.B(n_2135),
.C(n_2119),
.D(n_2118),
.Y(n_2389)
);

NOR3xp33_ASAP7_75t_L g2390 ( 
.A(n_2383),
.B(n_1933),
.C(n_1992),
.Y(n_2390)
);

NOR3xp33_ASAP7_75t_L g2391 ( 
.A(n_2380),
.B(n_1933),
.C(n_1992),
.Y(n_2391)
);

AND2x2_ASAP7_75t_L g2392 ( 
.A(n_2381),
.B(n_2384),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2387),
.B(n_2110),
.Y(n_2393)
);

NOR3xp33_ASAP7_75t_SL g2394 ( 
.A(n_2386),
.B(n_1995),
.C(n_1987),
.Y(n_2394)
);

INVx1_ASAP7_75t_SL g2395 ( 
.A(n_2380),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2395),
.B(n_2000),
.Y(n_2396)
);

AOI221xp5_ASAP7_75t_L g2397 ( 
.A1(n_2390),
.A2(n_2076),
.B1(n_1979),
.B2(n_2004),
.C(n_2140),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2392),
.B(n_2110),
.Y(n_2398)
);

NAND3xp33_ASAP7_75t_L g2399 ( 
.A(n_2391),
.B(n_1979),
.C(n_2004),
.Y(n_2399)
);

NAND3xp33_ASAP7_75t_SL g2400 ( 
.A(n_2389),
.B(n_2002),
.C(n_1933),
.Y(n_2400)
);

NOR3xp33_ASAP7_75t_SL g2401 ( 
.A(n_2388),
.B(n_1968),
.C(n_1966),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2398),
.Y(n_2402)
);

NOR3xp33_ASAP7_75t_L g2403 ( 
.A(n_2397),
.B(n_2393),
.C(n_2394),
.Y(n_2403)
);

INVxp67_ASAP7_75t_L g2404 ( 
.A(n_2396),
.Y(n_2404)
);

INVx1_ASAP7_75t_SL g2405 ( 
.A(n_2399),
.Y(n_2405)
);

AOI22xp5_ASAP7_75t_L g2406 ( 
.A1(n_2402),
.A2(n_2403),
.B1(n_2405),
.B2(n_2404),
.Y(n_2406)
);

AO21x2_ASAP7_75t_L g2407 ( 
.A1(n_2406),
.A2(n_2400),
.B(n_2401),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2407),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2407),
.Y(n_2409)
);

AOI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_2408),
.A2(n_2002),
.B(n_2140),
.Y(n_2410)
);

XNOR2xp5_ASAP7_75t_L g2411 ( 
.A(n_2409),
.B(n_2004),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2411),
.A2(n_2002),
.B(n_2140),
.Y(n_2412)
);

AOI222xp33_ASAP7_75t_L g2413 ( 
.A1(n_2410),
.A2(n_2058),
.B1(n_2070),
.B2(n_2057),
.C1(n_2064),
.C2(n_2110),
.Y(n_2413)
);

INVxp67_ASAP7_75t_SL g2414 ( 
.A(n_2412),
.Y(n_2414)
);

AOI221xp5_ASAP7_75t_L g2415 ( 
.A1(n_2414),
.A2(n_2413),
.B1(n_2058),
.B2(n_2064),
.C(n_2137),
.Y(n_2415)
);

AOI211xp5_ASAP7_75t_L g2416 ( 
.A1(n_2415),
.A2(n_1948),
.B(n_2064),
.C(n_2118),
.Y(n_2416)
);


endmodule