module fake_jpeg_8448_n_112 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_112);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

OR2x2_ASAP7_75t_SL g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_3),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_24),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_SL g42 ( 
.A(n_26),
.Y(n_42)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_12),
.B1(n_16),
.B2(n_22),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_49),
.B1(n_25),
.B2(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_50),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_12),
.B1(n_16),
.B2(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_20),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_44),
.A2(n_30),
.B(n_34),
.C(n_25),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_55),
.B1(n_56),
.B2(n_39),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_58),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_37),
.C(n_41),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_63),
.Y(n_73)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_11),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_6),
.C(n_8),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_21),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_18),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_18),
.C(n_10),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_10),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_48),
.B(n_38),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_73),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_64),
.B1(n_18),
.B2(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_56),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_80),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_55),
.Y(n_80)
);

XOR2x2_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_18),
.Y(n_81)
);

NAND2xp67_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_86),
.B(n_73),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_94),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_83),
.B1(n_78),
.B2(n_68),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_87),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_97),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_67),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_96),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_92),
.Y(n_103)
);

NOR2xp67_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_101),
.B(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_101),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_107),
.B(n_106),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_108),
.B(n_67),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_64),
.Y(n_112)
);


endmodule