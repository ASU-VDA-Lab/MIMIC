module fake_jpeg_2003_n_607 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_607);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_607;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_17),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_57),
.B(n_64),
.Y(n_136)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_76),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_47),
.B(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_68),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_69),
.B(n_84),
.Y(n_177)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_72),
.Y(n_162)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_74),
.Y(n_172)
);

CKINVDCx6p67_ASAP7_75t_R g75 ( 
.A(n_21),
.Y(n_75)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_75),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_37),
.B(n_9),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

BUFx12f_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_95),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_82),
.Y(n_141)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_39),
.B(n_9),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_39),
.A2(n_10),
.B(n_18),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_85),
.B(n_89),
.Y(n_168)
);

BUFx2_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_87),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

BUFx2_ASAP7_75t_SL g123 ( 
.A(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_43),
.B(n_10),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_90),
.Y(n_133)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_101),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_50),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_44),
.A2(n_8),
.B1(n_18),
.B2(n_17),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_26),
.B1(n_40),
.B2(n_34),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_8),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_45),
.B(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_77),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_106),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_19),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_40),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_79),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_115),
.A2(n_119),
.B1(n_129),
.B2(n_134),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_118),
.B(n_130),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_75),
.A2(n_24),
.B1(n_29),
.B2(n_48),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_51),
.B1(n_33),
.B2(n_29),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_46),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_132),
.B(n_135),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_70),
.B(n_26),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_55),
.A2(n_33),
.B1(n_49),
.B2(n_38),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_140),
.A2(n_142),
.B1(n_146),
.B2(n_155),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_65),
.A2(n_29),
.B1(n_32),
.B2(n_41),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_100),
.A2(n_29),
.B1(n_33),
.B2(n_53),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_78),
.A2(n_32),
.B1(n_41),
.B2(n_49),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_83),
.A2(n_51),
.B1(n_53),
.B2(n_38),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_157),
.A2(n_164),
.B1(n_41),
.B2(n_32),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_109),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_160),
.B(n_165),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_87),
.A2(n_32),
.B1(n_41),
.B2(n_49),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_34),
.Y(n_165)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_91),
.C(n_73),
.Y(n_191)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_178),
.B(n_192),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_112),
.B(n_63),
.Y(n_180)
);

OAI21xp33_ASAP7_75t_L g253 ( 
.A1(n_180),
.A2(n_191),
.B(n_206),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_121),
.B(n_68),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_181),
.B(n_204),
.Y(n_244)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_182),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_185),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_122),
.A2(n_63),
.B(n_86),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_186),
.A2(n_213),
.B(n_214),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_187),
.B(n_196),
.Y(n_246)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_138),
.Y(n_188)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_80),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_193),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_194),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_67),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_195),
.B(n_209),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_197),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_198),
.A2(n_90),
.B1(n_158),
.B2(n_144),
.Y(n_257)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_131),
.Y(n_199)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_200),
.Y(n_287)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_143),
.B(n_61),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_202),
.Y(n_249)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_113),
.B(n_104),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_112),
.B(n_58),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_141),
.B(n_48),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_122),
.B(n_81),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_210),
.B(n_215),
.Y(n_272)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_211),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_124),
.A2(n_96),
.B1(n_105),
.B2(n_111),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_212),
.A2(n_235),
.B1(n_1),
.B2(n_2),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_115),
.A2(n_119),
.B(n_136),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_120),
.A2(n_98),
.B(n_88),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_159),
.B(n_48),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_0),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_216),
.B(n_220),
.Y(n_270)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_114),
.Y(n_217)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_217),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_218),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_126),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_0),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_147),
.B(n_88),
.C(n_108),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_221),
.B(n_127),
.C(n_169),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g222 ( 
.A1(n_151),
.A2(n_98),
.B(n_71),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_223),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_174),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_114),
.Y(n_224)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_173),
.B(n_97),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_231),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_150),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_228),
.Y(n_280)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_227),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_140),
.B(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_31),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_229),
.B(n_241),
.Y(n_292)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_153),
.B(n_93),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_156),
.Y(n_232)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_232),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_176),
.A2(n_110),
.B1(n_94),
.B2(n_53),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_133),
.Y(n_236)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_117),
.Y(n_237)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_139),
.B(n_1),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_142),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_127),
.A2(n_60),
.B(n_27),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_31),
.Y(n_263)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_149),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_240),
.Y(n_265)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_123),
.A2(n_35),
.B(n_27),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_176),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_243),
.B(n_249),
.Y(n_314)
);

OAI32xp33_ASAP7_75t_L g251 ( 
.A1(n_178),
.A2(n_155),
.A3(n_164),
.B1(n_163),
.B2(n_145),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_251),
.B(n_255),
.Y(n_351)
);

OAI32xp33_ASAP7_75t_L g256 ( 
.A1(n_192),
.A2(n_163),
.A3(n_145),
.B1(n_158),
.B2(n_139),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_214),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_257),
.A2(n_290),
.B1(n_199),
.B2(n_184),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_263),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_228),
.A2(n_144),
.B1(n_169),
.B2(n_149),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_267),
.A2(n_274),
.B1(n_239),
.B2(n_180),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_233),
.A2(n_53),
.B1(n_38),
.B2(n_31),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_271),
.A2(n_278),
.B1(n_285),
.B2(n_295),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_L g274 ( 
.A1(n_213),
.A2(n_38),
.B1(n_35),
.B2(n_27),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_208),
.A2(n_238),
.B1(n_209),
.B2(n_220),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_35),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_281),
.B(n_283),
.C(n_221),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_207),
.B(n_35),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_216),
.A2(n_35),
.B1(n_11),
.B2(n_12),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_200),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_180),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_226),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_189),
.B(n_18),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_297),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_183),
.B(n_196),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_190),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_186),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_300),
.B(n_294),
.Y(n_385)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_250),
.Y(n_301)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_302),
.A2(n_346),
.B1(n_347),
.B2(n_350),
.Y(n_377)
);

OAI21xp33_ASAP7_75t_SL g359 ( 
.A1(n_303),
.A2(n_325),
.B(n_275),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_278),
.B1(n_258),
.B2(n_263),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_304),
.A2(n_311),
.B1(n_318),
.B2(n_335),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_286),
.Y(n_305)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_305),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_248),
.B(n_206),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_308),
.B(n_314),
.Y(n_373)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_309),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_202),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_310),
.B(n_312),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_280),
.A2(n_224),
.B1(n_236),
.B2(n_217),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_270),
.B(n_202),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g313 ( 
.A(n_246),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_313),
.B(n_323),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_315),
.B(n_269),
.Y(n_394)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_317),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_258),
.A2(n_230),
.B1(n_188),
.B2(n_179),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_276),
.A2(n_179),
.B(n_206),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_319),
.A2(n_330),
.B(n_345),
.Y(n_388)
);

INVx8_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_321),
.Y(n_376)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_322),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_287),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_248),
.B(n_193),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_326),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_264),
.B(n_182),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_247),
.Y(n_327)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_327),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_197),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_337),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_263),
.A2(n_187),
.B(n_184),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_268),
.B(n_275),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_272),
.A2(n_211),
.B(n_234),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_244),
.B(n_185),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_266),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_334),
.Y(n_380)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_247),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_243),
.A2(n_194),
.B1(n_237),
.B2(n_232),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_201),
.C(n_203),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_341),
.C(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_245),
.B(n_283),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_255),
.B(n_256),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_342),
.Y(n_367)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_262),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_339),
.B(n_340),
.Y(n_387)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_262),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_259),
.C(n_277),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_295),
.B(n_205),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_273),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_344),
.Y(n_375)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_253),
.A2(n_232),
.B(n_219),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_271),
.A2(n_240),
.B1(n_227),
.B2(n_242),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_251),
.A2(n_205),
.B1(n_2),
.B2(n_3),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_285),
.A2(n_205),
.B1(n_7),
.B2(n_11),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_348),
.A2(n_265),
.B1(n_288),
.B2(n_261),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_259),
.B(n_18),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_352),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_265),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_268),
.B(n_7),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_352),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_356),
.B(n_363),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_359),
.A2(n_365),
.B1(n_381),
.B2(n_345),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_360),
.A2(n_372),
.B(n_374),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_361),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_314),
.B(n_277),
.C(n_261),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_362),
.B(n_378),
.C(n_394),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_349),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_337),
.B(n_260),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_364),
.B(n_386),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_317),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_370),
.B(n_326),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_304),
.A2(n_252),
.B(n_260),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_303),
.A2(n_252),
.B(n_291),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_315),
.B(n_254),
.C(n_293),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_338),
.A2(n_298),
.B1(n_266),
.B2(n_282),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_330),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_382),
.B(n_343),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g386 ( 
.A(n_310),
.B(n_282),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_351),
.A2(n_298),
.B1(n_296),
.B2(n_279),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_390),
.A2(n_393),
.B1(n_335),
.B2(n_316),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_254),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_309),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_351),
.A2(n_291),
.B1(n_269),
.B2(n_293),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_294),
.C(n_286),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_395),
.B(n_397),
.C(n_398),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_336),
.B(n_284),
.C(n_4),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_312),
.B(n_284),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_307),
.A2(n_3),
.B(n_4),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_350),
.B(n_301),
.Y(n_429)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_401),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_373),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_425),
.Y(n_440)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_387),
.Y(n_404)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_405),
.B(n_411),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_406),
.A2(n_407),
.B1(n_427),
.B2(n_428),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_381),
.A2(n_391),
.B1(n_377),
.B2(n_374),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_387),
.Y(n_408)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_380),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_355),
.B(n_328),
.Y(n_412)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_375),
.Y(n_413)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g470 ( 
.A(n_414),
.Y(n_470)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_415),
.B(n_416),
.Y(n_443)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_369),
.B(n_333),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_417),
.B(n_370),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_377),
.A2(n_307),
.B1(n_302),
.B2(n_306),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_418),
.A2(n_423),
.B1(n_430),
.B2(n_390),
.Y(n_457)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_419),
.B(n_426),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_355),
.B(n_308),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_422),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_367),
.A2(n_306),
.B1(n_300),
.B2(n_318),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_378),
.B(n_341),
.C(n_319),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_420),
.C(n_403),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_373),
.B(n_329),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_380),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_358),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_391),
.A2(n_347),
.B1(n_346),
.B2(n_342),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_429),
.A2(n_431),
.B1(n_432),
.B2(n_433),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_367),
.A2(n_311),
.B1(n_348),
.B2(n_327),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_358),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_382),
.A2(n_322),
.B1(n_334),
.B2(n_323),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_434),
.A2(n_437),
.B1(n_438),
.B2(n_439),
.Y(n_463)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_372),
.A2(n_344),
.B1(n_340),
.B2(n_339),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_364),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_444),
.B(n_460),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_445),
.B(n_415),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_449),
.B(n_451),
.C(n_453),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_361),
.C(n_398),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_362),
.C(n_395),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_402),
.B(n_353),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_454),
.B(n_429),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_386),
.C(n_353),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_455),
.B(n_458),
.C(n_469),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_407),
.A2(n_406),
.B1(n_428),
.B2(n_413),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_456),
.A2(n_459),
.B1(n_461),
.B2(n_464),
.Y(n_492)
);

AO21x1_ASAP7_75t_L g495 ( 
.A1(n_457),
.A2(n_466),
.B(n_409),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_410),
.B(n_357),
.C(n_393),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_414),
.A2(n_357),
.B1(n_376),
.B2(n_379),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_410),
.B(n_379),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_422),
.A2(n_363),
.B1(n_360),
.B2(n_392),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_412),
.A2(n_356),
.B1(n_389),
.B2(n_368),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_427),
.A2(n_388),
.B1(n_365),
.B2(n_389),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_388),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_408),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_423),
.A2(n_354),
.B1(n_368),
.B2(n_383),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_468),
.A2(n_471),
.B1(n_474),
.B2(n_416),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_418),
.B(n_397),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_434),
.A2(n_354),
.B1(n_383),
.B2(n_399),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_332),
.C(n_366),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_440),
.C(n_444),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_435),
.A2(n_366),
.B1(n_320),
.B2(n_305),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_433),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_476),
.B(n_487),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_473),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_490),
.Y(n_517)
);

MAJx2_ASAP7_75t_L g526 ( 
.A(n_479),
.B(n_500),
.C(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_481),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_483),
.B(n_499),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_426),
.C(n_411),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_484),
.B(n_489),
.C(n_493),
.Y(n_511)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_443),
.Y(n_485)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_485),
.Y(n_531)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_452),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_488),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_436),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_449),
.B(n_436),
.C(n_430),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_474),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_441),
.B(n_405),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_491),
.B(n_494),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_453),
.B(n_401),
.C(n_409),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_439),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_495),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_455),
.B(n_438),
.C(n_400),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_496),
.B(n_505),
.C(n_472),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_497),
.A2(n_498),
.B1(n_475),
.B2(n_13),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_440),
.B(n_437),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_447),
.B(n_441),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_501),
.A2(n_503),
.B(n_471),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_432),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_502),
.B(n_504),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_442),
.A2(n_431),
.B(n_419),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_454),
.B(n_320),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_469),
.B(n_4),
.C(n_5),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_14),
.Y(n_506)
);

OA21x2_ASAP7_75t_SL g507 ( 
.A1(n_503),
.A2(n_465),
.B(n_472),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_527),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g508 ( 
.A(n_479),
.B(n_467),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_SL g534 ( 
.A(n_508),
.B(n_525),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_456),
.B1(n_468),
.B2(n_446),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_510),
.A2(n_515),
.B1(n_495),
.B2(n_493),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_478),
.A2(n_446),
.B1(n_470),
.B2(n_448),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_520),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_490),
.A2(n_457),
.B1(n_463),
.B2(n_470),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_483),
.B(n_458),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_519),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_480),
.B(n_462),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_448),
.Y(n_521)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_521),
.Y(n_536)
);

INVx13_ASAP7_75t_L g522 ( 
.A(n_498),
.Y(n_522)
);

INVxp33_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_524),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_500),
.B(n_499),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_477),
.B(n_475),
.C(n_461),
.Y(n_527)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_528),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_480),
.B(n_13),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_506),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_477),
.C(n_484),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_540),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_539),
.A2(n_517),
.B1(n_515),
.B2(n_510),
.Y(n_567)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_523),
.Y(n_541)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_541),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_511),
.B(n_513),
.C(n_516),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_542),
.B(n_546),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_509),
.A2(n_492),
.B(n_489),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_543),
.A2(n_509),
.B(n_524),
.Y(n_555)
);

CKINVDCx14_ASAP7_75t_R g546 ( 
.A(n_512),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_530),
.B(n_531),
.Y(n_548)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_548),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_513),
.B(n_496),
.C(n_482),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_549),
.B(n_550),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_482),
.C(n_505),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_520),
.B(n_4),
.C(n_5),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_551),
.B(n_552),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_519),
.B(n_5),
.C(n_6),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_530),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_531),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_534),
.B(n_525),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_560),
.Y(n_572)
);

AO21x1_ASAP7_75t_L g575 ( 
.A1(n_555),
.A2(n_533),
.B(n_561),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_557),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_537),
.B(n_518),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_558),
.B(n_561),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_521),
.Y(n_559)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_559),
.Y(n_578)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_508),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_533),
.A2(n_517),
.B1(n_522),
.B2(n_529),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_535),
.B(n_544),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_563),
.B(n_567),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_544),
.B(n_514),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_568),
.B(n_571),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_SL g570 ( 
.A(n_542),
.B(n_532),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_570),
.A2(n_543),
.B(n_548),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_526),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_564),
.B(n_550),
.C(n_549),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_573),
.B(n_580),
.Y(n_589)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_575),
.A2(n_568),
.B(n_571),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_538),
.Y(n_580)
);

AOI21xp33_ASAP7_75t_L g592 ( 
.A1(n_581),
.A2(n_554),
.B(n_526),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_562),
.B(n_547),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_582),
.B(n_583),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_569),
.B(n_536),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_559),
.B(n_547),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g594 ( 
.A1(n_584),
.A2(n_585),
.B(n_540),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g585 ( 
.A1(n_555),
.A2(n_552),
.B(n_534),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_579),
.B(n_567),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_586),
.B(n_588),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_587),
.A2(n_590),
.B(n_592),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_579),
.B(n_563),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_573),
.B(n_556),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_577),
.A2(n_566),
.B1(n_551),
.B2(n_560),
.Y(n_591)
);

AO221x1_ASAP7_75t_L g597 ( 
.A1(n_591),
.A2(n_575),
.B1(n_576),
.B2(n_572),
.C(n_578),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_594),
.B(n_581),
.C(n_585),
.Y(n_595)
);

NOR2x1_ASAP7_75t_L g600 ( 
.A(n_595),
.B(n_597),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_589),
.A2(n_574),
.B(n_572),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_599),
.B(n_588),
.C(n_586),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_601),
.A2(n_598),
.B1(n_593),
.B2(n_13),
.Y(n_603)
);

BUFx24_ASAP7_75t_SL g602 ( 
.A(n_596),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g604 ( 
.A(n_602),
.B(n_13),
.C(n_6),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_603),
.A2(n_604),
.B(n_600),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_605),
.B(n_6),
.C(n_596),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_606),
.B(n_6),
.Y(n_607)
);


endmodule