module real_aes_2992_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_832, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_832;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_649;
wire n_397;
wire n_162;
wire n_293;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g230 ( .A(n_0), .B(n_167), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_1), .B(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g139 ( .A(n_2), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_3), .B(n_143), .Y(n_188) );
NAND2xp33_ASAP7_75t_SL g250 ( .A(n_4), .B(n_149), .Y(n_250) );
INVx1_ASAP7_75t_L g242 ( .A(n_5), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_6), .B(n_193), .Y(n_460) );
INVx1_ASAP7_75t_L g504 ( .A(n_7), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_8), .Y(n_106) );
AND2x2_ASAP7_75t_L g186 ( .A(n_9), .B(n_172), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_10), .Y(n_496) );
INVx2_ASAP7_75t_L g131 ( .A(n_11), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g469 ( .A(n_13), .Y(n_469) );
AOI221x1_ASAP7_75t_L g245 ( .A1(n_14), .A2(n_151), .B1(n_246), .B2(n_248), .C(n_249), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_15), .B(n_143), .Y(n_210) );
INVx1_ASAP7_75t_L g114 ( .A(n_16), .Y(n_114) );
INVx1_ASAP7_75t_L g467 ( .A(n_17), .Y(n_467) );
INVx1_ASAP7_75t_SL g563 ( .A(n_18), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_19), .B(n_144), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_20), .A2(n_151), .B(n_190), .Y(n_189) );
AOI221xp5_ASAP7_75t_SL g219 ( .A1(n_21), .A2(n_38), .B1(n_143), .B2(n_151), .C(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_22), .B(n_167), .Y(n_191) );
AOI33xp33_ASAP7_75t_L g513 ( .A1(n_23), .A2(n_50), .A3(n_136), .B1(n_156), .B2(n_514), .B3(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g490 ( .A(n_24), .Y(n_490) );
INVx1_ASAP7_75t_L g117 ( .A(n_25), .Y(n_117) );
OA21x2_ASAP7_75t_L g130 ( .A1(n_26), .A2(n_88), .B(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g173 ( .A(n_26), .B(n_88), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_27), .B(n_165), .Y(n_214) );
INVxp67_ASAP7_75t_L g244 ( .A(n_28), .Y(n_244) );
AND2x2_ASAP7_75t_L g183 ( .A(n_29), .B(n_171), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_30), .B(n_134), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_31), .A2(n_151), .B(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_32), .B(n_165), .Y(n_221) );
AOI222xp33_ASAP7_75t_SL g99 ( .A1(n_33), .A2(n_100), .B1(n_116), .B2(n_806), .C1(n_808), .C2(n_824), .Y(n_99) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_33), .A2(n_49), .B1(n_649), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g816 ( .A(n_33), .Y(n_816) );
AND2x2_ASAP7_75t_L g141 ( .A(n_34), .B(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g149 ( .A(n_34), .B(n_139), .Y(n_149) );
INVx1_ASAP7_75t_L g155 ( .A(n_34), .Y(n_155) );
OR2x6_ASAP7_75t_L g112 ( .A(n_35), .B(n_113), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_36), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_37), .B(n_134), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_39), .A2(n_193), .B1(n_226), .B2(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_40), .B(n_539), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g150 ( .A1(n_41), .A2(n_79), .B1(n_151), .B2(n_153), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_42), .B(n_144), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_43), .B(n_167), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_44), .B(n_129), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_45), .B(n_144), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_46), .Y(n_534) );
AND2x2_ASAP7_75t_L g233 ( .A(n_47), .B(n_171), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_48), .B(n_171), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_49), .Y(n_649) );
HB1xp67_ASAP7_75t_SL g720 ( .A(n_49), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_51), .B(n_144), .Y(n_482) );
INVx1_ASAP7_75t_L g137 ( .A(n_52), .Y(n_137) );
INVx1_ASAP7_75t_L g146 ( .A(n_52), .Y(n_146) );
AND2x2_ASAP7_75t_L g483 ( .A(n_53), .B(n_171), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_54), .A2(n_72), .B1(n_134), .B2(n_153), .C(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_55), .B(n_134), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_56), .B(n_143), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_57), .B(n_226), .Y(n_498) );
AOI21xp5_ASAP7_75t_SL g523 ( .A1(n_58), .A2(n_153), .B(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g174 ( .A(n_59), .B(n_171), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_60), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_61), .B(n_165), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_62), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_SL g215 ( .A(n_63), .B(n_172), .Y(n_215) );
INVx1_ASAP7_75t_L g463 ( .A(n_64), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_65), .A2(n_151), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g481 ( .A(n_66), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_67), .B(n_165), .Y(n_192) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_68), .B(n_129), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_69), .A2(n_153), .B(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g142 ( .A(n_70), .Y(n_142) );
INVx1_ASAP7_75t_L g148 ( .A(n_70), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_71), .B(n_134), .Y(n_516) );
AND2x2_ASAP7_75t_L g565 ( .A(n_73), .B(n_248), .Y(n_565) );
INVx1_ASAP7_75t_L g465 ( .A(n_74), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_75), .A2(n_153), .B(n_562), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_76), .A2(n_128), .B(n_153), .C(n_536), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g133 ( .A1(n_77), .A2(n_82), .B1(n_134), .B2(n_143), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_78), .B(n_143), .Y(n_169) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_81), .B(n_248), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_83), .A2(n_153), .B1(n_511), .B2(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_84), .B(n_167), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_85), .B(n_167), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g797 ( .A1(n_86), .A2(n_117), .B1(n_798), .B2(n_802), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_87), .A2(n_151), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g525 ( .A(n_89), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_90), .B(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g517 ( .A(n_91), .B(n_248), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_92), .A2(n_488), .B(n_489), .C(n_491), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_93), .B(n_143), .Y(n_232) );
INVxp67_ASAP7_75t_L g247 ( .A(n_94), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_95), .B(n_165), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_96), .A2(n_151), .B(n_212), .Y(n_211) );
BUFx2_ASAP7_75t_L g107 ( .A(n_97), .Y(n_107) );
BUFx2_ASAP7_75t_SL g828 ( .A(n_97), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_98), .B(n_144), .Y(n_526) );
BUFx4f_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_104), .B(n_107), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_SL g807 ( .A(n_105), .B(n_107), .Y(n_807) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_105), .A2(n_826), .B(n_829), .Y(n_825) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_R g821 ( .A(n_109), .Y(n_821) );
BUFx2_ASAP7_75t_L g830 ( .A(n_109), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
OR2x6_ASAP7_75t_SL g450 ( .A(n_110), .B(n_111), .Y(n_450) );
AND2x6_ASAP7_75t_SL g796 ( .A(n_110), .B(n_112), .Y(n_796) );
OR2x2_ASAP7_75t_L g805 ( .A(n_110), .B(n_112), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_118), .B(n_797), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_450), .B1(n_451), .B2(n_793), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g798 ( .A1(n_121), .A2(n_452), .B1(n_799), .B2(n_800), .Y(n_798) );
AND3x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_321), .C(n_395), .Y(n_121) );
NOR3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_263), .C(n_294), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_196), .B(n_205), .C(n_234), .Y(n_123) );
AOI21x1_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_175), .B(n_194), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_125), .A2(n_297), .B1(n_303), .B2(n_306), .Y(n_296) );
AND2x2_ASAP7_75t_L g430 ( .A(n_125), .B(n_198), .Y(n_430) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_159), .Y(n_125) );
BUFx2_ASAP7_75t_L g201 ( .A(n_126), .Y(n_201) );
AND2x2_ASAP7_75t_L g289 ( .A(n_126), .B(n_160), .Y(n_289) );
AND2x2_ASAP7_75t_L g360 ( .A(n_126), .B(n_204), .Y(n_360) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_127), .Y(n_254) );
AOI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B(n_158), .Y(n_127) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_128), .A2(n_509), .B(n_517), .Y(n_508) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_128), .A2(n_509), .B(n_517), .Y(n_580) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_129), .A2(n_210), .B(n_211), .Y(n_209) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_129), .A2(n_502), .B(n_506), .Y(n_501) );
BUFx4f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx3_ASAP7_75t_L g226 ( .A(n_130), .Y(n_226) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_131), .B(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g193 ( .A(n_131), .B(n_173), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_150), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_134), .A2(n_153), .B1(n_241), .B2(n_243), .Y(n_240) );
INVx1_ASAP7_75t_L g499 ( .A(n_134), .Y(n_499) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_140), .Y(n_134) );
INVx1_ASAP7_75t_L g532 ( .A(n_135), .Y(n_532) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_138), .Y(n_135) );
OR2x6_ASAP7_75t_L g464 ( .A(n_136), .B(n_157), .Y(n_464) );
INVxp33_ASAP7_75t_L g514 ( .A(n_136), .Y(n_514) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g152 ( .A(n_137), .B(n_139), .Y(n_152) );
AND2x4_ASAP7_75t_L g165 ( .A(n_137), .B(n_147), .Y(n_165) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g533 ( .A(n_140), .Y(n_533) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x6_ASAP7_75t_L g151 ( .A(n_141), .B(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
AND2x6_ASAP7_75t_L g167 ( .A(n_142), .B(n_145), .Y(n_167) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_149), .Y(n_143) );
INVx1_ASAP7_75t_L g251 ( .A(n_144), .Y(n_251) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_147), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx5_ASAP7_75t_L g168 ( .A(n_149), .Y(n_168) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_149), .Y(n_491) );
AND2x4_ASAP7_75t_L g153 ( .A(n_152), .B(n_154), .Y(n_153) );
INVxp67_ASAP7_75t_L g497 ( .A(n_153), .Y(n_497) );
NOR2x1p5_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
INVx1_ASAP7_75t_L g515 ( .A(n_156), .Y(n_515) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g253 ( .A(n_159), .B(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g195 ( .A(n_160), .B(n_185), .Y(n_195) );
OR2x2_ASAP7_75t_L g203 ( .A(n_160), .B(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g258 ( .A(n_160), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g305 ( .A(n_160), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_160), .B(n_204), .Y(n_313) );
AND2x2_ASAP7_75t_L g350 ( .A(n_160), .B(n_254), .Y(n_350) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_160), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_160), .B(n_184), .Y(n_391) );
AO21x2_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_170), .B(n_174), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_169), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_166), .B(n_168), .Y(n_163) );
INVxp67_ASAP7_75t_L g470 ( .A(n_165), .Y(n_470) );
INVxp67_ASAP7_75t_L g468 ( .A(n_167), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_168), .A2(n_180), .B(n_181), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_168), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_168), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_168), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_168), .A2(n_230), .B(n_231), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_168), .B(n_193), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_168), .A2(n_464), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g503 ( .A1(n_168), .A2(n_464), .B(n_504), .C(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g511 ( .A(n_168), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_168), .A2(n_464), .B(n_525), .C(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_168), .A2(n_537), .B(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g562 ( .A1(n_168), .A2(n_464), .B(n_563), .C(n_564), .Y(n_562) );
AO21x2_ASAP7_75t_L g176 ( .A1(n_170), .A2(n_177), .B(n_183), .Y(n_176) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_177), .B(n_183), .Y(n_204) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_170), .A2(n_559), .B(n_565), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
OA21x2_ASAP7_75t_L g218 ( .A1(n_171), .A2(n_219), .B(n_223), .Y(n_218) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g292 ( .A(n_175), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_175), .B(n_253), .Y(n_348) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_175), .Y(n_449) );
AND2x4_ASAP7_75t_L g175 ( .A(n_176), .B(n_184), .Y(n_175) );
AND2x2_ASAP7_75t_L g194 ( .A(n_176), .B(n_195), .Y(n_194) );
OR2x2_ASAP7_75t_L g274 ( .A(n_176), .B(n_185), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_176), .B(n_305), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_178), .B(n_182), .Y(n_177) );
AND2x2_ASAP7_75t_L g341 ( .A(n_184), .B(n_258), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_184), .B(n_253), .Y(n_397) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g199 ( .A(n_185), .Y(n_199) );
AND2x2_ASAP7_75t_L g268 ( .A(n_185), .B(n_259), .Y(n_268) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_185), .Y(n_288) );
AND2x4_ASAP7_75t_L g295 ( .A(n_185), .B(n_204), .Y(n_295) );
AND2x2_ASAP7_75t_SL g442 ( .A(n_185), .B(n_254), .Y(n_442) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_193), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_193), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_193), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_193), .B(n_247), .Y(n_246) );
NOR3xp33_ASAP7_75t_L g249 ( .A(n_193), .B(n_250), .C(n_251), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_193), .A2(n_523), .B(n_527), .Y(n_522) );
INVx1_ASAP7_75t_L g421 ( .A(n_194), .Y(n_421) );
INVx1_ASAP7_75t_L g363 ( .A(n_195), .Y(n_363) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_200), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
OR2x2_ASAP7_75t_L g285 ( .A(n_199), .B(n_203), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_199), .B(n_254), .Y(n_378) );
AND2x2_ASAP7_75t_L g380 ( .A(n_199), .B(n_202), .Y(n_380) );
AOI32xp33_ASAP7_75t_L g446 ( .A1(n_199), .A2(n_262), .A3(n_417), .B1(n_447), .B2(n_449), .Y(n_446) );
AND2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
AND2x2_ASAP7_75t_L g272 ( .A(n_201), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g390 ( .A(n_201), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g413 ( .A(n_201), .B(n_274), .Y(n_413) );
AND2x2_ASAP7_75t_L g440 ( .A(n_201), .B(n_341), .Y(n_440) );
AND2x2_ASAP7_75t_L g366 ( .A(n_202), .B(n_254), .Y(n_366) );
AND2x2_ASAP7_75t_L g441 ( .A(n_202), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
NOR2x1p5_ASAP7_75t_L g299 ( .A(n_207), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g317 ( .A(n_207), .Y(n_317) );
OR2x2_ASAP7_75t_L g345 ( .A(n_207), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x4_ASAP7_75t_SL g262 ( .A(n_208), .B(n_239), .Y(n_262) );
AND2x4_ASAP7_75t_L g278 ( .A(n_208), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g281 ( .A(n_208), .B(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g309 ( .A(n_208), .B(n_218), .Y(n_309) );
OR2x2_ASAP7_75t_L g334 ( .A(n_208), .B(n_283), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_208), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_208), .B(n_218), .Y(n_369) );
INVx2_ASAP7_75t_L g385 ( .A(n_208), .Y(n_385) );
AND2x2_ASAP7_75t_L g400 ( .A(n_208), .B(n_238), .Y(n_400) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_208), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_208), .Y(n_429) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_215), .Y(n_208) );
AND2x2_ASAP7_75t_L g293 ( .A(n_216), .B(n_278), .Y(n_293) );
AND2x2_ASAP7_75t_L g314 ( .A(n_216), .B(n_262), .Y(n_314) );
INVx1_ASAP7_75t_L g346 ( .A(n_216), .Y(n_346) );
AND2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_224), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g237 ( .A(n_218), .Y(n_237) );
INVx2_ASAP7_75t_L g283 ( .A(n_218), .Y(n_283) );
BUFx3_ASAP7_75t_L g300 ( .A(n_218), .Y(n_300) );
AND2x2_ASAP7_75t_L g339 ( .A(n_218), .B(n_224), .Y(n_339) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_218), .Y(n_437) );
INVx2_ASAP7_75t_L g252 ( .A(n_224), .Y(n_252) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_224), .Y(n_261) );
INVx1_ASAP7_75t_L g277 ( .A(n_224), .Y(n_277) );
OR2x2_ASAP7_75t_L g282 ( .A(n_224), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g302 ( .A(n_224), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_224), .B(n_279), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_224), .B(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_233), .Y(n_225) );
INVx4_ASAP7_75t_L g248 ( .A(n_226), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_226), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_232), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_235), .A2(n_253), .B(n_255), .Y(n_234) );
AND2x2_ASAP7_75t_SL g235 ( .A(n_236), .B(n_238), .Y(n_235) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_236), .Y(n_445) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVxp67_ASAP7_75t_SL g271 ( .A(n_237), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_237), .B(n_277), .Y(n_319) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_237), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_238), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g324 ( .A(n_238), .B(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g375 ( .A(n_238), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_238), .A2(n_380), .B1(n_381), .B2(n_386), .C(n_389), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_238), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_252), .Y(n_238) );
INVx3_ASAP7_75t_L g279 ( .A(n_239), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_239), .B(n_283), .Y(n_383) );
AND2x2_ASAP7_75t_L g412 ( .A(n_239), .B(n_385), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_239), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_245), .Y(n_239) );
INVx3_ASAP7_75t_L g476 ( .A(n_248), .Y(n_476) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_248), .A2(n_476), .B1(n_487), .B2(n_492), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_251), .A2(n_463), .B1(n_464), .B2(n_465), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_251), .B(n_490), .Y(n_489) );
AND2x2_ASAP7_75t_L g320 ( .A(n_253), .B(n_295), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_253), .A2(n_273), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g257 ( .A(n_254), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g266 ( .A(n_254), .Y(n_266) );
OR2x2_ASAP7_75t_L g312 ( .A(n_254), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_254), .B(n_295), .Y(n_404) );
OR2x2_ASAP7_75t_L g436 ( .A(n_254), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g448 ( .A(n_254), .B(n_354), .Y(n_448) );
INVxp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx2_ASAP7_75t_L g326 ( .A(n_257), .Y(n_326) );
INVx3_ASAP7_75t_SL g392 ( .A(n_258), .Y(n_392) );
INVxp67_ASAP7_75t_L g342 ( .A(n_260), .Y(n_342) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AOI322xp5_ASAP7_75t_L g264 ( .A1(n_262), .A2(n_265), .A3(n_269), .B1(n_272), .B2(n_275), .C1(n_280), .C2(n_284), .Y(n_264) );
INVx1_ASAP7_75t_SL g353 ( .A(n_262), .Y(n_353) );
AND2x4_ASAP7_75t_L g438 ( .A(n_262), .B(n_325), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_286), .Y(n_263) );
NOR2x1_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
OR2x2_ASAP7_75t_L g291 ( .A(n_266), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g387 ( .A(n_266), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g415 ( .A(n_266), .B(n_268), .Y(n_415) );
AOI32xp33_ASAP7_75t_L g416 ( .A1(n_266), .A2(n_267), .A3(n_417), .B1(n_419), .B2(n_422), .Y(n_416) );
OR2x2_ASAP7_75t_L g420 ( .A(n_266), .B(n_313), .Y(n_420) );
NAND3xp33_ASAP7_75t_L g376 ( .A(n_267), .B(n_292), .C(n_377), .Y(n_376) );
OAI22xp33_ASAP7_75t_SL g396 ( .A1(n_267), .A2(n_333), .B1(n_397), .B2(n_398), .Y(n_396) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g399 ( .A(n_270), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_274), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OAI322xp33_ASAP7_75t_L g322 ( .A1(n_278), .A2(n_282), .A3(n_291), .B1(n_323), .B2(n_326), .C1(n_327), .C2(n_328), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_278), .B(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_278), .B(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g301 ( .A(n_279), .B(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g333 ( .A(n_279), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_279), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g394 ( .A(n_282), .Y(n_394) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_283), .Y(n_325) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .B(n_293), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_289), .B(n_337), .Y(n_336) );
AOI322xp5_ASAP7_75t_SL g431 ( .A1(n_289), .A2(n_295), .A3(n_412), .B1(n_430), .B2(n_432), .C1(n_435), .C2(n_438), .Y(n_431) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_296), .B(n_310), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_295), .B(n_305), .Y(n_327) );
INVx2_ASAP7_75t_SL g337 ( .A(n_295), .Y(n_337) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_SL g362 ( .A(n_301), .Y(n_362) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_302), .Y(n_332) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g407 ( .A(n_308), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g361 ( .A(n_309), .B(n_362), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_314), .B1(n_315), .B2(n_320), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR4xp75_ASAP7_75t_L g321 ( .A(n_322), .B(n_335), .C(n_355), .D(n_371), .Y(n_321) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_330), .B(n_333), .Y(n_329) );
INVxp67_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_333), .A2(n_410), .B1(n_413), .B2(n_414), .Y(n_409) );
OR2x2_ASAP7_75t_L g374 ( .A(n_334), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g418 ( .A(n_334), .Y(n_418) );
OAI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B1(n_340), .B2(n_342), .C(n_343), .Y(n_335) );
INVx2_ASAP7_75t_L g354 ( .A(n_339), .Y(n_354) );
AND2x2_ASAP7_75t_L g411 ( .A(n_339), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B1(n_349), .B2(n_351), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g406 ( .A(n_350), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_351), .A2(n_357), .B1(n_373), .B2(n_376), .Y(n_372) );
INVx1_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
OAI221xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_361), .B1(n_363), .B2(n_364), .C(n_832), .Y(n_355) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
OR2x2_ASAP7_75t_L g423 ( .A(n_362), .B(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_379), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_392), .B(n_393), .Y(n_389) );
NOR3xp33_ASAP7_75t_SL g395 ( .A(n_396), .B(n_401), .C(n_425), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_402), .B(n_416), .Y(n_401) );
O2A1O1Ixp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B(n_407), .C(n_409), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g417 ( .A(n_408), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx1_ASAP7_75t_SL g422 ( .A(n_423), .Y(n_422) );
NAND4xp25_ASAP7_75t_SL g425 ( .A(n_426), .B(n_431), .C(n_439), .D(n_446), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_441), .B(n_443), .Y(n_439) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
CKINVDCx11_ASAP7_75t_R g801 ( .A(n_450), .Y(n_801) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI211x1_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_649), .B(n_650), .C(n_790), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND4x1_ASAP7_75t_L g790 ( .A(n_454), .B(n_651), .C(n_791), .D(n_792), .Y(n_790) );
NAND3x1_ASAP7_75t_L g813 ( .A(n_454), .B(n_651), .C(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_617), .Y(n_454) );
AOI211xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_540), .B(n_552), .C(n_593), .Y(n_455) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_472), .B(n_518), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_SL g540 ( .A1(n_458), .A2(n_541), .B(n_546), .C(n_551), .Y(n_540) );
NAND2x1_ASAP7_75t_L g670 ( .A(n_458), .B(n_671), .Y(n_670) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_458), .B(n_690), .Y(n_761) );
AND2x2_ASAP7_75t_L g780 ( .A(n_458), .B(n_520), .Y(n_780) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx3_ASAP7_75t_L g557 ( .A(n_459), .Y(n_557) );
AND2x2_ASAP7_75t_L g628 ( .A(n_459), .B(n_558), .Y(n_628) );
AND2x2_ASAP7_75t_L g633 ( .A(n_459), .B(n_529), .Y(n_633) );
NOR2x1_ASAP7_75t_SL g749 ( .A(n_459), .B(n_520), .Y(n_749) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_466), .B(n_471), .Y(n_461) );
INVxp67_ASAP7_75t_L g488 ( .A(n_464), .Y(n_488) );
INVx2_ASAP7_75t_L g539 ( .A(n_464), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_469), .B2(n_470), .Y(n_466) );
INVx1_ASAP7_75t_SL g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_500), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g664 ( .A(n_474), .B(n_598), .Y(n_664) );
AND2x2_ASAP7_75t_L g781 ( .A(n_474), .B(n_622), .Y(n_781) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_475), .B(n_550), .Y(n_549) );
INVx2_ASAP7_75t_L g570 ( .A(n_475), .Y(n_570) );
AND2x2_ASAP7_75t_L g578 ( .A(n_475), .B(n_579), .Y(n_578) );
NOR2xp67_ASAP7_75t_L g716 ( .A(n_475), .B(n_484), .Y(n_716) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_483), .Y(n_475) );
AO21x2_ASAP7_75t_L g601 ( .A1(n_476), .A2(n_477), .B(n_483), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
AND2x2_ASAP7_75t_L g668 ( .A(n_484), .B(n_508), .Y(n_668) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g544 ( .A(n_485), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g548 ( .A(n_485), .Y(n_548) );
INVx1_ASAP7_75t_L g568 ( .A(n_485), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_485), .B(n_601), .Y(n_625) );
AND2x2_ASAP7_75t_L g674 ( .A(n_485), .B(n_501), .Y(n_674) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_497), .B1(n_498), .B2(n_499), .Y(n_493) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g629 ( .A(n_500), .B(n_624), .Y(n_629) );
AND2x2_ASAP7_75t_L g685 ( .A(n_500), .B(n_568), .Y(n_685) );
AND2x2_ASAP7_75t_L g700 ( .A(n_500), .B(n_614), .Y(n_700) );
AND2x2_ASAP7_75t_L g737 ( .A(n_500), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g753 ( .A(n_500), .Y(n_753) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
INVx2_ASAP7_75t_L g545 ( .A(n_501), .Y(n_545) );
INVx1_ASAP7_75t_L g550 ( .A(n_501), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_501), .B(n_580), .Y(n_583) );
INVx1_ASAP7_75t_L g597 ( .A(n_501), .Y(n_597) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_501), .Y(n_607) );
INVxp67_ASAP7_75t_L g623 ( .A(n_501), .Y(n_623) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g542 ( .A(n_508), .Y(n_542) );
AND2x4_ASAP7_75t_L g569 ( .A(n_508), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_510), .B(n_516), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g551 ( .A(n_518), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_518), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_SL g572 ( .A(n_519), .B(n_573), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_519), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_519), .B(n_586), .Y(n_729) );
HB1xp67_ASAP7_75t_L g767 ( .A(n_519), .Y(n_767) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_528), .Y(n_519) );
INVx2_ASAP7_75t_L g592 ( .A(n_520), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_520), .B(n_529), .Y(n_603) );
INVx4_ASAP7_75t_L g611 ( .A(n_520), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_520), .B(n_587), .Y(n_647) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_520), .Y(n_660) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AND2x4_ASAP7_75t_L g638 ( .A(n_528), .B(n_611), .Y(n_638) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x4_ASAP7_75t_L g589 ( .A(n_529), .B(n_557), .Y(n_589) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_529), .Y(n_610) );
INVx2_ASAP7_75t_L g659 ( .A(n_529), .Y(n_659) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
NOR3xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .C(n_534), .Y(n_531) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_542), .B(n_547), .Y(n_648) );
NAND2x1_ASAP7_75t_SL g762 ( .A(n_542), .B(n_544), .Y(n_762) );
OR2x2_ASAP7_75t_L g641 ( .A(n_543), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g744 ( .A(n_543), .Y(n_744) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g634 ( .A(n_544), .B(n_569), .Y(n_634) );
AND2x2_ASAP7_75t_L g750 ( .A(n_544), .B(n_743), .Y(n_750) );
OAI221xp5_ASAP7_75t_L g758 ( .A1(n_546), .A2(n_759), .B1(n_762), .B2(n_763), .C(n_765), .Y(n_758) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_547), .A2(n_703), .B1(n_705), .B2(n_707), .Y(n_702) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_548), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g616 ( .A(n_548), .Y(n_616) );
BUFx2_ASAP7_75t_L g697 ( .A(n_548), .Y(n_697) );
AND2x2_ASAP7_75t_L g667 ( .A(n_549), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_553), .B(n_571), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_566), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g640 ( .A(n_556), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_556), .B(n_766), .C(n_767), .D(n_768), .Y(n_765) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
INVx1_ASAP7_75t_L g575 ( .A(n_557), .Y(n_575) );
AND2x2_ASAP7_75t_L g658 ( .A(n_557), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g574 ( .A(n_558), .Y(n_574) );
INVx2_ASAP7_75t_L g588 ( .A(n_558), .Y(n_588) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_558), .Y(n_615) );
INVx1_ASAP7_75t_L g632 ( .A(n_558), .Y(n_632) );
HB1xp67_ASAP7_75t_L g672 ( .A(n_558), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_561), .Y(n_559) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx1_ASAP7_75t_L g779 ( .A(n_567), .Y(n_779) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g577 ( .A(n_568), .Y(n_577) );
AND2x2_ASAP7_75t_L g673 ( .A(n_569), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g773 ( .A(n_569), .B(n_774), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B1(n_581), .B2(n_584), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_573), .B(n_638), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_573), .B(n_737), .Y(n_736) );
AND2x4_ASAP7_75t_L g754 ( .A(n_573), .B(n_732), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_573), .A2(n_609), .B(n_731), .Y(n_784) );
AND2x4_ASAP7_75t_SL g573 ( .A(n_574), .B(n_575), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_574), .B(n_658), .Y(n_695) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_574), .Y(n_711) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
AND2x2_ASAP7_75t_L g581 ( .A(n_577), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g598 ( .A(n_579), .Y(n_598) );
AND2x2_ASAP7_75t_L g622 ( .A(n_579), .B(n_623), .Y(n_622) );
AND2x4_ASAP7_75t_L g743 ( .A(n_579), .B(n_600), .Y(n_743) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_580), .B(n_601), .Y(n_642) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g718 ( .A(n_583), .B(n_625), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_590), .Y(n_584) );
INVx1_ASAP7_75t_L g699 ( .A(n_585), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g594 ( .A(n_586), .B(n_595), .C(n_599), .Y(n_594) );
AND2x2_ASAP7_75t_L g637 ( .A(n_586), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g666 ( .A(n_586), .B(n_609), .Y(n_666) );
AND2x2_ASAP7_75t_L g748 ( .A(n_586), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g774 ( .A(n_586), .Y(n_774) );
INVx1_ASAP7_75t_L g788 ( .A(n_586), .Y(n_788) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g591 ( .A(n_589), .B(n_592), .Y(n_591) );
INVx4_ASAP7_75t_L g747 ( .A(n_589), .Y(n_747) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g787 ( .A(n_591), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g690 ( .A(n_592), .Y(n_690) );
AO22x1_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_602), .B1(n_604), .B2(n_612), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_596), .B(n_600), .Y(n_680) );
INVx3_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
BUFx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx3_ASAP7_75t_L g614 ( .A(n_600), .Y(n_614) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g692 ( .A(n_601), .B(n_607), .Y(n_692) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_601), .Y(n_739) );
AOI31xp33_ASAP7_75t_L g643 ( .A1(n_602), .A2(n_644), .A3(n_646), .B(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_603), .A2(n_620), .B1(n_626), .B2(n_629), .Y(n_619) );
AND2x2_ASAP7_75t_L g703 ( .A(n_603), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g710 ( .A(n_603), .B(n_711), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_609), .B(n_764), .Y(n_763) );
AND2x4_ASAP7_75t_SL g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g639 ( .A(n_611), .B(n_640), .Y(n_639) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_611), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_616), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
AND2x2_ASAP7_75t_L g734 ( .A(n_614), .B(n_674), .Y(n_734) );
INVx1_ASAP7_75t_L g769 ( .A(n_614), .Y(n_769) );
AND2x2_ASAP7_75t_L g719 ( .A(n_615), .B(n_658), .Y(n_719) );
BUFx2_ASAP7_75t_L g764 ( .A(n_615), .Y(n_764) );
AND2x2_ASAP7_75t_L g707 ( .A(n_616), .B(n_708), .Y(n_707) );
NOR3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_635), .C(n_643), .Y(n_617) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_619), .B(n_630), .Y(n_618) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2x1p5_ASAP7_75t_L g621 ( .A(n_622), .B(n_624), .Y(n_621) );
AND2x2_ASAP7_75t_L g696 ( .A(n_622), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_SL g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_628), .B(n_638), .Y(n_661) );
AND2x2_ASAP7_75t_L g683 ( .A(n_628), .B(n_660), .Y(n_683) );
AND2x2_ASAP7_75t_SL g731 ( .A(n_628), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .Y(n_630) );
AND2x2_ASAP7_75t_L g786 ( .A(n_631), .B(n_660), .Y(n_786) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x2_ASAP7_75t_L g760 ( .A(n_632), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g677 ( .A(n_633), .Y(n_677) );
AND2x2_ASAP7_75t_L g777 ( .A(n_633), .B(n_660), .Y(n_777) );
AOI21xp33_ASAP7_75t_R g635 ( .A1(n_636), .A2(n_639), .B(n_641), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_637), .B(n_741), .Y(n_740) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_638), .Y(n_645) );
INVx1_ASAP7_75t_L g708 ( .A(n_642), .Y(n_708) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_644), .A2(n_662), .B1(n_676), .B2(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g676 ( .A(n_647), .B(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_649), .B(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_649), .B(n_756), .Y(n_755) );
NOR2xp67_ASAP7_75t_SL g791 ( .A(n_649), .B(n_722), .Y(n_791) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_720), .B(n_721), .C(n_755), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_686), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_675), .C(n_681), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_662), .B(n_665), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_661), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_657), .A2(n_696), .B1(n_699), .B2(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_L g733 ( .A(n_659), .Y(n_733) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g725 ( .A(n_664), .B(n_714), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_669), .B2(n_673), .Y(n_665) );
INVx1_ASAP7_75t_L g679 ( .A(n_668), .Y(n_679) );
AND2x4_ASAP7_75t_L g691 ( .A(n_668), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g727 ( .A(n_670), .Y(n_727) );
INVx1_ASAP7_75t_L g704 ( .A(n_671), .Y(n_704) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_673), .A2(n_683), .B1(n_731), .B2(n_734), .Y(n_730) );
INVxp67_ASAP7_75t_L g775 ( .A(n_674), .Y(n_775) );
NOR2x1_ASAP7_75t_L g689 ( .A(n_677), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
INVxp33_ASAP7_75t_L g789 ( .A(n_680), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g686 ( .A(n_687), .B(n_701), .Y(n_686) );
NAND2xp5_ASAP7_75t_SL g687 ( .A(n_688), .B(n_698), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B1(n_693), .B2(n_696), .Y(n_688) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
BUFx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_702), .B(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B1(n_717), .B2(n_719), .Y(n_709) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g766 ( .A(n_714), .Y(n_766) );
INVxp67_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g814 ( .A(n_723), .B(n_757), .Y(n_814) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_735), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_726), .B(n_730), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NAND4xp25_ASAP7_75t_SL g735 ( .A(n_736), .B(n_740), .C(n_745), .D(n_751), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g778 ( .A(n_743), .B(n_779), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_748), .B(n_750), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g792 ( .A(n_756), .Y(n_792) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR3x1_ASAP7_75t_L g757 ( .A(n_758), .B(n_770), .C(n_782), .Y(n_757) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_775), .B(n_776), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_773), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_780), .B2(n_781), .Y(n_776) );
INVx1_ASAP7_75t_L g783 ( .A(n_781), .Y(n_783) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B(n_785), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B(n_789), .Y(n_785) );
CKINVDCx11_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
CKINVDCx6p67_ASAP7_75t_R g799 ( .A(n_794), .Y(n_799) );
INVx3_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_SL g803 ( .A(n_804), .Y(n_803) );
INVx3_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVxp67_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_819), .B(n_822), .Y(n_809) );
OAI22xp5_ASAP7_75t_SL g810 ( .A1(n_811), .A2(n_815), .B1(n_817), .B2(n_818), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVxp67_ASAP7_75t_SL g817 ( .A(n_813), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_815), .Y(n_818) );
INVx1_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_SL g820 ( .A(n_821), .Y(n_820) );
NOR2xp33_ASAP7_75t_SL g822 ( .A(n_821), .B(n_823), .Y(n_822) );
INVx1_ASAP7_75t_SL g824 ( .A(n_825), .Y(n_824) );
CKINVDCx11_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
CKINVDCx8_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
endmodule