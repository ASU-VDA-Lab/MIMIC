module fake_jpeg_10968_n_472 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_23),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_53),
.B(n_69),
.Y(n_119)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx6p67_ASAP7_75t_R g107 ( 
.A(n_54),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_21),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_92),
.Y(n_112)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_15),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_68),
.B(n_77),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_43),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_73),
.B(n_90),
.Y(n_99)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_84),
.B(n_91),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_31),
.B(n_13),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_89),
.B(n_12),
.Y(n_105)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_41),
.B(n_13),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_95),
.Y(n_118)
);

NAND2xp33_ASAP7_75t_SL g94 ( 
.A(n_18),
.B(n_0),
.Y(n_94)
);

NOR2x1_ASAP7_75t_R g116 ( 
.A(n_94),
.B(n_73),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g96 ( 
.A(n_28),
.Y(n_96)
);

HAxp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_28),
.CON(n_110),
.SN(n_110)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_31),
.B1(n_28),
.B2(n_42),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_103),
.A2(n_126),
.B1(n_133),
.B2(n_138),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_105),
.B(n_27),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_110),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_24),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_66),
.A2(n_45),
.B1(n_42),
.B2(n_36),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_128),
.B1(n_132),
.B2(n_140),
.Y(n_166)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_39),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_125),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_67),
.A2(n_39),
.B1(n_18),
.B2(n_30),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_32),
.B1(n_45),
.B2(n_34),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_58),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_78),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_62),
.B(n_30),
.C(n_40),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_72),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_L g138 ( 
.A1(n_79),
.A2(n_46),
.B1(n_40),
.B2(n_37),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_85),
.A2(n_46),
.B1(n_37),
.B2(n_35),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_52),
.A2(n_35),
.B1(n_29),
.B2(n_27),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_149),
.B1(n_24),
.B2(n_54),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_57),
.A2(n_29),
.B1(n_11),
.B2(n_24),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_71),
.Y(n_150)
);

NAND2x1_ASAP7_75t_L g226 ( 
.A(n_150),
.B(n_152),
.Y(n_226)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_64),
.B1(n_60),
.B2(n_95),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_153),
.A2(n_175),
.B1(n_184),
.B2(n_186),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_97),
.B(n_51),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_154),
.B(n_180),
.C(n_63),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_155),
.B(n_190),
.Y(n_224)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_158),
.Y(n_227)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_159),
.Y(n_232)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_11),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_163),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_11),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_98),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_164),
.B(n_173),
.Y(n_229)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_117),
.Y(n_171)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_171),
.Y(n_219)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_172),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_174),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_81),
.B1(n_80),
.B2(n_91),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_0),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_176),
.B(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_100),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_1),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_185),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_102),
.B(n_61),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_120),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_181),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_110),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_140),
.A2(n_87),
.B1(n_86),
.B2(n_27),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_125),
.B(n_1),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_193),
.Y(n_238)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_141),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_189),
.Y(n_240)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_113),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_191),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_192),
.A2(n_199),
.B1(n_2),
.B2(n_4),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_132),
.A2(n_87),
.B1(n_86),
.B2(n_82),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_148),
.B1(n_101),
.B2(n_115),
.Y(n_212)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_195),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_107),
.B(n_61),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_106),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

INVx11_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_1),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_2),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_99),
.B(n_107),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_205),
.B(n_209),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_150),
.B(n_111),
.C(n_104),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_206),
.B(n_222),
.C(n_233),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_156),
.A2(n_139),
.B1(n_115),
.B2(n_145),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_208),
.A2(n_189),
.B1(n_174),
.B2(n_183),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_212),
.A2(n_215),
.B1(n_228),
.B2(n_192),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_179),
.A2(n_145),
.B1(n_129),
.B2(n_127),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_150),
.B(n_142),
.C(n_129),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_179),
.A2(n_131),
.B1(n_139),
.B2(n_142),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_63),
.C(n_124),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_199),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_237),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_156),
.A2(n_131),
.B(n_4),
.C(n_5),
.Y(n_236)
);

O2A1O1Ixp33_ASAP7_75t_L g262 ( 
.A1(n_236),
.A2(n_180),
.B(n_187),
.C(n_191),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_154),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_4),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_213),
.Y(n_246)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_184),
.B(n_193),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_248),
.A2(n_263),
.B(n_270),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_153),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_166),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_252),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_253),
.B(n_255),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_254),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_220),
.Y(n_257)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_257),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_165),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_259),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_222),
.B(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_227),
.Y(n_260)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_260),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_154),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_264),
.C(n_279),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_262),
.B(n_285),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_234),
.A2(n_180),
.B(n_181),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_170),
.C(n_167),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_195),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_265),
.B(n_277),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g266 ( 
.A(n_233),
.B(n_172),
.CI(n_160),
.CON(n_266),
.SN(n_266)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_266),
.B(n_281),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_267),
.B(n_272),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_159),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_269),
.B(n_271),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_224),
.A2(n_190),
.B(n_157),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_158),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_245),
.A2(n_151),
.B1(n_8),
.B2(n_9),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx11_ASAP7_75t_L g274 ( 
.A(n_221),
.Y(n_274)
);

BUFx24_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_215),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_275),
.A2(n_204),
.B1(n_217),
.B2(n_221),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_5),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_238),
.B(n_8),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_280),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_223),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_232),
.Y(n_282)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_228),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_283),
.B(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_205),
.A2(n_206),
.B(n_245),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_211),
.B(n_219),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_299),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_210),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_331)
);

MAJx2_ASAP7_75t_L g293 ( 
.A(n_251),
.B(n_212),
.C(n_204),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_201),
.C(n_214),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_286),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_302),
.A2(n_273),
.B1(n_254),
.B2(n_262),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_247),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_308),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_269),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_258),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_317),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_318),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_257),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_283),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_251),
.B(n_202),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_319),
.B(n_276),
.C(n_270),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_289),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_329),
.C(n_343),
.Y(n_358)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_325),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_318),
.A2(n_250),
.B1(n_268),
.B2(n_249),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_326),
.A2(n_340),
.B1(n_315),
.B2(n_295),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_327),
.A2(n_352),
.B1(n_301),
.B2(n_295),
.Y(n_357)
);

OAI32xp33_ASAP7_75t_L g328 ( 
.A1(n_298),
.A2(n_271),
.A3(n_285),
.B1(n_246),
.B2(n_266),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_328),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_276),
.Y(n_329)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_314),
.Y(n_334)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_334),
.Y(n_371)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_314),
.Y(n_335)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_264),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_338),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_307),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_266),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_339),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_301),
.A2(n_275),
.B1(n_248),
.B2(n_256),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_261),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_341),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g342 ( 
.A(n_310),
.B(n_276),
.CI(n_279),
.CON(n_342),
.SN(n_342)
);

MAJIxp5_ASAP7_75t_SL g356 ( 
.A(n_342),
.B(n_287),
.C(n_293),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_287),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_351),
.C(n_322),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_312),
.A2(n_256),
.B(n_236),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_345),
.A2(n_346),
.B(n_292),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_290),
.A2(n_281),
.B(n_221),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_292),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_347),
.B(n_353),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_290),
.A2(n_291),
.B(n_305),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_348),
.A2(n_291),
.B(n_296),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_284),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_350),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_282),
.C(n_280),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_315),
.A2(n_278),
.B1(n_260),
.B2(n_252),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_292),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_356),
.B(n_341),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_374),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_313),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_373),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_361),
.B(n_370),
.Y(n_396)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_324),
.Y(n_362)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_363),
.A2(n_352),
.B1(n_326),
.B2(n_328),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_300),
.C(n_306),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_379),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_339),
.A2(n_296),
.B1(n_303),
.B2(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_367),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_327),
.A2(n_303),
.B1(n_320),
.B2(n_322),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_380),
.C(n_351),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_333),
.A2(n_292),
.B(n_320),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_331),
.B(n_302),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_349),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_331),
.B(n_344),
.C(n_336),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_377),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_378),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_392),
.C(n_395),
.Y(n_413)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_355),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_386),
.B(n_388),
.Y(n_419)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_366),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_362),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_389),
.A2(n_399),
.B1(n_402),
.B2(n_387),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_376),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_390),
.B(n_398),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_363),
.A2(n_333),
.B1(n_348),
.B2(n_350),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_391),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_329),
.C(n_323),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_393),
.B(n_359),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_394),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_371),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_358),
.B(n_346),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_358),
.Y(n_408)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_396),
.A2(n_374),
.B(n_360),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_404),
.B(n_408),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_401),
.A2(n_360),
.B(n_361),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_406),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_401),
.A2(n_370),
.B(n_367),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_401),
.A2(n_397),
.B(n_384),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_409),
.B(n_410),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_369),
.B(n_356),
.C(n_380),
.D(n_375),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_384),
.A2(n_345),
.B(n_373),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_411),
.A2(n_412),
.B1(n_402),
.B2(n_399),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_381),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_395),
.C(n_383),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_R g433 ( 
.A(n_416),
.B(n_342),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_421),
.B(n_423),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_422),
.B(n_428),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_392),
.C(n_400),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_408),
.B(n_354),
.C(n_391),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_424),
.B(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_407),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_414),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_429),
.B(n_430),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_365),
.C(n_357),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_420),
.B(n_387),
.C(n_372),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_418),
.C(n_417),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_433),
.B(n_411),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_420),
.A2(n_371),
.B1(n_342),
.B2(n_332),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_434),
.A2(n_325),
.B1(n_297),
.B2(n_204),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_445),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_431),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_439),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_424),
.A2(n_409),
.B(n_410),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_441),
.B(n_442),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_446),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_428),
.A2(n_418),
.B(n_415),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_419),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_443),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_421),
.B(n_337),
.C(n_335),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_438),
.B(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_449),
.B(n_435),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_436),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_452),
.C(n_453),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_444),
.A2(n_423),
.B(n_432),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_451),
.A2(n_455),
.B(n_223),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_427),
.C(n_430),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_434),
.C(n_297),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_448),
.A2(n_443),
.B(n_446),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_457),
.B(n_459),
.Y(n_465)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_458),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_452),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_460),
.B(n_450),
.Y(n_466)
);

OA21x2_ASAP7_75t_SL g461 ( 
.A1(n_454),
.A2(n_216),
.B(n_218),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_461),
.A2(n_453),
.B(n_216),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_463),
.B(n_466),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_462),
.C(n_456),
.Y(n_467)
);

AOI321xp33_ASAP7_75t_L g469 ( 
.A1(n_467),
.A2(n_464),
.A3(n_447),
.B1(n_240),
.B2(n_242),
.C(n_218),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_468),
.C(n_447),
.Y(n_470)
);

A2O1A1Ixp33_ASAP7_75t_R g471 ( 
.A1(n_470),
.A2(n_242),
.B(n_225),
.C(n_243),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_225),
.Y(n_472)
);


endmodule