module fake_jpeg_4441_n_229 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_36),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_31),
.B(n_0),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_43),
.Y(n_69)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_22),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_49),
.Y(n_65)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_7),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_19),
.B1(n_17),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_25),
.B1(n_21),
.B2(n_28),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_56),
.A2(n_50),
.B1(n_73),
.B2(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_58),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_37),
.B1(n_31),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_77),
.B1(n_47),
.B2(n_16),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_31),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_68),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_63),
.B(n_75),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_38),
.C(n_31),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_47),
.Y(n_97)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_31),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_19),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_72),
.B1(n_78),
.B2(n_16),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_36),
.B1(n_33),
.B2(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_36),
.B1(n_33),
.B2(n_17),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_15),
.B1(n_27),
.B2(n_22),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_43),
.A2(n_32),
.B1(n_33),
.B2(n_30),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_42),
.B(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_22),
.Y(n_94)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_54),
.B1(n_77),
.B2(n_71),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_56),
.B1(n_70),
.B2(n_80),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_53),
.B(n_49),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_95),
.Y(n_118)
);

NOR2x1p5_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_32),
.Y(n_91)
);

XOR2x1_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_72),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_62),
.A2(n_28),
.B(n_25),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_97),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_55),
.Y(n_117)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_21),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_98),
.B(n_104),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_59),
.B1(n_65),
.B2(n_61),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_73),
.B1(n_65),
.B2(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_64),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_59),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_108),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_111),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_119),
.B1(n_123),
.B2(n_125),
.Y(n_136)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

OA21x2_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_79),
.B(n_68),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_88),
.CON(n_142),
.SN(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_91),
.B1(n_89),
.B2(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_126),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_69),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_88),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_130),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_89),
.B1(n_96),
.B2(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_141),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_143),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_100),
.B1(n_102),
.B2(n_93),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_137),
.A2(n_139),
.B1(n_151),
.B2(n_116),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_144),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_93),
.B1(n_85),
.B2(n_81),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_20),
.B(n_81),
.Y(n_141)
);

XOR2x2_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_126),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_130),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_153),
.C(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_108),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_83),
.B1(n_95),
.B2(n_67),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_67),
.C(n_21),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_20),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_115),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_131),
.B1(n_150),
.B2(n_137),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_168),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_124),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_164),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_122),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_112),
.B(n_129),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_170),
.B(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_106),
.C(n_113),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_145),
.B1(n_139),
.B2(n_132),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_30),
.Y(n_173)
);

AO221x1_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_156),
.B1(n_26),
.B2(n_30),
.C(n_157),
.Y(n_182)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_133),
.B(n_141),
.C(n_136),
.D(n_152),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_179),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_151),
.B1(n_133),
.B2(n_144),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_176),
.Y(n_195)
);

OAI321xp33_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_147),
.A3(n_149),
.B1(n_154),
.B2(n_153),
.C(n_30),
.Y(n_180)
);

AOI31xp67_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_26),
.A3(n_24),
.B(n_167),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_186),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_147),
.B1(n_149),
.B2(n_20),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_183),
.B(n_164),
.C(n_159),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_179),
.C(n_24),
.Y(n_204)
);

AOI21x1_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_167),
.B(n_171),
.Y(n_189)
);

NOR2xp67_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_24),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_187),
.A2(n_184),
.B(n_181),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_190),
.A2(n_192),
.B(n_193),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_176),
.A2(n_161),
.B(n_169),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_196),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_158),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_8),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_178),
.A2(n_168),
.B1(n_1),
.B2(n_2),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_0),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_185),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_208),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_181),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_177),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_24),
.C(n_0),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_207),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_206),
.C(n_196),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_24),
.C(n_26),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_213),
.C(n_8),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_195),
.A3(n_199),
.B1(n_2),
.B2(n_3),
.C1(n_5),
.C2(n_6),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_214),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_215),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_1),
.B(n_5),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_207),
.C(n_3),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_9),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_220),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_224),
.A3(n_225),
.B1(n_14),
.B2(n_10),
.C1(n_11),
.C2(n_13),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_215),
.B1(n_212),
.B2(n_11),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_9),
.A3(n_10),
.B1(n_13),
.B2(n_14),
.C1(n_215),
.C2(n_210),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_10),
.Y(n_229)
);


endmodule