module fake_aes_7282_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_5), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
BUFx3_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_10), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_15), .A2(n_9), .B(n_1), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_16), .B(n_0), .Y(n_19) );
A2O1A1Ixp33_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_1), .B(n_2), .C(n_3), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_14), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g22 ( .A1(n_15), .A2(n_5), .B(n_6), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_21), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
AND2x4_ASAP7_75t_L g26 ( .A(n_25), .B(n_20), .Y(n_26) );
BUFx2_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_11), .Y(n_28) );
OAI21xp33_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_24), .B(n_23), .Y(n_29) );
OAI222xp33_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_11), .B1(n_12), .B2(n_13), .C1(n_14), .C2(n_15), .Y(n_30) );
NAND2xp5_ASAP7_75t_SL g31 ( .A(n_29), .B(n_28), .Y(n_31) );
AOI221xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_28), .B1(n_26), .B2(n_27), .C(n_24), .Y(n_32) );
AOI32xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_28), .A3(n_12), .B1(n_26), .B2(n_16), .Y(n_33) );
CKINVDCx16_ASAP7_75t_R g34 ( .A(n_31), .Y(n_34) );
AO22x2_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_26), .B1(n_29), .B2(n_18), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_27), .B1(n_17), .B2(n_33), .Y(n_36) );
endmodule