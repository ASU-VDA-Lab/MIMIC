module fake_jpeg_13412_n_197 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_197);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_197;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_12),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_0),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_1),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_25),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_0),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_70),
.B1(n_63),
.B2(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_94),
.B1(n_95),
.B2(n_68),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_85),
.A2(n_70),
.B1(n_65),
.B2(n_81),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_88),
.A2(n_59),
.B1(n_56),
.B2(n_71),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_57),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_63),
.B1(n_75),
.B2(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_102),
.B1(n_74),
.B2(n_80),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_89),
.A2(n_75),
.B1(n_71),
.B2(n_56),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_108),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_73),
.B(n_62),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_114),
.B(n_7),
.Y(n_138)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_60),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_92),
.A2(n_64),
.B1(n_69),
.B2(n_73),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_112),
.A2(n_118),
.B1(n_79),
.B2(n_72),
.Y(n_123)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_66),
.B1(n_68),
.B2(n_5),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_29),
.Y(n_136)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_101),
.B(n_84),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_4),
.B(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_78),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_8),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_123),
.A2(n_125),
.B1(n_133),
.B2(n_115),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_124),
.A2(n_15),
.B1(n_16),
.B2(n_21),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_136),
.B(n_37),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

AO22x2_ASAP7_75t_L g131 ( 
.A1(n_121),
.A2(n_31),
.B1(n_53),
.B2(n_52),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_119),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_142),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_14),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_117),
.B(n_10),
.Y(n_140)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_113),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_107),
.B(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_39),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_147),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_13),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_152),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_34),
.B1(n_50),
.B2(n_20),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_127),
.A2(n_16),
.B1(n_23),
.B2(n_24),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_41),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_160),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_142),
.B1(n_131),
.B2(n_128),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_146),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_171),
.B(n_153),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_128),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_155),
.C(n_129),
.Y(n_182)
);

AO22x2_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_161),
.B1(n_155),
.B2(n_149),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_180),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_162),
.A2(n_144),
.B(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_177),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_163),
.A2(n_171),
.B1(n_137),
.B2(n_141),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_175),
.A2(n_169),
.B1(n_174),
.B2(n_165),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_185),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_183),
.A2(n_178),
.B(n_180),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_184),
.B(n_167),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_189),
.A2(n_187),
.B1(n_170),
.B2(n_172),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_186),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_168),
.B(n_159),
.C(n_54),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_193),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_195),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_196),
.B(n_48),
.Y(n_197)
);


endmodule