module real_jpeg_15964_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_620;
wire n_332;
wire n_366;
wire n_456;
wire n_578;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_411;
wire n_382;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_412;
wire n_405;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_531;
wire n_285;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_1),
.Y(n_108)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_1),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_1),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_1),
.Y(n_340)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_2),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_3),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_3),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_3),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_3),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_4),
.A2(n_124),
.B1(n_128),
.B2(n_133),
.Y(n_123)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_4),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_4),
.A2(n_133),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_4),
.A2(n_133),
.B1(n_372),
.B2(n_374),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_SL g583 ( 
.A1(n_4),
.A2(n_133),
.B1(n_247),
.B2(n_584),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_5),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_5),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_5),
.A2(n_232),
.B1(n_252),
.B2(n_257),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_5),
.A2(n_232),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_5),
.A2(n_151),
.B1(n_232),
.B2(n_245),
.Y(n_393)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_6),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_6),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_7),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_7),
.A2(n_74),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_7),
.A2(n_74),
.B1(n_347),
.B2(n_349),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_7),
.A2(n_74),
.B1(n_441),
.B2(n_444),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_114),
.B1(n_117),
.B2(n_118),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_8),
.A2(n_117),
.B1(n_216),
.B2(n_220),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_8),
.A2(n_117),
.B1(n_353),
.B2(n_356),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_8),
.A2(n_117),
.B1(n_569),
.B2(n_570),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_9),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_9),
.A2(n_173),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_9),
.A2(n_173),
.B1(n_573),
.B2(n_577),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_SL g616 ( 
.A1(n_9),
.A2(n_173),
.B1(n_617),
.B2(n_620),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_10),
.A2(n_158),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_10),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_10),
.A2(n_76),
.B1(n_162),
.B2(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_10),
.A2(n_162),
.B1(n_450),
.B2(n_452),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_10),
.A2(n_162),
.B1(n_462),
.B2(n_465),
.Y(n_461)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_11),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_11),
.A2(n_38),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_11),
.A2(n_38),
.B1(n_128),
.B2(n_433),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_11),
.A2(n_38),
.B1(n_528),
.B2(n_531),
.Y(n_527)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_13),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_13),
.A2(n_94),
.B(n_245),
.Y(n_278)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_13),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_13),
.B(n_80),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_13),
.A2(n_106),
.B1(n_485),
.B2(n_487),
.Y(n_484)
);

OAI32xp33_ASAP7_75t_L g500 ( 
.A1(n_13),
.A2(n_501),
.A3(n_503),
.B1(n_506),
.B2(n_511),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_13),
.A2(n_316),
.B1(n_520),
.B2(n_522),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_14),
.A2(n_148),
.B1(n_151),
.B2(n_155),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_14),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_14),
.A2(n_155),
.B1(n_297),
.B2(n_302),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_14),
.A2(n_155),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_14),
.A2(n_155),
.B1(n_463),
.B2(n_486),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_15),
.A2(n_179),
.B1(n_182),
.B2(n_184),
.Y(n_178)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_15),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_15),
.A2(n_184),
.B1(n_380),
.B2(n_383),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_15),
.A2(n_184),
.B1(n_353),
.B2(n_590),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_15),
.A2(n_184),
.B1(n_629),
.B2(n_633),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_16),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_16),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_16),
.Y(n_222)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_16),
.Y(n_231)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_16),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_16),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_16),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_17),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_21),
.B(n_23),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_19),
.Y(n_150)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_19),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_644),
.B(n_647),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_559),
.B(n_637),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_397),
.B(n_554),
.Y(n_26)
);

NAND3xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_319),
.C(n_361),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_261),
.B(n_289),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_29),
.B(n_261),
.C(n_556),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_164),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_30),
.B(n_165),
.C(n_223),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_82),
.C(n_134),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_31),
.A2(n_134),
.B1(n_135),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_31),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_43),
.B1(n_71),
.B2(n_80),
.Y(n_31)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_32),
.Y(n_276)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_36),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_37),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_42),
.Y(n_143)
);

INVx3_ASAP7_75t_SL g250 ( 
.A(n_43),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_43),
.A2(n_80),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

OAI21xp33_ASAP7_75t_SL g612 ( 
.A1(n_43),
.A2(n_80),
.B(n_613),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_53),
.B(n_59),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g511 ( 
.A(n_44),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_52),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_63),
.Y(n_197)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_63),
.Y(n_214)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_66),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_67),
.Y(n_219)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_67),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_67),
.Y(n_425)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_67),
.Y(n_455)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_71),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_72),
.Y(n_502)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_73),
.Y(n_521)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_78),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_79),
.Y(n_256)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_79),
.Y(n_301)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_79),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_79),
.Y(n_576)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22x1_ASAP7_75t_SL g248 ( 
.A1(n_81),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_81),
.A2(n_250),
.B1(n_269),
.B2(n_276),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_81),
.A2(n_250),
.B1(n_269),
.B2(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_81),
.A2(n_250),
.B1(n_251),
.B2(n_352),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_81),
.A2(n_250),
.B1(n_296),
.B2(n_519),
.Y(n_518)
);

OAI22x1_ASAP7_75t_L g571 ( 
.A1(n_81),
.A2(n_250),
.B1(n_371),
.B2(n_572),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_81),
.A2(n_250),
.B1(n_572),
.B2(n_589),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_82),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_105),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_83),
.B(n_105),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_97),
.B2(n_101),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_90),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_92),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_95),
.Y(n_163)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_96),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_137),
.B(n_142),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_112),
.B1(n_122),
.B2(n_123),
.Y(n_105)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_106),
.A2(n_123),
.B1(n_169),
.B2(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_106),
.A2(n_178),
.B(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_106),
.A2(n_432),
.B1(n_437),
.B2(n_439),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_106),
.A2(n_461),
.B1(n_485),
.B2(n_491),
.Y(n_490)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_107),
.A2(n_167),
.B1(n_460),
.B2(n_469),
.Y(n_459)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_109),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_109),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_110),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_113),
.A2(n_167),
.B1(n_308),
.B2(n_314),
.Y(n_307)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_114),
.Y(n_444)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_114),
.Y(n_486)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g403 ( 
.A1(n_119),
.A2(n_404),
.A3(n_407),
.B1(n_411),
.B2(n_413),
.Y(n_403)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx5_ASAP7_75t_L g436 ( 
.A(n_121),
.Y(n_436)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_127),
.Y(n_419)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_127),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_132),
.Y(n_313)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g243 ( 
.A1(n_136),
.A2(n_156),
.B1(n_157),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_136),
.A2(n_147),
.B1(n_156),
.B2(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_136),
.A2(n_156),
.B1(n_244),
.B2(n_346),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_136),
.A2(n_156),
.B1(n_346),
.B2(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_136),
.A2(n_156),
.B1(n_393),
.B2(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_136),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_136),
.A2(n_156),
.B1(n_615),
.B2(n_616),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_136),
.A2(n_156),
.B1(n_616),
.B2(n_628),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_142),
.A2(n_581),
.B1(n_582),
.B2(n_583),
.Y(n_580)
);

OAI21xp5_ASAP7_75t_SL g645 ( 
.A1(n_142),
.A2(n_582),
.B(n_646),
.Y(n_645)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_143),
.Y(n_591)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_148),
.Y(n_620)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g635 ( 
.A(n_150),
.Y(n_635)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_153),
.Y(n_348)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_153),
.Y(n_350)
);

INVx8_ASAP7_75t_L g586 ( 
.A(n_153),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_156),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_223),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_185),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_166),
.A2(n_186),
.B(n_202),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_174),
.B2(n_177),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_167),
.A2(n_308),
.B1(n_440),
.B2(n_513),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_170),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_175),
.Y(n_491)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_176),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_202),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_194),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_187),
.A2(n_203),
.B1(n_215),
.B2(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_187),
.A2(n_203),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_187),
.A2(n_203),
.B1(n_422),
.B2(n_426),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_187),
.A2(n_203),
.B1(n_426),
.B2(n_449),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_187),
.A2(n_203),
.B1(n_449),
.B2(n_527),
.Y(n_526)
);

OA21x2_ASAP7_75t_L g565 ( 
.A1(n_187),
.A2(n_203),
.B(n_379),
.Y(n_565)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_188),
.A2(n_280),
.B1(n_281),
.B2(n_288),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_188),
.A2(n_195),
.B1(n_280),
.B2(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_188),
.B(n_316),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_188),
.A2(n_280),
.B1(n_281),
.B2(n_544),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_189),
.B(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_201),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_215),
.Y(n_202)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_203),
.Y(n_280)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_209),
.B1(n_212),
.B2(n_214),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_207),
.Y(n_505)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_213),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_221),
.Y(n_429)
);

BUFx12f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_222),
.Y(n_385)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_222),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_222),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_242),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_224),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_237),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_225),
.A2(n_226),
.B1(n_237),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_227),
.Y(n_288)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_231),
.Y(n_334)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_236),
.Y(n_532)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_238),
.Y(n_314)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_238),
.Y(n_513)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_241),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_248),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_243),
.Y(n_322)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_247),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_248),
.B(n_322),
.C(n_323),
.Y(n_321)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_256),
.Y(n_305)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_267),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_262),
.B(n_318),
.Y(n_317)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_267),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_277),
.C(n_279),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_279),
.Y(n_292)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_274),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_277),
.B(n_292),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_317),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_290),
.B(n_317),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.C(n_294),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_291),
.B(n_551),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_293),
.B(n_294),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_306),
.C(n_315),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_295),
.B(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx6_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_304),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_306),
.A2(n_307),
.B1(n_315),
.B2(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_313),
.Y(n_468)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_315),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_316),
.B(n_412),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_SL g422 ( 
.A1(n_316),
.A2(n_411),
.B(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_316),
.B(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_316),
.B(n_507),
.Y(n_506)
);

A2O1A1O1Ixp25_ASAP7_75t_L g554 ( 
.A1(n_319),
.A2(n_361),
.B(n_555),
.C(n_557),
.D(n_558),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_360),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_320),
.B(n_360),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_342),
.B1(n_358),
.B2(n_359),
.Y(n_324)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_325),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_359),
.C(n_396),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_335),
.B1(n_336),
.B2(n_341),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_326),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_336),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_327),
.Y(n_378)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_330),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_334),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_335),
.A2(n_336),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_335),
.A2(n_392),
.B(n_394),
.Y(n_601)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_342),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_364),
.C(n_365),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_351),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_345),
.Y(n_365)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_347),
.Y(n_570)
);

INVx6_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_349),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_350),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_352),
.Y(n_369)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_395),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_362),
.B(n_395),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_363),
.B(n_604),
.C(n_605),
.Y(n_603)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_387),
.Y(n_366)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_367),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_377),
.B(n_386),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_377),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_386),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_386),
.A2(n_597),
.B1(n_600),
.B2(n_608),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_387),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_394),
.Y(n_387)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

AOI21x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_549),
.B(n_553),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_534),
.B(n_548),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_496),
.B(n_533),
.Y(n_399)
);

OAI21x1_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_457),
.B(n_495),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_430),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_402),
.B(n_430),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_420),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_403),
.A2(n_420),
.B1(n_421),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_445),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_431),
.B(n_447),
.C(n_456),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_432),
.Y(n_469)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_448),
.B2(n_456),
.Y(n_445)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_446),
.Y(n_456)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_472),
.B(n_494),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_470),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_459),
.B(n_470),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g472 ( 
.A1(n_473),
.A2(n_489),
.B(n_493),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_484),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_482),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_492),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_497),
.B(n_498),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_516),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_499),
.B(n_517),
.C(n_526),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_512),
.B1(n_514),
.B2(n_515),
.Y(n_499)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_500),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_500),
.B(n_515),
.Y(n_542)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_512),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_517),
.A2(n_518),
.B1(n_525),
.B2(n_526),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_527),
.Y(n_544)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_535),
.B(n_547),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_535),
.B(n_547),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_536),
.A2(n_537),
.B1(n_540),
.B2(n_541),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_536),
.B(n_543),
.C(n_545),
.Y(n_552)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_542),
.A2(n_543),
.B1(n_545),
.B2(n_546),
.Y(n_541)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_542),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_543),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_550),
.B(n_552),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_552),
.Y(n_553)
);

NOR3xp33_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_609),
.C(n_625),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_602),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_562),
.A2(n_640),
.B(n_641),
.Y(n_639)
);

NOR2x1_ASAP7_75t_L g562 ( 
.A(n_563),
.B(n_595),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_563),
.B(n_595),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_578),
.Y(n_563)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_566),
.C(n_571),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_565),
.A2(n_588),
.B1(n_592),
.B2(n_593),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_565),
.Y(n_593)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_565),
.B(n_571),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_565),
.B(n_580),
.C(n_622),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_566),
.A2(n_567),
.B1(n_579),
.B2(n_594),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_566),
.A2(n_567),
.B1(n_598),
.B2(n_599),
.Y(n_597)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_567),
.B(n_579),
.C(n_624),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_568),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_574),
.Y(n_573)
);

INVx6_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx6_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_579),
.Y(n_594)
);

XNOR2x1_ASAP7_75t_L g579 ( 
.A(n_580),
.B(n_587),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_583),
.Y(n_615)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_588),
.Y(n_592)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_589),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_592),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_596),
.B(n_600),
.C(n_601),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_597),
.Y(n_608)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_598),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_601),
.B(n_607),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_606),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_603),
.B(n_606),
.Y(n_640)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

A2O1A1O1Ixp25_ASAP7_75t_L g638 ( 
.A1(n_610),
.A2(n_626),
.B(n_639),
.C(n_642),
.D(n_643),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_623),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_611),
.B(n_623),
.Y(n_642)
);

BUFx24_ASAP7_75t_SL g650 ( 
.A(n_611),
.Y(n_650)
);

FAx1_ASAP7_75t_SL g611 ( 
.A(n_612),
.B(n_614),
.CI(n_621),
.CON(n_611),
.SN(n_611)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_612),
.B(n_614),
.C(n_621),
.Y(n_636)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_627),
.B(n_636),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_627),
.B(n_636),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_627),
.B(n_645),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_645),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_628),
.Y(n_646)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_648),
.Y(n_647)
);


endmodule