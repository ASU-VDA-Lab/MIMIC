module fake_jpeg_29066_n_186 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_186);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_186;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_26),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

BUFx6f_ASAP7_75t_SL g75 ( 
.A(n_69),
.Y(n_75)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_79),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_1),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_51),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_87),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_64),
.B1(n_63),
.B2(n_47),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_93),
.B1(n_54),
.B2(n_72),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_64),
.B1(n_47),
.B2(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_53),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_72),
.Y(n_116)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_97),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_116),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_84),
.A2(n_70),
.B(n_57),
.C(n_62),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_106),
.B(n_21),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_58),
.B(n_49),
.Y(n_106)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_110),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_71),
.B1(n_66),
.B2(n_60),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_48),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_138),
.C(n_22),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_50),
.B1(n_48),
.B2(n_68),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_125),
.B1(n_128),
.B2(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_1),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_134),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_133),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_101),
.A2(n_2),
.B1(n_4),
.B2(n_7),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_14),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_45),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_33),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_17),
.Y(n_138)
);

OA22x2_ASAP7_75t_SL g139 ( 
.A1(n_115),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_35),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_141),
.B(n_28),
.Y(n_156)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_148),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_150),
.C(n_155),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_24),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_154),
.B(n_159),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_44),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_30),
.B(n_31),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_160),
.B(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_151),
.A2(n_119),
.B(n_37),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_165),
.A2(n_151),
.B1(n_142),
.B2(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_152),
.B(n_155),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_173),
.B(n_174),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_177),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_176),
.C(n_175),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_180),
.B(n_162),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_170),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_182),
.B(n_163),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_166),
.A3(n_147),
.B1(n_175),
.B2(n_178),
.C1(n_161),
.C2(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_150),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_169),
.Y(n_186)
);


endmodule