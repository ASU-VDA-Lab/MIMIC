module real_jpeg_28110_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_0),
.A2(n_28),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_21),
.B1(n_23),
.B2(n_28),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_1),
.B(n_21),
.Y(n_42)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_21),
.B1(n_23),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_30),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_96)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_21),
.B1(n_23),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g51 ( 
.A1(n_6),
.A2(n_52),
.B(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_25),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_25),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_6),
.A2(n_41),
.B1(n_45),
.B2(n_103),
.Y(n_106)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_9),
.A2(n_21),
.B1(n_23),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_11),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_78),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_76),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_48),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_15),
.B(n_48),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_31),
.C(n_38),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_16),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_16)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_17),
.A2(n_18),
.B1(n_27),
.B2(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_24),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_18),
.B(n_56),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_18)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

OAI32xp33_ASAP7_75t_L g86 ( 
.A1(n_19),
.A2(n_23),
.A3(n_25),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_20),
.B(n_21),
.Y(n_88)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_21),
.B(n_108),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_25),
.B(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI32xp33_ASAP7_75t_L g68 ( 
.A1(n_26),
.A2(n_36),
.A3(n_52),
.B1(n_55),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_29),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_51),
.B1(n_57),
.B2(n_59),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_36),
.B(n_52),
.C(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_52),
.Y(n_58)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_45),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_41),
.A2(n_43),
.B1(n_45),
.B2(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_41),
.A2(n_45),
.B1(n_96),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_42),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_45),
.B(n_56),
.Y(n_108)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_67),
.B1(n_74),
.B2(n_75),
.Y(n_48)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_92),
.B(n_111),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_89),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_89),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_99)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_100),
.B(n_110),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_99),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_109),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_102),
.B(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);


endmodule