module fake_netlist_6_4242_n_1611 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1611);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1611;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_30),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_2),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_39),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_72),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_27),
.Y(n_160)
);

BUFx10_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_5),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_97),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_74),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_18),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_33),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_15),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_26),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_117),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_71),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_9),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_115),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_33),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_22),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_52),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_80),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_133),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_46),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_38),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_57),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_34),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_17),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_137),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_26),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_20),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_81),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_87),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_100),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_92),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_107),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_67),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_55),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_120),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_136),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_49),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_15),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_96),
.Y(n_214)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_56),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_108),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_3),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_50),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_34),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_16),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_127),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_122),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_88),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_7),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_126),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_44),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_124),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_29),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_48),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_145),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_104),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_51),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_73),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_58),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_78),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_64),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_9),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_4),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_36),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_95),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_47),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_147),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_21),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_19),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_82),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_35),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_62),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_76),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_43),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_60),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_22),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_61),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_99),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_143),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_4),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_106),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_116),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_37),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_21),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_89),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_20),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_42),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_6),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_30),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_119),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_86),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_11),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_68),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_29),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_38),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_23),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_90),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_25),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_70),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_102),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_24),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_103),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_113),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_114),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_75),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_59),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_3),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_125),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_5),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_98),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_151),
.Y(n_303)
);

INVxp33_ASAP7_75t_SL g304 ( 
.A(n_164),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_267),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_189),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_156),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_191),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_152),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_236),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_193),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_221),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_196),
.B(n_0),
.Y(n_314)
);

BUFx10_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_174),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_152),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_174),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_156),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_183),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_183),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_198),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_202),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_271),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_246),
.B(n_1),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_266),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_203),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_175),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_157),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_204),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_209),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_160),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_159),
.Y(n_337)
);

INVxp67_ASAP7_75t_SL g338 ( 
.A(n_223),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_223),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_159),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_180),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_210),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_181),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_186),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_211),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_246),
.B(n_1),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_187),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_188),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_194),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_199),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_200),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_213),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_227),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_231),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_249),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_266),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_212),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_252),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_224),
.B(n_6),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_164),
.Y(n_361)
);

BUFx2_ASAP7_75t_SL g362 ( 
.A(n_185),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_257),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_268),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_185),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_270),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_226),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_228),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_234),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_238),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_240),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_190),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_258),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_247),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_272),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_310),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_305),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_305),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_317),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_358),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_316),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_316),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_333),
.Y(n_387)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_315),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_333),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_318),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_341),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_313),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_341),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_362),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_302),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_339),
.B(n_217),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_303),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_306),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_344),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_315),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_339),
.B(n_158),
.Y(n_405)
);

OAI21x1_ASAP7_75t_L g406 ( 
.A1(n_328),
.A2(n_299),
.B(n_155),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_315),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_361),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_258),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_348),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_308),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_348),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_312),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_329),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_323),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_346),
.A2(n_299),
.B(n_162),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_352),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_307),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_352),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_325),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_330),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_334),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_374),
.B(n_265),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_314),
.B(n_304),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_335),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_320),
.B(n_322),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_354),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_342),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_320),
.B(n_265),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_345),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

CKINVDCx11_ASAP7_75t_R g446 ( 
.A(n_377),
.Y(n_446)
);

BUFx10_ASAP7_75t_L g447 ( 
.A(n_436),
.Y(n_447)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

NOR2x1p5_ASAP7_75t_L g450 ( 
.A(n_399),
.B(n_311),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_357),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_400),
.B(n_359),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_388),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_411),
.B(n_153),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_411),
.B(n_322),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_435),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_421),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_377),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_417),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_438),
.Y(n_461)
);

INVxp33_ASAP7_75t_L g462 ( 
.A(n_398),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_400),
.B(n_365),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_438),
.Y(n_464)
);

INVxp33_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

BUFx6f_ASAP7_75t_SL g466 ( 
.A(n_416),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_380),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_405),
.B(n_153),
.Y(n_468)
);

AND2x6_ASAP7_75t_L g469 ( 
.A(n_411),
.B(n_153),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_380),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_389),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_404),
.B(n_368),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_435),
.B(n_404),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_382),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_435),
.B(n_376),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_416),
.B(n_369),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_414),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_435),
.A2(n_442),
.B1(n_424),
.B2(n_406),
.Y(n_484)
);

AND2x6_ASAP7_75t_L g485 ( 
.A(n_435),
.B(n_153),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_417),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_404),
.B(n_370),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_408),
.B(n_414),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_381),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_327),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_427),
.B(n_332),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_383),
.Y(n_493)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_427),
.B(n_405),
.C(n_410),
.Y(n_494)
);

OR2x6_ASAP7_75t_L g495 ( 
.A(n_416),
.B(n_362),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_383),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_408),
.B(n_371),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_416),
.B(n_372),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_412),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_381),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_383),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_414),
.B(n_163),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_383),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_416),
.B(n_360),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_417),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_417),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_402),
.B(n_375),
.Y(n_508)
);

AND3x2_ASAP7_75t_L g509 ( 
.A(n_382),
.B(n_173),
.C(n_356),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_383),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_413),
.A2(n_326),
.B1(n_251),
.B2(n_237),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_414),
.B(n_376),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_442),
.B(n_364),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_383),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_415),
.B(n_419),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_415),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_419),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_386),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_421),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_386),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_408),
.B(n_248),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_386),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_410),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_397),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_386),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_445),
.B(n_163),
.Y(n_530)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_406),
.A2(n_215),
.B1(n_292),
.B2(n_300),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_386),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_406),
.A2(n_215),
.B1(n_278),
.B2(n_274),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_425),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_425),
.B(n_163),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_426),
.B(n_327),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_424),
.B(n_363),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_423),
.B(n_343),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_386),
.Y(n_540)
);

BUFx10_ASAP7_75t_L g541 ( 
.A(n_429),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_386),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_433),
.B(n_307),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_425),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_390),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_397),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_390),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_390),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_424),
.B(n_321),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_425),
.B(n_163),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_418),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_434),
.B(n_219),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_321),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_390),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_431),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_441),
.A2(n_237),
.B1(n_251),
.B2(n_244),
.Y(n_559)
);

BUFx2_ASAP7_75t_L g560 ( 
.A(n_395),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_390),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_432),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_432),
.B(n_367),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_395),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_418),
.B(n_219),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_418),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_418),
.B(n_254),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_L g568 ( 
.A(n_444),
.B(n_331),
.C(n_277),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_443),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_418),
.Y(n_570)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_445),
.B(n_331),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_445),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_384),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_384),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_453),
.B(n_158),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_516),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_451),
.B(n_241),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_SL g578 ( 
.A(n_512),
.B(n_340),
.C(n_337),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_463),
.B(n_165),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

O2A1O1Ixp33_ASAP7_75t_L g581 ( 
.A1(n_452),
.A2(n_445),
.B(n_440),
.C(n_439),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_539),
.B(n_165),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_491),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_505),
.B(n_167),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_566),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_494),
.B(n_167),
.Y(n_586)
);

OR2x6_ASAP7_75t_L g587 ( 
.A(n_560),
.B(n_273),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_481),
.B(n_378),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_558),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_558),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_481),
.B(n_379),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_573),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_505),
.A2(n_262),
.B1(n_192),
.B2(n_184),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_526),
.B(n_367),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_483),
.B(n_379),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_562),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_482),
.B(n_170),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_562),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_170),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_478),
.A2(n_179),
.B1(n_205),
.B2(n_206),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_574),
.Y(n_601)
);

O2A1O1Ixp5_ASAP7_75t_L g602 ( 
.A1(n_478),
.A2(n_269),
.B(n_208),
.C(n_207),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_552),
.A2(n_197),
.B1(n_243),
.B2(n_295),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_456),
.B(n_177),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_456),
.B(n_177),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_574),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_513),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_554),
.B(n_219),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

INVxp67_ASAP7_75t_R g610 ( 
.A(n_564),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_461),
.B(n_178),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_526),
.B(n_366),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_464),
.B(n_178),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_467),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_513),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_552),
.A2(n_243),
.B1(n_197),
.B2(n_149),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_499),
.B(n_233),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

NOR3xp33_ASAP7_75t_L g619 ( 
.A(n_559),
.B(n_222),
.C(n_229),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_514),
.B(n_233),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_446),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_466),
.A2(n_373),
.B1(n_256),
.B2(n_260),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_473),
.B(n_487),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_497),
.B(n_440),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_470),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_472),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_555),
.B(n_281),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_555),
.B(n_286),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_514),
.B(n_286),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_514),
.B(n_545),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_556),
.B(n_288),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_447),
.B(n_288),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_476),
.B(n_477),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_480),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_491),
.B(n_393),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_470),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_448),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_489),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_479),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_548),
.B(n_290),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_495),
.B(n_166),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_448),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_479),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_447),
.B(n_290),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_447),
.B(n_492),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_500),
.B(n_439),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_517),
.B(n_294),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_518),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_519),
.B(n_525),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_479),
.B(n_161),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_532),
.B(n_394),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_543),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_537),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_484),
.A2(n_534),
.B1(n_531),
.B2(n_538),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_459),
.B(n_171),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_571),
.A2(n_428),
.B(n_409),
.C(n_403),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_554),
.B(n_279),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_SL g658 ( 
.A(n_541),
.B(n_161),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_541),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_541),
.Y(n_660)
);

AND2x4_ASAP7_75t_SL g661 ( 
.A(n_495),
.B(n_161),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_537),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_466),
.A2(n_264),
.B1(n_261),
.B2(n_297),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_508),
.B(n_294),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_552),
.A2(n_538),
.B1(n_469),
.B2(n_455),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_568),
.B(n_296),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_475),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_527),
.B(n_396),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_548),
.B(n_296),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_572),
.B(n_428),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_488),
.A2(n_225),
.B(n_230),
.C(n_235),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_462),
.B(n_396),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_572),
.B(n_409),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_547),
.Y(n_675)
);

BUFx2_ASAP7_75t_L g676 ( 
.A(n_490),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_547),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_462),
.B(n_275),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_550),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_550),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_552),
.A2(n_168),
.B1(n_301),
.B2(n_169),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_465),
.B(n_154),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_501),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_446),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_563),
.Y(n_685)
);

AO221x1_ASAP7_75t_L g686 ( 
.A1(n_449),
.A2(n_279),
.B1(n_176),
.B2(n_182),
.C(n_195),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_572),
.B(n_403),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_458),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_563),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_523),
.B(n_567),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_563),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_455),
.B(n_469),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_465),
.B(n_276),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_557),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_469),
.B(n_409),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_557),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_561),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_469),
.B(n_255),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_450),
.B(n_392),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_521),
.B(n_232),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_469),
.B(n_488),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_538),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_485),
.B(n_454),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_538),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_495),
.A2(n_284),
.B1(n_216),
.B2(n_201),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_536),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_493),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_485),
.A2(n_468),
.B1(n_530),
.B2(n_553),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_577),
.B(n_474),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_675),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_SL g712 ( 
.A1(n_690),
.A2(n_536),
.B(n_553),
.C(n_524),
.Y(n_712)
);

OAI21xp33_ASAP7_75t_L g713 ( 
.A1(n_577),
.A2(n_280),
.B(n_172),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_654),
.A2(n_496),
.B(n_493),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_656),
.A2(n_496),
.B(n_504),
.Y(n_715)
);

O2A1O1Ixp33_ASAP7_75t_SL g716 ( 
.A1(n_623),
.A2(n_593),
.B(n_702),
.C(n_579),
.Y(n_716)
);

AND2x2_ASAP7_75t_SL g717 ( 
.A(n_603),
.B(n_468),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_635),
.Y(n_718)
);

NOR2x1_ASAP7_75t_L g719 ( 
.A(n_639),
.B(n_474),
.Y(n_719)
);

AOI21x1_ASAP7_75t_L g720 ( 
.A1(n_608),
.A2(n_533),
.B(n_522),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_671),
.A2(n_687),
.B(n_674),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_584),
.A2(n_583),
.B(n_580),
.C(n_576),
.Y(n_722)
);

O2A1O1Ixp5_ASAP7_75t_L g723 ( 
.A1(n_575),
.A2(n_608),
.B(n_657),
.C(n_602),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_635),
.Y(n_724)
);

AO21x1_ASAP7_75t_L g725 ( 
.A1(n_703),
.A2(n_565),
.B(n_503),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_598),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_R g727 ( 
.A(n_688),
.B(n_521),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_578),
.B(n_253),
.C(n_263),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_598),
.Y(n_729)
);

BUFx8_ASAP7_75t_L g730 ( 
.A(n_676),
.Y(n_730)
);

INVx5_ASAP7_75t_L g731 ( 
.A(n_641),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_598),
.Y(n_732)
);

AO22x1_ASAP7_75t_L g733 ( 
.A1(n_665),
.A2(n_171),
.B1(n_172),
.B2(n_280),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_630),
.A2(n_503),
.B(n_565),
.C(n_498),
.Y(n_734)
);

AOI21xp5_ASAP7_75t_L g735 ( 
.A1(n_704),
.A2(n_535),
.B(n_486),
.Y(n_735)
);

AOI22x1_ASAP7_75t_L g736 ( 
.A1(n_707),
.A2(n_504),
.B1(n_502),
.B2(n_544),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_621),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_705),
.B(n_529),
.C(n_502),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_675),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_643),
.Y(n_740)
);

BUFx12f_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

BUFx12f_ASAP7_75t_L g742 ( 
.A(n_637),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_673),
.B(n_669),
.Y(n_743)
);

NAND2x1p5_ASAP7_75t_L g744 ( 
.A(n_607),
.B(n_609),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_615),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_509),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_665),
.B(n_632),
.Y(n_747)
);

NAND3xp33_ASAP7_75t_L g748 ( 
.A(n_681),
.B(n_515),
.C(n_510),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_677),
.Y(n_749)
);

CKINVDCx8_ASAP7_75t_R g750 ( 
.A(n_587),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_581),
.A2(n_520),
.B(n_510),
.Y(n_751)
);

AOI21x1_ASAP7_75t_L g752 ( 
.A1(n_657),
.A2(n_520),
.B(n_524),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_627),
.A2(n_522),
.B(n_529),
.C(n_544),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_677),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_653),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_604),
.B(n_485),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_685),
.A2(n_528),
.B1(n_546),
.B2(n_542),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_639),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_604),
.B(n_605),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_588),
.A2(n_540),
.B(n_570),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_591),
.A2(n_540),
.B(n_570),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_595),
.A2(n_570),
.B(n_546),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_659),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_605),
.B(n_506),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_633),
.A2(n_570),
.B(n_546),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_649),
.A2(n_542),
.B(n_449),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_692),
.A2(n_279),
.B1(n_528),
.B2(n_511),
.Y(n_767)
);

A2O1A1Ixp33_ASAP7_75t_L g768 ( 
.A1(n_627),
.A2(n_507),
.B(n_506),
.C(n_460),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_642),
.B(n_232),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_594),
.B(n_283),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_660),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_663),
.B(n_232),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_640),
.B(n_218),
.C(n_239),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_646),
.A2(n_385),
.B(n_384),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_618),
.B(n_385),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_679),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_585),
.A2(n_283),
.B(n_291),
.C(n_289),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_666),
.A2(n_530),
.B(n_298),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_666),
.A2(n_259),
.B1(n_245),
.B2(n_250),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_680),
.A2(n_530),
.B(n_242),
.Y(n_780)
);

AND2x2_ASAP7_75t_SL g781 ( 
.A(n_603),
.B(n_285),
.Y(n_781)
);

AO21x2_ASAP7_75t_L g782 ( 
.A1(n_686),
.A2(n_530),
.B(n_63),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_626),
.B(n_291),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_638),
.B(n_289),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_680),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_589),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_700),
.B(n_285),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_648),
.B(n_8),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_645),
.A2(n_144),
.B1(n_142),
.B2(n_134),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_652),
.B(n_8),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_691),
.Y(n_791)
);

AOI21x1_ASAP7_75t_L g792 ( 
.A1(n_651),
.A2(n_131),
.B(n_129),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_632),
.B(n_11),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_695),
.Y(n_794)
);

BUFx4f_ASAP7_75t_L g795 ( 
.A(n_641),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_698),
.A2(n_91),
.B(n_84),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_698),
.A2(n_83),
.B(n_69),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_634),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_683),
.Y(n_799)
);

BUFx12f_ASAP7_75t_L g800 ( 
.A(n_587),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_592),
.A2(n_65),
.B(n_13),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_697),
.A2(n_12),
.B(n_13),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_644),
.B(n_12),
.Y(n_803)
);

OR2x6_ASAP7_75t_SL g804 ( 
.A(n_655),
.B(n_14),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_662),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_708),
.A2(n_16),
.B(n_18),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_696),
.A2(n_19),
.B(n_24),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_600),
.A2(n_25),
.B(n_28),
.C(n_31),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_31),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_693),
.A2(n_36),
.B(n_37),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_645),
.B(n_631),
.Y(n_811)
);

OR2x6_ASAP7_75t_SL g812 ( 
.A(n_616),
.B(n_39),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_611),
.B(n_40),
.Y(n_813)
);

AND2x2_ASAP7_75t_SL g814 ( 
.A(n_616),
.B(n_40),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_SL g815 ( 
.A(n_650),
.B(n_45),
.Y(n_815)
);

INVx11_ASAP7_75t_L g816 ( 
.A(n_610),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_612),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_611),
.B(n_41),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_628),
.A2(n_619),
.B1(n_586),
.B2(n_667),
.Y(n_819)
);

AOI21x1_ASAP7_75t_L g820 ( 
.A1(n_601),
.A2(n_614),
.B(n_668),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_628),
.A2(n_667),
.B1(n_596),
.B2(n_590),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_586),
.A2(n_617),
.B1(n_597),
.B2(n_613),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_613),
.B(n_599),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_620),
.A2(n_629),
.B(n_582),
.C(n_706),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_606),
.Y(n_825)
);

AOI21x1_ASAP7_75t_L g826 ( 
.A1(n_606),
.A2(n_625),
.B(n_636),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_641),
.A2(n_709),
.B1(n_599),
.B2(n_661),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_647),
.B(n_668),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_664),
.B(n_622),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_587),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_709),
.A2(n_661),
.B1(n_647),
.B2(n_682),
.Y(n_831)
);

A2O1A1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_682),
.A2(n_672),
.B(n_699),
.C(n_658),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_670),
.B(n_678),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_694),
.B(n_701),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_577),
.A2(n_623),
.B(n_627),
.C(n_628),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_635),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_594),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_SL g838 ( 
.A(n_577),
.B(n_466),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_635),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_634),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_594),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_577),
.B(n_623),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_577),
.B(n_623),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_676),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_577),
.B(n_451),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_635),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_583),
.B(n_689),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_639),
.B(n_659),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_598),
.B(n_577),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_577),
.B(n_623),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_624),
.A2(n_457),
.B(n_478),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_654),
.A2(n_577),
.B1(n_623),
.B2(n_681),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_577),
.B(n_451),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_624),
.A2(n_457),
.B(n_478),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_577),
.A2(n_623),
.B1(n_654),
.B2(n_463),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_598),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_577),
.B(n_451),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_621),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_842),
.B(n_843),
.Y(n_859)
);

AO31x2_ASAP7_75t_L g860 ( 
.A1(n_725),
.A2(n_753),
.A3(n_852),
.B(n_768),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_743),
.B(n_770),
.Y(n_861)
);

OAI21x1_ASAP7_75t_L g862 ( 
.A1(n_720),
.A2(n_752),
.B(n_820),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_850),
.B(n_845),
.Y(n_863)
);

AO31x2_ASAP7_75t_L g864 ( 
.A1(n_835),
.A2(n_831),
.A3(n_832),
.B(n_809),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_726),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_853),
.A2(n_857),
.B(n_747),
.C(n_855),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_837),
.B(n_841),
.Y(n_867)
);

NOR3xp33_ASAP7_75t_L g868 ( 
.A(n_759),
.B(n_823),
.C(n_834),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_805),
.Y(n_869)
);

AOI21xp33_ASAP7_75t_L g870 ( 
.A1(n_819),
.A2(n_818),
.B(n_813),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_844),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_826),
.A2(n_736),
.B(n_751),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_828),
.B(n_822),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_724),
.B(n_811),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_749),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_825),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_833),
.A2(n_793),
.B1(n_803),
.B2(n_829),
.Y(n_877)
);

OAI21x1_ASAP7_75t_SL g878 ( 
.A1(n_801),
.A2(n_797),
.B(n_796),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_798),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_724),
.B(n_764),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_851),
.A2(n_854),
.B(n_721),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_840),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_715),
.A2(n_714),
.B(n_735),
.Y(n_883)
);

AO21x1_ASAP7_75t_L g884 ( 
.A1(n_801),
.A2(n_806),
.B(n_802),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_824),
.A2(n_722),
.B(n_821),
.C(n_717),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_726),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_SL g887 ( 
.A1(n_827),
.A2(n_797),
.B(n_796),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_716),
.A2(n_710),
.B(n_756),
.Y(n_888)
);

AO21x1_ASAP7_75t_L g889 ( 
.A1(n_838),
.A2(n_849),
.B(n_810),
.Y(n_889)
);

OAI21xp5_ASAP7_75t_L g890 ( 
.A1(n_748),
.A2(n_723),
.B(n_738),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_755),
.B(n_814),
.Y(n_891)
);

BUFx4f_ASAP7_75t_SL g892 ( 
.A(n_742),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_726),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_718),
.B(n_836),
.Y(n_894)
);

OAI21x1_ASAP7_75t_L g895 ( 
.A1(n_766),
.A2(n_761),
.B(n_760),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_754),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_SL g897 ( 
.A1(n_745),
.A2(n_790),
.B(n_788),
.Y(n_897)
);

OAI21x1_ASAP7_75t_L g898 ( 
.A1(n_762),
.A2(n_774),
.B(n_765),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_776),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_840),
.B(n_799),
.Y(n_900)
);

OAI21x1_ASAP7_75t_L g901 ( 
.A1(n_734),
.A2(n_711),
.B(n_739),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_817),
.B(n_781),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_839),
.B(n_846),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_785),
.A2(n_794),
.B(n_791),
.Y(n_904)
);

NAND2x1_ASAP7_75t_L g905 ( 
.A(n_729),
.B(n_856),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_780),
.A2(n_712),
.B(n_748),
.Y(n_906)
);

NAND2x1_ASAP7_75t_L g907 ( 
.A(n_729),
.B(n_856),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_730),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_713),
.B(n_755),
.Y(n_909)
);

OAI222xp33_ASAP7_75t_L g910 ( 
.A1(n_779),
.A2(n_812),
.B1(n_808),
.B2(n_789),
.C1(n_750),
.C2(n_807),
.Y(n_910)
);

AOI21xp33_ASAP7_75t_L g911 ( 
.A1(n_838),
.A2(n_775),
.B(n_778),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_847),
.B(n_755),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_729),
.Y(n_913)
);

OAI21x1_ASAP7_75t_L g914 ( 
.A1(n_744),
.A2(n_757),
.B(n_792),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_732),
.B(n_786),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_767),
.A2(n_778),
.B(n_783),
.Y(n_916)
);

OR2x6_ASAP7_75t_SL g917 ( 
.A(n_740),
.B(n_784),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_786),
.B(n_847),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_786),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_856),
.B(n_719),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_L g921 ( 
.A(n_815),
.B(n_728),
.C(n_733),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_787),
.B(n_773),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_795),
.A2(n_731),
.B1(n_848),
.B2(n_830),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_758),
.B(n_746),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_731),
.B(n_758),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_772),
.A2(n_769),
.B(n_777),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_795),
.A2(n_746),
.B(n_815),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_758),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_848),
.A2(n_804),
.B1(n_763),
.B2(n_771),
.Y(n_929)
);

NAND2x1_ASAP7_75t_L g930 ( 
.A(n_763),
.B(n_816),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_741),
.B(n_800),
.Y(n_931)
);

AOI21xp33_ASAP7_75t_L g932 ( 
.A1(n_782),
.A2(n_730),
.B(n_737),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_858),
.A2(n_852),
.B(n_855),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_727),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_727),
.Y(n_935)
);

OAI22x1_ASAP7_75t_L g936 ( 
.A1(n_845),
.A2(n_853),
.B1(n_857),
.B2(n_747),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_726),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_720),
.A2(n_752),
.B(n_820),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_825),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_851),
.A2(n_854),
.B(n_654),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_851),
.A2(n_854),
.B(n_654),
.Y(n_941)
);

AND2x2_ASAP7_75t_SL g942 ( 
.A(n_814),
.B(n_853),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_845),
.B(n_853),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_805),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_845),
.B(n_853),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_743),
.B(n_847),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_726),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_844),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_852),
.A2(n_855),
.B(n_714),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_740),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_840),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_842),
.B(n_843),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_842),
.B(n_843),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_726),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_842),
.B(n_843),
.Y(n_955)
);

AOI221x1_ASAP7_75t_L g956 ( 
.A1(n_845),
.A2(n_853),
.B1(n_857),
.B2(n_747),
.C(n_852),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_726),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_805),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_842),
.B(n_843),
.Y(n_959)
);

AO21x1_ASAP7_75t_L g960 ( 
.A1(n_852),
.A2(n_747),
.B(n_845),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_743),
.B(n_770),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_743),
.B(n_770),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_720),
.A2(n_752),
.B(n_820),
.Y(n_963)
);

NAND2x1p5_ASAP7_75t_L g964 ( 
.A(n_724),
.B(n_726),
.Y(n_964)
);

NOR2x1_ASAP7_75t_SL g965 ( 
.A(n_726),
.B(n_729),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_720),
.A2(n_752),
.B(n_820),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_842),
.B(n_843),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_845),
.A2(n_857),
.B(n_853),
.C(n_747),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_845),
.B(n_853),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_726),
.Y(n_970)
);

BUFx6f_ASAP7_75t_SL g971 ( 
.A(n_771),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_852),
.A2(n_855),
.B(n_714),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_825),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_805),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_842),
.B(n_843),
.Y(n_975)
);

OAI21x1_ASAP7_75t_SL g976 ( 
.A1(n_801),
.A2(n_797),
.B(n_796),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_743),
.B(n_847),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_845),
.A2(n_857),
.B(n_853),
.C(n_747),
.Y(n_978)
);

BUFx2_ASAP7_75t_R g979 ( 
.A(n_812),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_851),
.A2(n_854),
.B(n_654),
.Y(n_980)
);

AND2x2_ASAP7_75t_SL g981 ( 
.A(n_814),
.B(n_853),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_943),
.B(n_863),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_863),
.B(n_968),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_951),
.B(n_871),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_912),
.B(n_946),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_882),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_869),
.Y(n_987)
);

CKINVDCx16_ASAP7_75t_R g988 ( 
.A(n_950),
.Y(n_988)
);

O2A1O1Ixp5_ASAP7_75t_L g989 ( 
.A1(n_978),
.A2(n_960),
.B(n_884),
.C(n_870),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_942),
.A2(n_981),
.B1(n_936),
.B2(n_945),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_944),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_887),
.A2(n_881),
.B(n_949),
.Y(n_992)
);

O2A1O1Ixp5_ASAP7_75t_SL g993 ( 
.A1(n_870),
.A2(n_932),
.B(n_911),
.C(n_972),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_958),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_859),
.B(n_952),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_951),
.B(n_930),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_969),
.A2(n_933),
.B1(n_921),
.B2(n_877),
.Y(n_997)
);

HB1xp67_ASAP7_75t_L g998 ( 
.A(n_879),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_866),
.B(n_946),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_897),
.B(n_873),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_933),
.A2(n_902),
.B1(n_972),
.B2(n_949),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_977),
.B(n_925),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_859),
.B(n_952),
.Y(n_1003)
);

INVx2_ASAP7_75t_SL g1004 ( 
.A(n_867),
.Y(n_1004)
);

INVx3_ASAP7_75t_SL g1005 ( 
.A(n_935),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_974),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_L g1007 ( 
.A(n_868),
.B(n_953),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_875),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_948),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_896),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_913),
.B(n_954),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_953),
.B(n_955),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_893),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_885),
.A2(n_975),
.B(n_967),
.C(n_955),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_899),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_861),
.B(n_961),
.Y(n_1016)
);

INVx2_ASAP7_75t_SL g1017 ( 
.A(n_950),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_891),
.A2(n_977),
.B1(n_976),
.B2(n_878),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_959),
.A2(n_967),
.B1(n_975),
.B2(n_873),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_893),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_962),
.A2(n_927),
.B1(n_959),
.B2(n_909),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_927),
.A2(n_922),
.B1(n_911),
.B2(n_874),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_893),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_971),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_900),
.Y(n_1025)
);

INVx3_ASAP7_75t_SL g1026 ( 
.A(n_924),
.Y(n_1026)
);

INVx6_ASAP7_75t_L g1027 ( 
.A(n_924),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_916),
.A2(n_922),
.B(n_874),
.C(n_926),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_908),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_894),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_L g1031 ( 
.A(n_956),
.B(n_916),
.C(n_980),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_894),
.Y(n_1032)
);

CKINVDCx8_ASAP7_75t_R g1033 ( 
.A(n_924),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_903),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_970),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_918),
.Y(n_1036)
);

OAI21xp33_ASAP7_75t_L g1037 ( 
.A1(n_979),
.A2(n_903),
.B(n_934),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_918),
.B(n_979),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_929),
.A2(n_923),
.B1(n_880),
.B2(n_924),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_971),
.Y(n_1040)
);

INVx5_ASAP7_75t_L g1041 ( 
.A(n_970),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_928),
.B(n_919),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_929),
.A2(n_923),
.B1(n_880),
.B2(n_889),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_925),
.B(n_915),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_892),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_876),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_864),
.B(n_915),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_917),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_905),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_865),
.Y(n_1050)
);

AND2x6_ASAP7_75t_L g1051 ( 
.A(n_865),
.B(n_886),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_864),
.B(n_920),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_940),
.A2(n_941),
.B(n_906),
.C(n_883),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_864),
.B(n_920),
.Y(n_1054)
);

AOI222xp33_ASAP7_75t_L g1055 ( 
.A1(n_910),
.A2(n_931),
.B1(n_890),
.B2(n_939),
.C1(n_973),
.C2(n_965),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_932),
.A2(n_964),
.B1(n_937),
.B2(n_957),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_890),
.B(n_947),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_886),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_913),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_937),
.B(n_957),
.Y(n_1060)
);

INVx4_ASAP7_75t_L g1061 ( 
.A(n_954),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_907),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_947),
.B(n_860),
.Y(n_1063)
);

INVxp67_ASAP7_75t_L g1064 ( 
.A(n_904),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_901),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_914),
.A2(n_895),
.B(n_898),
.C(n_862),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_938),
.B(n_966),
.Y(n_1067)
);

CKINVDCx11_ASAP7_75t_R g1068 ( 
.A(n_963),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_887),
.A2(n_881),
.B(n_949),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_950),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_871),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_887),
.A2(n_881),
.B(n_949),
.Y(n_1072)
);

BUFx4f_ASAP7_75t_L g1073 ( 
.A(n_924),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_893),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_890),
.A2(n_872),
.B(n_888),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_943),
.B(n_863),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_943),
.A2(n_968),
.B1(n_978),
.B2(n_866),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_951),
.B(n_871),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_968),
.A2(n_853),
.B(n_857),
.C(n_845),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_869),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_SL g1081 ( 
.A(n_950),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_943),
.B(n_863),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_968),
.A2(n_853),
.B(n_857),
.C(n_845),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_871),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_887),
.A2(n_881),
.B(n_949),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_882),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_887),
.A2(n_881),
.B(n_949),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_912),
.B(n_946),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_871),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_887),
.A2(n_881),
.B(n_949),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_964),
.Y(n_1091)
);

HB1xp67_ASAP7_75t_L g1092 ( 
.A(n_951),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_893),
.Y(n_1093)
);

OR2x2_ASAP7_75t_L g1094 ( 
.A(n_863),
.B(n_459),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_951),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_943),
.B(n_942),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_863),
.B(n_459),
.Y(n_1097)
);

OAI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_943),
.A2(n_845),
.B1(n_857),
.B2(n_853),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_968),
.A2(n_853),
.B(n_857),
.C(n_845),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_943),
.B(n_863),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_871),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_869),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_871),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_943),
.B(n_863),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_943),
.A2(n_845),
.B1(n_857),
.B2(n_853),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_943),
.B(n_845),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_893),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_943),
.B(n_853),
.C(n_845),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_871),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_943),
.A2(n_845),
.B(n_857),
.C(n_853),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_871),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_869),
.Y(n_1112)
);

HB1xp67_ASAP7_75t_L g1113 ( 
.A(n_951),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_893),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1059),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_1073),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1109),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_SL g1118 ( 
.A1(n_1106),
.A2(n_1108),
.B1(n_1077),
.B2(n_1096),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1108),
.A2(n_1077),
.B1(n_1098),
.B2(n_1076),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_987),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1092),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_1113),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_991),
.Y(n_1123)
);

CKINVDCx11_ASAP7_75t_R g1124 ( 
.A(n_1029),
.Y(n_1124)
);

BUFx6f_ASAP7_75t_L g1125 ( 
.A(n_1073),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1095),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1006),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_1033),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1105),
.B(n_1110),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1105),
.B(n_1082),
.Y(n_1130)
);

AO21x1_ASAP7_75t_L g1131 ( 
.A1(n_1079),
.A2(n_1099),
.B(n_1083),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1100),
.B(n_1104),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1112),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1094),
.B(n_1097),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1065),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1003),
.A2(n_1012),
.B1(n_982),
.B2(n_995),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_984),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_994),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1001),
.B(n_983),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_1095),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_1004),
.B(n_1017),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_982),
.A2(n_995),
.B1(n_1025),
.B2(n_1019),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1080),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_990),
.A2(n_1021),
.B1(n_997),
.B2(n_1039),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1102),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1008),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_SL g1147 ( 
.A1(n_1038),
.A2(n_1081),
.B1(n_1069),
.B2(n_1072),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1010),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_992),
.A2(n_1085),
.B(n_1087),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1071),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1019),
.B(n_1030),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1015),
.Y(n_1152)
);

BUFx8_ASAP7_75t_L g1153 ( 
.A(n_1081),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1007),
.A2(n_999),
.B1(n_1022),
.B2(n_1000),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_SL g1155 ( 
.A1(n_1090),
.A2(n_1048),
.B1(n_988),
.B2(n_1016),
.Y(n_1155)
);

HB1xp67_ASAP7_75t_L g1156 ( 
.A(n_986),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1046),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1042),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1063),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1036),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1032),
.B(n_1034),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1057),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_1067),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1014),
.B(n_1044),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1089),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1052),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_998),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1009),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_1047),
.B(n_1054),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1031),
.A2(n_1037),
.B1(n_1018),
.B2(n_1055),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1078),
.B(n_1002),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1026),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1075),
.Y(n_1173)
);

AOI222xp33_ASAP7_75t_L g1174 ( 
.A1(n_1037),
.A2(n_985),
.B1(n_1088),
.B2(n_1002),
.C1(n_1031),
.C2(n_1086),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1055),
.A2(n_1044),
.B1(n_1043),
.B2(n_1039),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1060),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1058),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_1041),
.B(n_1074),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1043),
.A2(n_1056),
.B1(n_1027),
.B2(n_996),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_989),
.B(n_1028),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_985),
.B(n_1088),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1084),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1091),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1064),
.Y(n_1184)
);

AO21x1_ASAP7_75t_L g1185 ( 
.A1(n_993),
.A2(n_1035),
.B(n_1011),
.Y(n_1185)
);

BUFx10_ASAP7_75t_L g1186 ( 
.A(n_1024),
.Y(n_1186)
);

OA21x2_ASAP7_75t_L g1187 ( 
.A1(n_1053),
.A2(n_1066),
.B(n_1068),
.Y(n_1187)
);

AOI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1051),
.A2(n_1074),
.B(n_1035),
.Y(n_1188)
);

NOR2x1_ASAP7_75t_SL g1189 ( 
.A(n_1074),
.B(n_1070),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1051),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1051),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1013),
.Y(n_1192)
);

NAND2x1p5_ASAP7_75t_L g1193 ( 
.A(n_1061),
.B(n_1114),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1013),
.Y(n_1194)
);

BUFx10_ASAP7_75t_L g1195 ( 
.A(n_1040),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1101),
.Y(n_1196)
);

OAI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1103),
.A2(n_1111),
.B(n_1045),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1020),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1005),
.B(n_1050),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1020),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1023),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_1023),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1049),
.A2(n_1062),
.B(n_1093),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1107),
.Y(n_1204)
);

BUFx6f_ASAP7_75t_L g1205 ( 
.A(n_1114),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1114),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1049),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1062),
.A2(n_943),
.B1(n_1105),
.B2(n_845),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1001),
.B(n_983),
.Y(n_1209)
);

NAND2x1p5_ASAP7_75t_L g1210 ( 
.A(n_1073),
.B(n_999),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1109),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1073),
.Y(n_1212)
);

AO21x1_ASAP7_75t_L g1213 ( 
.A1(n_1098),
.A2(n_853),
.B(n_845),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_1073),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1098),
.A2(n_943),
.B1(n_853),
.B2(n_857),
.Y(n_1215)
);

HB1xp67_ASAP7_75t_L g1216 ( 
.A(n_1092),
.Y(n_1216)
);

BUFx2_ASAP7_75t_R g1217 ( 
.A(n_1045),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1024),
.Y(n_1218)
);

OR2x2_ASAP7_75t_L g1219 ( 
.A(n_1094),
.B(n_1097),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1106),
.B(n_943),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1106),
.B(n_943),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1092),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1073),
.B(n_999),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_1059),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1151),
.B(n_1136),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1210),
.Y(n_1226)
);

INVxp67_ASAP7_75t_R g1227 ( 
.A(n_1198),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1135),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1169),
.B(n_1166),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1126),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1169),
.B(n_1159),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1163),
.Y(n_1232)
);

BUFx4f_ASAP7_75t_SL g1233 ( 
.A(n_1200),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1163),
.Y(n_1234)
);

AO21x2_ASAP7_75t_L g1235 ( 
.A1(n_1149),
.A2(n_1142),
.B(n_1180),
.Y(n_1235)
);

INVx4_ASAP7_75t_L g1236 ( 
.A(n_1212),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1173),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1139),
.B(n_1209),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1184),
.Y(n_1239)
);

BUFx4f_ASAP7_75t_SL g1240 ( 
.A(n_1200),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1140),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1139),
.B(n_1209),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1162),
.B(n_1142),
.Y(n_1243)
);

OR2x2_ASAP7_75t_L g1244 ( 
.A(n_1164),
.B(n_1175),
.Y(n_1244)
);

BUFx4f_ASAP7_75t_L g1245 ( 
.A(n_1210),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1129),
.B(n_1175),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1223),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1129),
.B(n_1138),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1121),
.Y(n_1249)
);

OR2x6_ASAP7_75t_L g1250 ( 
.A(n_1187),
.B(n_1223),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1119),
.B(n_1118),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1143),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1130),
.B(n_1161),
.Y(n_1253)
);

INVxp33_ASAP7_75t_L g1254 ( 
.A(n_1168),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1122),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1145),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1146),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1148),
.Y(n_1258)
);

AO21x2_ASAP7_75t_L g1259 ( 
.A1(n_1131),
.A2(n_1213),
.B(n_1185),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1134),
.B(n_1219),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1152),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1144),
.B(n_1160),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1179),
.A2(n_1208),
.B(n_1157),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1176),
.B(n_1147),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1216),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_1170),
.B(n_1222),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1167),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1187),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1187),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1215),
.A2(n_1154),
.B(n_1170),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1177),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1158),
.B(n_1120),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1123),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1154),
.A2(n_1188),
.B(n_1190),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1127),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1133),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1190),
.A2(n_1203),
.B(n_1198),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1156),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1137),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1212),
.B(n_1116),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1132),
.B(n_1183),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1171),
.B(n_1155),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1215),
.B(n_1221),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1172),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1181),
.B(n_1201),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1191),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1203),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1194),
.B(n_1174),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1117),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1116),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1178),
.A2(n_1193),
.B(n_1128),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1211),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1192),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1125),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1220),
.A2(n_1141),
.B(n_1189),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1172),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1228),
.Y(n_1297)
);

INVx1_ASAP7_75t_SL g1298 ( 
.A(n_1233),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1231),
.B(n_1224),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1253),
.B(n_1196),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1253),
.B(n_1115),
.Y(n_1301)
);

BUFx4_ASAP7_75t_R g1302 ( 
.A(n_1296),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1231),
.B(n_1115),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1270),
.A2(n_1128),
.B1(n_1197),
.B2(n_1153),
.Y(n_1304)
);

BUFx2_ASAP7_75t_L g1305 ( 
.A(n_1229),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1240),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1260),
.B(n_1182),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1238),
.B(n_1202),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1251),
.A2(n_1270),
.B1(n_1246),
.B2(n_1283),
.Y(n_1309)
);

AND2x4_ASAP7_75t_L g1310 ( 
.A(n_1232),
.B(n_1234),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1229),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1235),
.B(n_1128),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1242),
.B(n_1202),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1242),
.B(n_1205),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1287),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1235),
.B(n_1150),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1248),
.B(n_1230),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1261),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1261),
.B(n_1206),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1237),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1261),
.B(n_1207),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1249),
.B(n_1199),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1235),
.B(n_1252),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1254),
.B(n_1283),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1235),
.B(n_1214),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1252),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1285),
.B(n_1217),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1250),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1269),
.B(n_1165),
.Y(n_1329)
);

NOR2x1_ASAP7_75t_L g1330 ( 
.A(n_1259),
.B(n_1165),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1256),
.B(n_1214),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1255),
.B(n_1199),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1251),
.A2(n_1153),
.B1(n_1125),
.B2(n_1124),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1256),
.B(n_1257),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1309),
.A2(n_1246),
.B1(n_1244),
.B2(n_1264),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1305),
.B(n_1269),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1305),
.B(n_1268),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1324),
.B(n_1265),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1311),
.B(n_1268),
.Y(n_1339)
);

NAND4xp25_ASAP7_75t_L g1340 ( 
.A(n_1309),
.B(n_1225),
.C(n_1262),
.D(n_1243),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1317),
.B(n_1225),
.Y(n_1341)
);

OAI221xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1304),
.A2(n_1244),
.B1(n_1266),
.B2(n_1282),
.C(n_1262),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1325),
.B(n_1250),
.Y(n_1343)
);

OAI221xp5_ASAP7_75t_L g1344 ( 
.A1(n_1333),
.A2(n_1282),
.B1(n_1266),
.B2(n_1243),
.C(n_1264),
.Y(n_1344)
);

AOI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1300),
.A2(n_1267),
.B1(n_1271),
.B2(n_1241),
.C(n_1278),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1325),
.B(n_1250),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1330),
.A2(n_1274),
.B(n_1245),
.Y(n_1347)
);

NAND3xp33_ASAP7_75t_L g1348 ( 
.A(n_1330),
.B(n_1288),
.C(n_1241),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1323),
.B(n_1250),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1301),
.B(n_1271),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1322),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1307),
.B(n_1263),
.Y(n_1352)
);

NOR3xp33_ASAP7_75t_SL g1353 ( 
.A(n_1332),
.B(n_1204),
.C(n_1290),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1299),
.B(n_1263),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1299),
.B(n_1263),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1316),
.B(n_1288),
.C(n_1292),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1303),
.B(n_1239),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1303),
.B(n_1295),
.Y(n_1358)
);

OAI221xp5_ASAP7_75t_L g1359 ( 
.A1(n_1316),
.A2(n_1247),
.B1(n_1226),
.B2(n_1245),
.C(n_1289),
.Y(n_1359)
);

OAI21xp33_ASAP7_75t_L g1360 ( 
.A1(n_1312),
.A2(n_1281),
.B(n_1226),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1321),
.B(n_1257),
.Y(n_1361)
);

OAI221xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1312),
.A2(n_1289),
.B1(n_1247),
.B2(n_1226),
.C(n_1279),
.Y(n_1362)
);

NAND3xp33_ASAP7_75t_L g1363 ( 
.A(n_1329),
.B(n_1281),
.C(n_1273),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1331),
.A2(n_1259),
.B1(n_1272),
.B2(n_1276),
.C(n_1273),
.Y(n_1364)
);

OAI221xp5_ASAP7_75t_L g1365 ( 
.A1(n_1327),
.A2(n_1247),
.B1(n_1245),
.B2(n_1284),
.C(n_1236),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1302),
.A2(n_1258),
.B1(n_1286),
.B2(n_1290),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1308),
.B(n_1227),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1298),
.A2(n_1125),
.B1(n_1280),
.B2(n_1294),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1319),
.B(n_1275),
.Y(n_1369)
);

AOI221xp5_ASAP7_75t_L g1370 ( 
.A1(n_1331),
.A2(n_1259),
.B1(n_1272),
.B2(n_1276),
.C(n_1293),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1329),
.B(n_1153),
.C(n_1286),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1313),
.B(n_1227),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1337),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1337),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1343),
.B(n_1328),
.Y(n_1375)
);

AND2x2_ASAP7_75t_SL g1376 ( 
.A(n_1335),
.B(n_1328),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1352),
.B(n_1318),
.Y(n_1377)
);

OR2x2_ASAP7_75t_L g1378 ( 
.A(n_1354),
.B(n_1315),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1336),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1341),
.B(n_1355),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1364),
.B(n_1334),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1370),
.B(n_1334),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1339),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1349),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1336),
.Y(n_1385)
);

INVx3_ASAP7_75t_L g1386 ( 
.A(n_1343),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1342),
.A2(n_1274),
.B(n_1291),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1358),
.B(n_1259),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1346),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1351),
.B(n_1326),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1369),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1361),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1357),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1363),
.B(n_1326),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1363),
.B(n_1297),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1367),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1372),
.B(n_1320),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1394),
.Y(n_1398)
);

OR2x6_ASAP7_75t_SL g1399 ( 
.A(n_1388),
.B(n_1356),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1380),
.B(n_1338),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1389),
.B(n_1372),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1394),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1389),
.B(n_1356),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1395),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1395),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1379),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1388),
.A2(n_1381),
.B(n_1382),
.C(n_1387),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1379),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1380),
.B(n_1393),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1389),
.B(n_1348),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1373),
.Y(n_1411)
);

AND2x2_ASAP7_75t_SL g1412 ( 
.A(n_1376),
.B(n_1345),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1385),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1386),
.B(n_1360),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1386),
.B(n_1360),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1393),
.B(n_1350),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1386),
.B(n_1347),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1391),
.B(n_1313),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1378),
.B(n_1348),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1373),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1385),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1373),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1374),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1374),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1373),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1386),
.B(n_1347),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1386),
.B(n_1310),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1391),
.B(n_1314),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1375),
.B(n_1371),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1383),
.Y(n_1430)
);

INVxp33_ASAP7_75t_L g1431 ( 
.A(n_1397),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1390),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1411),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1403),
.B(n_1384),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1411),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1403),
.B(n_1384),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1403),
.B(n_1384),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1410),
.B(n_1396),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1410),
.B(n_1376),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1410),
.B(n_1384),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1419),
.B(n_1378),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1406),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1406),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1408),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1398),
.B(n_1378),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1414),
.B(n_1396),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1420),
.Y(n_1447)
);

AND2x2_ASAP7_75t_SL g1448 ( 
.A(n_1412),
.B(n_1376),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1420),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1408),
.Y(n_1450)
);

BUFx3_ASAP7_75t_L g1451 ( 
.A(n_1412),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1413),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1422),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1413),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1422),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1425),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1430),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1421),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1414),
.B(n_1415),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1419),
.B(n_1377),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1430),
.Y(n_1462)
);

NAND2xp67_ASAP7_75t_L g1463 ( 
.A(n_1417),
.B(n_1124),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1429),
.A2(n_1340),
.B1(n_1376),
.B2(n_1344),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1401),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1421),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1398),
.Y(n_1467)
);

AO221x1_ASAP7_75t_L g1468 ( 
.A1(n_1399),
.A2(n_1396),
.B1(n_1368),
.B2(n_1366),
.C(n_1392),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1423),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1429),
.B(n_1375),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1400),
.B(n_1306),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1423),
.Y(n_1472)
);

NAND2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1429),
.B(n_1277),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1415),
.B(n_1396),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1424),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1442),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1442),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1407),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1451),
.B(n_1432),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1439),
.B(n_1417),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1402),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1451),
.B(n_1218),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1472),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1439),
.B(n_1460),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1441),
.B(n_1402),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1443),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1443),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1439),
.B(n_1426),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1448),
.A2(n_1340),
.B1(n_1426),
.B2(n_1404),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1444),
.Y(n_1490)
);

BUFx3_ASAP7_75t_L g1491 ( 
.A(n_1465),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1460),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1465),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1444),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1450),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1471),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1450),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1470),
.B(n_1401),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1448),
.A2(n_1404),
.B1(n_1405),
.B2(n_1401),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1452),
.Y(n_1500)
);

NOR2xp33_ASAP7_75t_L g1501 ( 
.A(n_1463),
.B(n_1218),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1448),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1464),
.B(n_1409),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1427),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1452),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1464),
.B(n_1405),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1470),
.B(n_1438),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_1461),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1468),
.B(n_1399),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1468),
.B(n_1416),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1454),
.Y(n_1511)
);

NOR3xp33_ASAP7_75t_L g1512 ( 
.A(n_1478),
.B(n_1467),
.C(n_1438),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1484),
.B(n_1470),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1502),
.B(n_1463),
.Y(n_1514)
);

NOR4xp25_ASAP7_75t_SL g1515 ( 
.A(n_1503),
.B(n_1362),
.C(n_1459),
.D(n_1466),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1509),
.A2(n_1461),
.B1(n_1474),
.B2(n_1446),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1496),
.B(n_1186),
.Y(n_1517)
);

INVxp67_ASAP7_75t_L g1518 ( 
.A(n_1491),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1489),
.A2(n_1440),
.B1(n_1434),
.B2(n_1437),
.Y(n_1519)
);

NAND2xp33_ASAP7_75t_SL g1520 ( 
.A(n_1484),
.B(n_1353),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1506),
.A2(n_1445),
.B(n_1467),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1507),
.Y(n_1522)
);

NOR2x1_ASAP7_75t_L g1523 ( 
.A(n_1482),
.B(n_1454),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1496),
.B(n_1446),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1493),
.B(n_1491),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1507),
.Y(n_1526)
);

OAI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1510),
.A2(n_1382),
.B1(n_1381),
.B2(n_1387),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1492),
.B(n_1474),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1476),
.Y(n_1529)
);

OAI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1499),
.A2(n_1473),
.B1(n_1445),
.B2(n_1440),
.C(n_1437),
.Y(n_1530)
);

AOI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1492),
.A2(n_1436),
.B1(n_1434),
.B2(n_1359),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

AND2x2_ASAP7_75t_SL g1533 ( 
.A(n_1501),
.B(n_1436),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1508),
.B(n_1418),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1481),
.B(n_1428),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1480),
.B(n_1390),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1476),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1518),
.B(n_1480),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1518),
.B(n_1488),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1525),
.B(n_1488),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1532),
.B(n_1498),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1517),
.B(n_1498),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1521),
.B(n_1481),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1513),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1528),
.B(n_1504),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1485),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1529),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1522),
.B(n_1495),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1537),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1497),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1533),
.B(n_1427),
.Y(n_1554)
);

INVx1_ASAP7_75t_SL g1555 ( 
.A(n_1520),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1523),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1527),
.B(n_1511),
.Y(n_1557)
);

OAI221xp5_ASAP7_75t_L g1558 ( 
.A1(n_1544),
.A2(n_1519),
.B1(n_1530),
.B2(n_1512),
.C(n_1531),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1556),
.A2(n_1527),
.B(n_1512),
.C(n_1515),
.Y(n_1559)
);

OAI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1544),
.A2(n_1536),
.B(n_1534),
.Y(n_1560)
);

OAI21xp33_ASAP7_75t_SL g1561 ( 
.A1(n_1557),
.A2(n_1486),
.B(n_1477),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1548),
.A2(n_1490),
.B1(n_1505),
.B2(n_1500),
.C(n_1494),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_SL g1563 ( 
.A1(n_1555),
.A2(n_1542),
.B1(n_1539),
.B2(n_1538),
.Y(n_1563)
);

OAI211xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1540),
.A2(n_1490),
.B(n_1505),
.C(n_1500),
.Y(n_1564)
);

AOI21xp33_ASAP7_75t_L g1565 ( 
.A1(n_1547),
.A2(n_1535),
.B(n_1486),
.Y(n_1565)
);

AOI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1548),
.A2(n_1487),
.B(n_1477),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1543),
.B(n_1186),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1552),
.A2(n_1494),
.B1(n_1487),
.B2(n_1466),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1549),
.Y(n_1569)
);

AOI211x1_ASAP7_75t_SL g1570 ( 
.A1(n_1564),
.A2(n_1541),
.B(n_1545),
.C(n_1553),
.Y(n_1570)
);

NOR2x1_ASAP7_75t_L g1571 ( 
.A(n_1559),
.B(n_1551),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1563),
.B(n_1543),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1560),
.B(n_1547),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1566),
.B(n_1546),
.Y(n_1574)
);

XNOR2x1_ASAP7_75t_L g1575 ( 
.A(n_1569),
.B(n_1554),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1565),
.B(n_1550),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1567),
.B(n_1375),
.Y(n_1577)
);

NOR2x1_ASAP7_75t_L g1578 ( 
.A(n_1558),
.B(n_1483),
.Y(n_1578)
);

OAI322xp33_ASAP7_75t_L g1579 ( 
.A1(n_1568),
.A2(n_1483),
.A3(n_1473),
.B1(n_1459),
.B2(n_1469),
.C1(n_1475),
.C2(n_1472),
.Y(n_1579)
);

NAND4xp25_ASAP7_75t_SL g1580 ( 
.A(n_1571),
.B(n_1561),
.C(n_1562),
.D(n_1365),
.Y(n_1580)
);

AND4x1_ASAP7_75t_L g1581 ( 
.A(n_1572),
.B(n_1186),
.C(n_1195),
.D(n_1371),
.Y(n_1581)
);

INVx2_ASAP7_75t_SL g1582 ( 
.A(n_1575),
.Y(n_1582)
);

NOR2x1_ASAP7_75t_L g1583 ( 
.A(n_1573),
.B(n_1469),
.Y(n_1583)
);

NAND5xp2_ASAP7_75t_L g1584 ( 
.A(n_1574),
.B(n_1473),
.C(n_1475),
.D(n_1431),
.E(n_1195),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1576),
.Y(n_1585)
);

INVxp67_ASAP7_75t_SL g1586 ( 
.A(n_1582),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1583),
.Y(n_1587)
);

NOR2x1_ASAP7_75t_L g1588 ( 
.A(n_1585),
.B(n_1578),
.Y(n_1588)
);

NOR2x1_ASAP7_75t_L g1589 ( 
.A(n_1580),
.B(n_1579),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1581),
.A2(n_1577),
.B1(n_1570),
.B2(n_1473),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1584),
.A2(n_1435),
.B1(n_1453),
.B2(n_1462),
.Y(n_1591)
);

AOI221x1_ASAP7_75t_L g1592 ( 
.A1(n_1587),
.A2(n_1457),
.B1(n_1433),
.B2(n_1462),
.C(n_1458),
.Y(n_1592)
);

INVx1_ASAP7_75t_SL g1593 ( 
.A(n_1588),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1586),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1589),
.B(n_1195),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1590),
.A2(n_1435),
.B1(n_1453),
.B2(n_1462),
.Y(n_1596)
);

NOR3xp33_ASAP7_75t_L g1597 ( 
.A(n_1594),
.B(n_1595),
.C(n_1593),
.Y(n_1597)
);

NAND2xp33_ASAP7_75t_SL g1598 ( 
.A(n_1592),
.B(n_1204),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1596),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1597),
.Y(n_1600)
);

XOR2xp5_ASAP7_75t_L g1601 ( 
.A(n_1600),
.B(n_1599),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1601),
.A2(n_1598),
.B1(n_1591),
.B2(n_1447),
.Y(n_1602)
);

OA21x2_ASAP7_75t_L g1603 ( 
.A1(n_1601),
.A2(n_1435),
.B(n_1433),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1602),
.Y(n_1604)
);

OAI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1603),
.A2(n_1447),
.B(n_1433),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1604),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1605),
.A2(n_1447),
.B1(n_1458),
.B2(n_1457),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1606),
.A2(n_1453),
.B(n_1449),
.Y(n_1608)
);

BUFx2_ASAP7_75t_L g1609 ( 
.A(n_1608),
.Y(n_1609)
);

OAI221xp5_ASAP7_75t_R g1610 ( 
.A1(n_1609),
.A2(n_1607),
.B1(n_1455),
.B2(n_1458),
.C(n_1457),
.Y(n_1610)
);

AOI211xp5_ASAP7_75t_L g1611 ( 
.A1(n_1610),
.A2(n_1456),
.B(n_1455),
.C(n_1449),
.Y(n_1611)
);


endmodule