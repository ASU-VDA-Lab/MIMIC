module fake_jpeg_554_n_113 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_113);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_113;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_22),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_50),
.B(n_52),
.Y(n_58)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_36),
.B1(n_37),
.B2(n_31),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_40),
.B1(n_41),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_38),
.B1(n_33),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_52)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_34),
.C(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_30),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_46),
.B1(n_32),
.B2(n_4),
.Y(n_68)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_62),
.B(n_48),
.Y(n_67)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_48),
.B1(n_34),
.B2(n_53),
.Y(n_65)
);

AO21x2_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_68),
.B(n_63),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_6),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_1),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_69),
.B(n_3),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_14),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_61),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_55),
.C(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_75),
.C(n_76),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_61),
.B(n_54),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_71),
.B1(n_17),
.B2(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_80),
.Y(n_90)
);

AOI22x1_ASAP7_75t_SL g79 ( 
.A1(n_65),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_79)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_68),
.A2(n_3),
.B(n_5),
.Y(n_81)
);

OR2x2_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_6),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_20),
.B1(n_11),
.B2(n_13),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_88),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_71),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_94),
.Y(n_96)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_100),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_101),
.C(n_89),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_10),
.B1(n_15),
.B2(n_23),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_90),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_91),
.C(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_104),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_98),
.B1(n_99),
.B2(n_96),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_93),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_106),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_89),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_98),
.C(n_25),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_24),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_112),
.B(n_27),
.Y(n_113)
);


endmodule