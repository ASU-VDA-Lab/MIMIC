module fake_jpeg_15769_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_12),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_17),
.Y(n_37)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_30),
.B1(n_37),
.B2(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_20),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_36),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_65),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_70),
.Y(n_105)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_81),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_55),
.A2(n_30),
.B1(n_21),
.B2(n_19),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_76),
.A2(n_97),
.B1(n_106),
.B2(n_62),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_100),
.B1(n_103),
.B2(n_107),
.Y(n_119)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_86),
.Y(n_111)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_24),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_92),
.Y(n_117)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_43),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.C(n_16),
.Y(n_127)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_43),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_25),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_96),
.A2(n_108),
.B1(n_16),
.B2(n_22),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_19),
.B1(n_37),
.B2(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_27),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_18),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_27),
.B1(n_34),
.B2(n_23),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_45),
.B1(n_40),
.B2(n_42),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_68),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_60),
.A2(n_33),
.B1(n_40),
.B2(n_18),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_14),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_61),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_91),
.B1(n_87),
.B2(n_78),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_114),
.B(n_29),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_47),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_132),
.C(n_47),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_31),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_123),
.Y(n_156)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_131),
.Y(n_157)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_125),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_22),
.Y(n_168)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_106),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_93),
.B(n_47),
.C(n_44),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_75),
.B(n_47),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_35),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_79),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_70),
.B(n_16),
.C(n_22),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_136),
.Y(n_143)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_104),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_140),
.Y(n_151)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_142),
.B(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_119),
.A2(n_76),
.B1(n_97),
.B2(n_103),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_148),
.B1(n_150),
.B2(n_167),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_145),
.B(n_168),
.Y(n_198)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

AO22x2_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_96),
.B1(n_89),
.B2(n_109),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_163),
.B1(n_135),
.B2(n_126),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_85),
.B1(n_89),
.B2(n_61),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_108),
.B1(n_102),
.B2(n_101),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_149),
.A2(n_159),
.B1(n_169),
.B2(n_128),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_132),
.A2(n_123),
.B1(n_116),
.B2(n_129),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_153),
.B(n_174),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_126),
.B1(n_115),
.B2(n_137),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_105),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_164),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_129),
.A2(n_136),
.B1(n_121),
.B2(n_110),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_170),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_84),
.B1(n_48),
.B2(n_16),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_112),
.B(n_124),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_84),
.B1(n_44),
.B2(n_92),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_112),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_120),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_35),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_16),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_117),
.C(n_139),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_175),
.B(n_180),
.C(n_187),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_31),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_178),
.A2(n_197),
.B(n_199),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_168),
.B(n_140),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_183),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_191),
.B1(n_201),
.B2(n_206),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_161),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_195),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_156),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_147),
.A2(n_143),
.B1(n_144),
.B2(n_157),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_189),
.A2(n_163),
.B1(n_162),
.B2(n_31),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_137),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_173),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_28),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_156),
.B(n_147),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_35),
.B(n_1),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_200),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_158),
.A2(n_29),
.B1(n_18),
.B2(n_22),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_162),
.B1(n_165),
.B2(n_10),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_203),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_205),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_167),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_146),
.A2(n_128),
.B1(n_22),
.B2(n_29),
.Y(n_206)
);

O2A1O1Ixp33_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_31),
.B(n_28),
.C(n_2),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_151),
.B(n_163),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_166),
.B(n_13),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_208),
.B(n_169),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_149),
.B(n_31),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_28),
.C(n_1),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_184),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_211),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_213),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_153),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_226),
.C(n_227),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_217),
.B(n_186),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_148),
.B(n_163),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_224),
.B1(n_237),
.B2(n_238),
.Y(n_241)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_193),
.Y(n_223)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_223),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_28),
.C(n_10),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_228),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_28),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_230),
.C(n_226),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_180),
.B(n_9),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_177),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_231),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_9),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_199),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_207),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_182),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_179),
.B1(n_185),
.B2(n_189),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_249),
.B1(n_6),
.B2(n_7),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_175),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_229),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_185),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_244),
.A2(n_248),
.B(n_251),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_247),
.B(n_263),
.Y(n_268)
);

OA21x2_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_195),
.B(n_192),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_183),
.B1(n_203),
.B2(n_200),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_224),
.A2(n_176),
.B1(n_194),
.B2(n_204),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_221),
.B1(n_228),
.B2(n_237),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_190),
.B(n_176),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_194),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_256),
.C(n_260),
.Y(n_272)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_254),
.B(n_5),
.Y(n_283)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_257),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_216),
.B(n_212),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_233),
.B1(n_219),
.B2(n_222),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_235),
.A2(n_181),
.B(n_188),
.Y(n_259)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_215),
.B(n_188),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_220),
.A2(n_2),
.B(n_3),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_267),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_283),
.B(n_245),
.Y(n_297)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_274),
.A2(n_277),
.B1(n_284),
.B2(n_249),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_230),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_282),
.C(n_256),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_244),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_241),
.A2(n_218),
.B1(n_223),
.B2(n_5),
.Y(n_277)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_3),
.C(n_4),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_5),
.Y(n_280)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_281),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_5),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_239),
.B1(n_257),
.B2(n_254),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_285),
.A2(n_297),
.B1(n_248),
.B2(n_278),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_286),
.B(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_261),
.Y(n_288)
);

AND2x2_ASAP7_75t_SL g313 ( 
.A(n_288),
.B(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_261),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_242),
.C(n_272),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_264),
.A2(n_251),
.B(n_258),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_292),
.B(n_287),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_284),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_242),
.C(n_243),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_268),
.C(n_248),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_310),
.C(n_314),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_289),
.B1(n_294),
.B2(n_296),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_270),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_295),
.A2(n_267),
.B(n_282),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_293),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_272),
.C(n_275),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_315),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_290),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_290),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_262),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_298),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_285),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_6),
.C(n_7),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_318),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_323),
.C(n_324),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_297),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_286),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_294),
.B1(n_296),
.B2(n_291),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_300),
.B(n_312),
.Y(n_330)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_326),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_327),
.B(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_313),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_321),
.C(n_317),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_310),
.B1(n_314),
.B2(n_309),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_331),
.B(n_321),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_334),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_336),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_6),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);

OAI21x1_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_339),
.B(n_335),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_333),
.B(n_337),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_332),
.B(n_6),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_332),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_344),
.A2(n_7),
.B(n_338),
.Y(n_345)
);


endmodule