module fake_jpeg_224_n_167 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_167);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_38),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_2),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_47),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_55),
.Y(n_82)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_61),
.B1(n_42),
.B2(n_53),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_74),
.A2(n_75),
.B1(n_49),
.B2(n_5),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_61),
.B1(n_46),
.B2(n_50),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_54),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_64),
.B(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_47),
.B(n_44),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_66),
.B1(n_45),
.B2(n_41),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_45),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_72),
.A2(n_40),
.B1(n_50),
.B2(n_51),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_51),
.B1(n_49),
.B2(n_46),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_94),
.B1(n_9),
.B2(n_12),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_75),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_20),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_104),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_103),
.Y(n_108)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_23),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_21),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_118),
.B1(n_122),
.B2(n_117),
.Y(n_134)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_87),
.B(n_10),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_95),
.B(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_12),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_31),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_108),
.A2(n_92),
.B1(n_102),
.B2(n_13),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_132),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_92),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_107),
.C(n_118),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_27),
.B(n_37),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_19),
.B(n_28),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_26),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_136),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_24),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_143),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_116),
.C(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_147),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_146),
.A2(n_136),
.B1(n_132),
.B2(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_143),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_128),
.B(n_129),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_127),
.B1(n_135),
.B2(n_133),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_154),
.A2(n_140),
.B1(n_130),
.B2(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_142),
.B1(n_145),
.B2(n_124),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_158),
.Y(n_160)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_156),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_149),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_155),
.B(n_157),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_159),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_153),
.B(n_150),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_33),
.C(n_35),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_36),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_39),
.Y(n_167)
);


endmodule