module fake_jpeg_27565_n_308 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_308);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_308;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_33),
.B1(n_32),
.B2(n_18),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_47),
.B1(n_35),
.B2(n_40),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_45),
.B(n_53),
.Y(n_90)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_16),
.B1(n_31),
.B2(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_17),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_33),
.B1(n_20),
.B2(n_23),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_51),
.B1(n_40),
.B2(n_37),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_40),
.B1(n_37),
.B2(n_33),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g52 ( 
.A(n_34),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_54),
.B(n_31),
.Y(n_95)
);

CKINVDCx12_ASAP7_75t_R g60 ( 
.A(n_34),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_62),
.B(n_64),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_45),
.A2(n_33),
.B1(n_25),
.B2(n_24),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_74),
.B1(n_43),
.B2(n_56),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_75),
.Y(n_123)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_83),
.B1(n_51),
.B2(n_43),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_73),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_53),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_59),
.A2(n_35),
.B1(n_21),
.B2(n_22),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_34),
.C(n_38),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_21),
.B(n_22),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_76),
.B(n_95),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_79),
.B(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_91),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_82),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_23),
.B1(n_27),
.B2(n_20),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_42),
.Y(n_110)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_46),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_87),
.A2(n_93),
.B1(n_28),
.B2(n_26),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_88),
.B(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_16),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_18),
.B1(n_26),
.B2(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_16),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_42),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_21),
.B(n_18),
.C(n_19),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_49),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_112),
.B1(n_113),
.B2(n_72),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_16),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_75),
.C(n_94),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_96),
.B1(n_70),
.B2(n_82),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_91),
.B(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_56),
.B1(n_49),
.B2(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_38),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_56),
.B1(n_52),
.B2(n_36),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_61),
.B1(n_68),
.B2(n_64),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_102),
.B1(n_99),
.B2(n_101),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_80),
.B(n_38),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_42),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_127),
.A2(n_106),
.B(n_108),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_128),
.A2(n_145),
.B1(n_120),
.B2(n_114),
.Y(n_183)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_131),
.B(n_141),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_136),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_73),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_134),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_97),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_79),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_140),
.Y(n_168)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_84),
.C(n_85),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_149),
.B1(n_98),
.B2(n_107),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_65),
.C(n_34),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_138),
.B(n_65),
.C(n_30),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_101),
.A2(n_86),
.B1(n_89),
.B2(n_29),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_103),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_126),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_142),
.B(n_146),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_42),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_143),
.B(n_144),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_81),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_70),
.B(n_31),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_117),
.B(n_125),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_148),
.B(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_110),
.B1(n_125),
.B2(n_116),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_150),
.A2(n_152),
.B1(n_109),
.B2(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_78),
.Y(n_151)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_77),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_126),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_99),
.B(n_23),
.Y(n_156)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_169),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_161),
.A2(n_135),
.B(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_113),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_166),
.A2(n_170),
.B1(n_160),
.B2(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_107),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_170),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_171),
.A2(n_183),
.B1(n_137),
.B2(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_173),
.Y(n_215)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_155),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_177),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_104),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_178),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_104),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_127),
.B(n_156),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_106),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_181),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_138),
.C(n_143),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_192),
.A2(n_203),
.B(n_9),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_194),
.C(n_196),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_132),
.C(n_153),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_150),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_202),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_143),
.C(n_148),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_197),
.A2(n_213),
.B(n_182),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_199),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_163),
.B(n_152),
.Y(n_202)
);

XOR2x2_ASAP7_75t_L g203 ( 
.A(n_159),
.B(n_143),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_211),
.B1(n_157),
.B2(n_186),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_168),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_208),
.C(n_214),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_145),
.Y(n_206)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_30),
.C(n_9),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_209),
.B1(n_187),
.B2(n_184),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_128),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_20),
.B1(n_30),
.B2(n_27),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_160),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_0),
.B(n_1),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_65),
.Y(n_214)
);

A2O1A1Ixp33_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_188),
.B(n_161),
.C(n_183),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_225),
.B1(n_207),
.B2(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_206),
.A2(n_188),
.B1(n_172),
.B2(n_173),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_218),
.A2(n_222),
.B1(n_13),
.B2(n_12),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_219),
.A2(n_232),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_227),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_176),
.B1(n_162),
.B2(n_182),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_200),
.B1(n_195),
.B2(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_215),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_229),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_184),
.Y(n_229)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_189),
.Y(n_230)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_236),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_197),
.A2(n_0),
.B(n_1),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_235),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_192),
.A2(n_1),
.B(n_2),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_251),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_243),
.B1(n_252),
.B2(n_255),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_226),
.A2(n_208),
.B1(n_202),
.B2(n_209),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_194),
.C(n_193),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_253),
.C(n_233),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_213),
.B1(n_205),
.B2(n_212),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_216),
.B1(n_231),
.B2(n_222),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_214),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_250),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_212),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_15),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_221),
.B(n_228),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_14),
.C(n_13),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_254),
.B(n_239),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_216),
.B(n_255),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_219),
.B(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_261),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_224),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_265),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_267),
.B(n_270),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_269),
.Y(n_278)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_280),
.B(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_240),
.C(n_248),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_230),
.C(n_243),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_225),
.C(n_216),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_281),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_257),
.A2(n_244),
.B(n_236),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_239),
.C(n_251),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_264),
.B1(n_260),
.B2(n_256),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_290),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_291),
.B(n_3),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_256),
.B(n_13),
.Y(n_285)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

OAI211xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_12),
.B(n_11),
.C(n_10),
.Y(n_287)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_287),
.A2(n_289),
.A3(n_291),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_12),
.B1(n_10),
.B2(n_4),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_282),
.Y(n_290)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_2),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_298),
.B1(n_7),
.B2(n_5),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_278),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_273),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_277),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_3),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_295),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_301),
.A2(n_302),
.B(n_298),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_300),
.B(n_296),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_304),
.B(n_299),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_6),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_307),
.B(n_6),
.Y(n_308)
);


endmodule