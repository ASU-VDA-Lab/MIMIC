module fake_jpeg_16638_n_397 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_397);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_397;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g101 ( 
.A(n_44),
.Y(n_101)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_49),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_8),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_58),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_64),
.Y(n_97)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_8),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_7),
.Y(n_62)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx12f_ASAP7_75t_SL g69 ( 
.A(n_36),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_70),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_9),
.C(n_1),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_71),
.B(n_74),
.Y(n_85)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_36),
.B1(n_16),
.B2(n_18),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_79),
.A2(n_82),
.B1(n_88),
.B2(n_92),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_16),
.B1(n_30),
.B2(n_38),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_40),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_87),
.B(n_90),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_42),
.A2(n_30),
.B1(n_38),
.B2(n_18),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_40),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_23),
.B1(n_37),
.B2(n_28),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_91),
.A2(n_95),
.B1(n_103),
.B2(n_105),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_46),
.A2(n_23),
.B1(n_37),
.B2(n_28),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_32),
.B1(n_22),
.B2(n_21),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_94),
.A2(n_98),
.B1(n_102),
.B2(n_114),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_39),
.B1(n_24),
.B2(n_26),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_47),
.A2(n_39),
.B1(n_24),
.B2(n_26),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_100),
.B(n_73),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_44),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_44),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_51),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_106),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_52),
.A2(n_33),
.B1(n_22),
.B2(n_21),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_109),
.B1(n_120),
.B2(n_123),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_53),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_56),
.A2(n_33),
.B1(n_22),
.B2(n_21),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_48),
.A2(n_33),
.B1(n_22),
.B2(n_5),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_125),
.B1(n_76),
.B2(n_33),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_55),
.A2(n_11),
.B1(n_2),
.B2(n_5),
.Y(n_120)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_59),
.A2(n_12),
.B1(n_5),
.B2(n_6),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_65),
.A2(n_33),
.B1(n_22),
.B2(n_9),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_156),
.Y(n_187)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_136),
.A2(n_140),
.B1(n_151),
.B2(n_173),
.Y(n_199)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_6),
.B1(n_9),
.B2(n_13),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_142),
.A2(n_143),
.B1(n_166),
.B2(n_159),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_14),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_144),
.B(n_146),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_130),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_183),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_83),
.B(n_49),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_148),
.B(n_159),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_0),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_150),
.B(n_170),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_61),
.B1(n_45),
.B2(n_0),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_153),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_104),
.Y(n_157)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_0),
.B1(n_123),
.B2(n_105),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_122),
.B1(n_148),
.B2(n_145),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_0),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_94),
.A2(n_0),
.B(n_85),
.Y(n_160)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_160),
.B(n_172),
.C(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_78),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_168),
.Y(n_195)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_164),
.A2(n_122),
.B1(n_127),
.B2(n_174),
.Y(n_186)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_165),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_118),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_102),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_175),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_93),
.B(n_89),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_93),
.B(n_131),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_180),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_109),
.A2(n_117),
.B1(n_107),
.B2(n_112),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_80),
.Y(n_174)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_178),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_77),
.A2(n_106),
.B1(n_82),
.B2(n_119),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_177),
.A2(n_164),
.B1(n_139),
.B2(n_178),
.Y(n_224)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_81),
.B(n_115),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_81),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_119),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_186),
.A2(n_188),
.B1(n_191),
.B2(n_197),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_159),
.A2(n_154),
.B1(n_141),
.B2(n_163),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_193),
.B(n_203),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_201),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_148),
.B1(n_176),
.B2(n_159),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_198),
.B(n_223),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_149),
.Y(n_203)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_166),
.B(n_160),
.C(n_170),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_204),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_150),
.C(n_162),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_208),
.B(n_215),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g210 ( 
.A(n_144),
.B(n_134),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_210),
.B(n_218),
.C(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_143),
.B(n_155),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_213),
.B(n_221),
.Y(n_238)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_152),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_135),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_133),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_143),
.B(n_180),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_218),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_155),
.B(n_165),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_224),
.A2(n_153),
.B1(n_199),
.B2(n_222),
.Y(n_237)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_138),
.Y(n_225)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_137),
.Y(n_227)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_191),
.A2(n_139),
.B1(n_181),
.B2(n_182),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_232),
.A2(n_236),
.B1(n_237),
.B2(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_234),
.Y(n_271)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_235),
.B(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_198),
.A2(n_153),
.B1(n_223),
.B2(n_197),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_239),
.B(n_246),
.C(n_251),
.Y(n_291)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_194),
.Y(n_240)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_240),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_184),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_187),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_255),
.Y(n_288)
);

MAJx2_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_204),
.C(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_248),
.Y(n_276)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_249),
.Y(n_295)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_263),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_222),
.A2(n_195),
.B1(n_210),
.B2(n_193),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_205),
.B1(n_219),
.B2(n_211),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_253),
.A2(n_261),
.B1(n_265),
.B2(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_207),
.A2(n_196),
.B(n_230),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_264),
.B(n_270),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_206),
.A2(n_190),
.B1(n_230),
.B2(n_212),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_206),
.B(n_229),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_207),
.A2(n_217),
.B(n_216),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_217),
.A2(n_185),
.B1(n_203),
.B2(n_192),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_215),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_269),
.Y(n_292)
);

INVxp33_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_189),
.B(n_209),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_209),
.B(n_227),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_256),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_185),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_265),
.C(n_245),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g274 ( 
.A1(n_238),
.A2(n_200),
.A3(n_226),
.B1(n_228),
.B2(n_246),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_274),
.B(n_291),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_259),
.A2(n_200),
.B(n_228),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_279),
.A2(n_284),
.B(n_286),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_281),
.A2(n_282),
.B(n_289),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_253),
.B(n_252),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_259),
.A2(n_241),
.B(n_238),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_244),
.A2(n_236),
.B1(n_237),
.B2(n_232),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_290),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_258),
.B(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_261),
.B(n_269),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_293),
.A2(n_299),
.B1(n_271),
.B2(n_277),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_239),
.A2(n_266),
.B(n_240),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_231),
.B(n_284),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_277),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_234),
.A2(n_242),
.B1(n_254),
.B2(n_250),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_303),
.B(n_311),
.C(n_317),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_235),
.B1(n_249),
.B2(n_233),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_304),
.A2(n_309),
.B1(n_300),
.B2(n_298),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_262),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_325),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_282),
.A2(n_233),
.B1(n_257),
.B2(n_231),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_308),
.A2(n_314),
.B1(n_320),
.B2(n_323),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_286),
.A2(n_231),
.B1(n_283),
.B2(n_289),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_310),
.A2(n_324),
.B(n_296),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_273),
.C(n_280),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_278),
.Y(n_312)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_312),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_279),
.A2(n_290),
.B1(n_283),
.B2(n_287),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_294),
.B(n_274),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_280),
.B(n_281),
.C(n_293),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_302),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_318),
.Y(n_335)
);

AO21x2_ASAP7_75t_L g320 ( 
.A1(n_299),
.A2(n_301),
.B(n_272),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_288),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_292),
.B(n_288),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_328),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_272),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_295),
.Y(n_325)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_327),
.A2(n_320),
.B1(n_324),
.B2(n_307),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_276),
.B(n_297),
.C(n_295),
.Y(n_328)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_330),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_311),
.B(n_296),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_321),
.C(n_322),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_335),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_314),
.A2(n_300),
.B1(n_298),
.B2(n_275),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_337),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_341),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_320),
.A2(n_275),
.B1(n_324),
.B2(n_313),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_304),
.B1(n_313),
.B2(n_323),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_343),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_320),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_328),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_331),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_317),
.A2(n_309),
.B1(n_303),
.B2(n_305),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_346),
.A2(n_319),
.B1(n_318),
.B2(n_312),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_305),
.B(n_308),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_347),
.B(n_340),
.Y(n_358)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_339),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_348),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_335),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_351),
.B(n_334),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_356),
.C(n_358),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_357),
.A2(n_364),
.B1(n_353),
.B2(n_350),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_333),
.C(n_331),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_363),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_361),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_347),
.B(n_329),
.CI(n_346),
.CON(n_362),
.SN(n_362)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_362),
.B(n_352),
.CI(n_360),
.CON(n_371),
.SN(n_371)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_336),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_341),
.A2(n_344),
.B1(n_330),
.B2(n_338),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_367),
.A2(n_369),
.B(n_375),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_353),
.A2(n_348),
.B1(n_333),
.B2(n_329),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_368),
.A2(n_372),
.B1(n_357),
.B2(n_358),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_370),
.B(n_364),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_368),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_355),
.B1(n_359),
.B2(n_356),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_355),
.B(n_359),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_381),
.C(n_382),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_377),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_349),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_378),
.B(n_380),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_374),
.A2(n_362),
.B(n_354),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_373),
.B(n_362),
.C(n_354),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_379),
.A2(n_367),
.B1(n_372),
.B2(n_369),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_379),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_387),
.A2(n_383),
.B1(n_386),
.B2(n_375),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_366),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_389),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_382),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_391),
.A2(n_390),
.B(n_366),
.Y(n_392)
);

OAI311xp33_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_375),
.A3(n_391),
.B1(n_377),
.C1(n_384),
.Y(n_393)
);

NAND4xp25_ASAP7_75t_SL g394 ( 
.A(n_393),
.B(n_370),
.C(n_381),
.D(n_373),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_394),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_389),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_371),
.B(n_374),
.Y(n_397)
);


endmodule