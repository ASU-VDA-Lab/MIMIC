module fake_jpeg_19120_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_8),
.B(n_38),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_3),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

BUFx8_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_0),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_86),
.B(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_65),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_55),
.B(n_66),
.C(n_77),
.Y(n_101)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_92),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_49),
.B(n_64),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_100),
.Y(n_120)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_93),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_51),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_59),
.Y(n_129)
);

OA22x2_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_76),
.B1(n_73),
.B2(n_58),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_117),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_115),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_108),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_57),
.B1(n_74),
.B2(n_60),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_53),
.B1(n_69),
.B2(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_70),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_124),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_82),
.B1(n_50),
.B2(n_48),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_101),
.B(n_71),
.Y(n_122)
);

AOI32xp33_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_2),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_61),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_120),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_132),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_72),
.B(n_29),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_128),
.A2(n_32),
.B(n_10),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_133),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_135),
.Y(n_141)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_71),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_113),
.A2(n_69),
.B(n_62),
.C(n_68),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_140),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_114),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_39),
.B(n_17),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_126),
.B1(n_125),
.B2(n_117),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_147),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_148),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_146),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_139),
.Y(n_151)
);

OAI21x1_ASAP7_75t_L g152 ( 
.A1(n_151),
.A2(n_143),
.B(n_144),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_126),
.B(n_134),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_31),
.A3(n_21),
.B1(n_23),
.B2(n_24),
.C1(n_26),
.C2(n_27),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_110),
.B(n_40),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_41),
.Y(n_159)
);


endmodule