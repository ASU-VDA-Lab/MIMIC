module fake_netlist_1_12755_n_702 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_702);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_702;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_72), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_55), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_35), .Y(n_106) );
INVx2_ASAP7_75t_SL g107 ( .A(n_42), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_29), .B(n_53), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_70), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_65), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_12), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_83), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_89), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_20), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_40), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
BUFx10_ASAP7_75t_L g118 ( .A(n_30), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_26), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_34), .Y(n_121) );
BUFx10_ASAP7_75t_L g122 ( .A(n_33), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_36), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_103), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_84), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_100), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_78), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_17), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_18), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_7), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_15), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_91), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_92), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g136 ( .A(n_38), .Y(n_136) );
INVxp33_ASAP7_75t_L g137 ( .A(n_4), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_97), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_37), .Y(n_139) );
INVxp67_ASAP7_75t_L g140 ( .A(n_52), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_82), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_7), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_81), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_27), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_22), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_32), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_137), .B(n_0), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_105), .Y(n_149) );
NOR2x1_ASAP7_75t_L g150 ( .A(n_106), .B(n_0), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_107), .B(n_1), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_128), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_112), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_131), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_107), .B(n_2), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_128), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_146), .Y(n_160) );
OA21x2_ASAP7_75t_L g161 ( .A1(n_116), .A2(n_5), .B(n_6), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_117), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_120), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_131), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_118), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_126), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_154), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_149), .B(n_127), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_149), .B(n_133), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_160), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_152), .A2(n_119), .B1(n_146), .B2(n_136), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_154), .Y(n_178) );
INVx4_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_151), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_161), .Y(n_181) );
OR2x2_ASAP7_75t_L g182 ( .A(n_148), .B(n_115), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_155), .B(n_118), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
AND2x2_ASAP7_75t_SL g185 ( .A(n_161), .B(n_134), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_154), .Y(n_187) );
INVx3_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_155), .B(n_165), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_153), .B(n_145), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_154), .Y(n_191) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_168), .B(n_104), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_179), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_186), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_183), .B(n_155), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_183), .B(n_179), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_182), .A2(n_148), .B1(n_165), .B2(n_155), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_168), .Y(n_198) );
AO22x1_ASAP7_75t_L g199 ( .A1(n_168), .A2(n_150), .B1(n_148), .B2(n_157), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_172), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_183), .B(n_155), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_189), .B(n_165), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_189), .Y(n_205) );
AND2x6_ASAP7_75t_SL g206 ( .A(n_177), .B(n_157), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_189), .B(n_165), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_171), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_179), .B(n_165), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_182), .B(n_153), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_182), .A2(n_124), .B1(n_109), .B2(n_144), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_171), .Y(n_212) );
INVx1_ASAP7_75t_SL g213 ( .A(n_186), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_179), .A2(n_166), .B1(n_163), .B2(n_161), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_179), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_176), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_176), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_186), .B(n_163), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_180), .B(n_166), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_180), .B(n_174), .Y(n_221) );
NAND3xp33_ASAP7_75t_L g222 ( .A(n_174), .B(n_152), .C(n_159), .Y(n_222) );
OAI22xp33_ASAP7_75t_L g223 ( .A1(n_177), .A2(n_159), .B1(n_114), .B2(n_111), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_218), .A2(n_188), .B(n_181), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_213), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_219), .B(n_170), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_218), .A2(n_188), .B(n_181), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_210), .A2(n_185), .B(n_188), .C(n_181), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_197), .B(n_170), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_205), .B(n_173), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_204), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_199), .B(n_173), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_207), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_194), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_196), .A2(n_188), .B(n_181), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_209), .A2(n_188), .B(n_181), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_198), .B(n_190), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_221), .B(n_190), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_195), .B(n_185), .Y(n_240) );
AO32x1_ASAP7_75t_L g241 ( .A1(n_208), .A2(n_164), .A3(n_158), .B1(n_156), .B2(n_184), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_199), .B(n_185), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_203), .A2(n_200), .B(n_198), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_220), .B(n_185), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_200), .A2(n_187), .B(n_175), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_201), .B(n_187), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_192), .B(n_150), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_211), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_201), .A2(n_141), .B1(n_125), .B2(n_135), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_222), .B(n_130), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_202), .B(n_187), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_202), .A2(n_184), .B(n_178), .Y(n_253) );
AOI221xp5_ASAP7_75t_SL g254 ( .A1(n_232), .A2(n_239), .B1(n_223), .B2(n_248), .C(n_226), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_239), .A2(n_208), .B(n_217), .C(n_212), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_230), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_225), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_235), .B(n_206), .Y(n_258) );
NAND3xp33_ASAP7_75t_SL g259 ( .A(n_249), .B(n_104), .C(n_147), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_228), .A2(n_217), .B(n_192), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_250), .Y(n_261) );
NAND2xp33_ASAP7_75t_L g262 ( .A(n_245), .B(n_214), .Y(n_262) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_251), .A2(n_142), .B1(n_132), .B2(n_131), .C(n_140), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_224), .A2(n_169), .B(n_184), .Y(n_264) );
INVxp67_ASAP7_75t_L g265 ( .A(n_230), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_243), .A2(n_156), .B(n_158), .C(n_164), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_236), .A2(n_215), .B(n_216), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_238), .B(n_215), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_238), .Y(n_269) );
AOI221x1_ASAP7_75t_L g270 ( .A1(n_242), .A2(n_154), .B1(n_162), .B2(n_167), .C(n_191), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_227), .A2(n_216), .B(n_175), .Y(n_271) );
AO31x2_ASAP7_75t_L g272 ( .A1(n_240), .A2(n_169), .A3(n_184), .B(n_178), .Y(n_272) );
BUFx10_ASAP7_75t_L g273 ( .A(n_238), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_237), .A2(n_178), .B(n_175), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_231), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_229), .B(n_139), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_253), .A2(n_178), .B(n_175), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_275), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_256), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_240), .B1(n_234), .B2(n_233), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_270), .A2(n_246), .B(n_169), .Y(n_281) );
INVx2_ASAP7_75t_SL g282 ( .A(n_273), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_254), .A2(n_244), .B1(n_233), .B2(n_161), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_273), .B(n_244), .Y(n_284) );
CKINVDCx11_ASAP7_75t_R g285 ( .A(n_257), .Y(n_285) );
OA21x2_ASAP7_75t_L g286 ( .A1(n_255), .A2(n_252), .B(n_247), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_273), .Y(n_287) );
INVx6_ASAP7_75t_L g288 ( .A(n_269), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_258), .B(n_252), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_277), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_261), .Y(n_291) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_268), .B(n_247), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_265), .B(n_125), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_259), .B(n_161), .Y(n_294) );
BUFx6f_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
CKINVDCx11_ASAP7_75t_R g296 ( .A(n_263), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_272), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_264), .A2(n_169), .B(n_241), .Y(n_298) );
AND2x4_ASAP7_75t_SL g299 ( .A(n_284), .B(n_122), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_280), .B(n_260), .Y(n_300) );
AO21x2_ASAP7_75t_L g301 ( .A1(n_290), .A2(n_266), .B(n_264), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_296), .A2(n_262), .B1(n_276), .B2(n_131), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_290), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_297), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_295), .Y(n_306) );
INVx5_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_297), .Y(n_308) );
AOI21xp5_ASAP7_75t_SL g309 ( .A1(n_280), .A2(n_266), .B(n_143), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_295), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
AO21x1_ASAP7_75t_SL g312 ( .A1(n_287), .A2(n_283), .B(n_278), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_279), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_286), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_286), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_295), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_284), .B(n_272), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_281), .A2(n_274), .B(n_271), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_295), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_286), .Y(n_324) );
INVx5_ASAP7_75t_L g325 ( .A(n_307), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_310), .Y(n_327) );
OR2x6_ASAP7_75t_L g328 ( .A(n_309), .B(n_282), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g329 ( .A(n_299), .B(n_285), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_320), .B(n_286), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_311), .B(n_272), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_305), .B(n_272), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_308), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_308), .B(n_281), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_320), .B(n_286), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_320), .B(n_282), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_311), .B(n_283), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_302), .Y(n_339) );
NOR2xp33_ASAP7_75t_R g340 ( .A(n_307), .B(n_291), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_313), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_313), .Y(n_342) );
OR2x2_ASAP7_75t_L g343 ( .A(n_314), .B(n_287), .Y(n_343) );
NAND2x1_ASAP7_75t_L g344 ( .A(n_302), .B(n_298), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_304), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_317), .B(n_298), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_303), .A2(n_294), .B1(n_288), .B2(n_292), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_323), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_317), .B(n_298), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_303), .A2(n_289), .B1(n_288), .B2(n_262), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_318), .B(n_281), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_314), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_318), .B(n_298), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_323), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_324), .B(n_323), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_310), .Y(n_358) );
NAND2x1p5_ASAP7_75t_SL g359 ( .A(n_306), .B(n_158), .Y(n_359) );
INVx3_ASAP7_75t_L g360 ( .A(n_319), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_292), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_316), .B(n_292), .Y(n_362) );
AOI222xp33_ASAP7_75t_L g363 ( .A1(n_299), .A2(n_288), .B1(n_293), .B2(n_122), .C1(n_129), .C2(n_135), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_300), .B(n_294), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_319), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_306), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_326), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_337), .B(n_306), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_326), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_346), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_337), .B(n_335), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_335), .B(n_315), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_346), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_325), .B(n_307), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_325), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_333), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_358), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_335), .B(n_315), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_330), .B(n_315), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_341), .B(n_300), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_330), .B(n_322), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_357), .B(n_322), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_341), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_357), .B(n_322), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_338), .B(n_312), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_342), .B(n_301), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_348), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_332), .B(n_301), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_350), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_325), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_334), .B(n_319), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_338), .B(n_312), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_354), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_354), .B(n_301), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_331), .B(n_301), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_361), .B(n_319), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_361), .B(n_319), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_356), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_347), .B(n_319), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_325), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_336), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_332), .Y(n_408) );
AND2x4_ASAP7_75t_L g409 ( .A(n_334), .B(n_319), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_348), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_347), .B(n_321), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_347), .B(n_321), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_331), .Y(n_413) );
INVxp67_ASAP7_75t_L g414 ( .A(n_358), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_336), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_351), .B(n_355), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_336), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_339), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_339), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_351), .B(n_321), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_351), .B(n_321), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_355), .B(n_321), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_362), .B(n_307), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_339), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_345), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_345), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_362), .B(n_307), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_364), .B(n_299), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_362), .B(n_307), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_366), .B(n_307), .Y(n_430) );
NAND4xp25_ASAP7_75t_L g431 ( .A(n_363), .B(n_129), .C(n_108), .D(n_156), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_364), .B(n_288), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_368), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_408), .B(n_343), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_374), .B(n_334), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_368), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_395), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_395), .B(n_329), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_370), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_373), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_408), .B(n_343), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_372), .B(n_327), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_370), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_375), .Y(n_445) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_431), .A2(n_363), .B(n_349), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_379), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_373), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_372), .B(n_327), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_413), .B(n_366), .Y(n_450) );
NAND2x1p5_ASAP7_75t_L g451 ( .A(n_395), .B(n_325), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_416), .B(n_345), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_373), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_413), .B(n_334), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_379), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_416), .B(n_367), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_386), .B(n_352), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_382), .B(n_367), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_371), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_386), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_382), .B(n_367), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_423), .B(n_325), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_374), .B(n_353), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_395), .B(n_325), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_381), .B(n_353), .Y(n_465) );
NAND2x1_ASAP7_75t_L g466 ( .A(n_378), .B(n_328), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_381), .B(n_353), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_388), .B(n_349), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_384), .B(n_353), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_406), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_377), .B(n_340), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_384), .B(n_344), .Y(n_472) );
AND2x4_ASAP7_75t_L g473 ( .A(n_406), .B(n_360), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_369), .B(n_344), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_388), .B(n_328), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_369), .B(n_328), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_420), .B(n_360), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_398), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_420), .B(n_360), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_420), .B(n_411), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_423), .B(n_360), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_398), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_411), .B(n_328), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_380), .B(n_328), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_380), .B(n_328), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_400), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_400), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_431), .B(n_6), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_412), .B(n_365), .Y(n_489) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_406), .B(n_365), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_404), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_387), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_412), .B(n_365), .Y(n_493) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_371), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_421), .B(n_365), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_421), .B(n_359), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_422), .B(n_359), .Y(n_497) );
NOR2xp33_ASAP7_75t_SL g498 ( .A(n_377), .B(n_288), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_404), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g500 ( .A(n_378), .B(n_428), .C(n_390), .D(n_397), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_387), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_414), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_405), .B(n_158), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_387), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_414), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_422), .B(n_359), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_405), .B(n_164), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_385), .B(n_8), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_385), .B(n_8), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_385), .B(n_9), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_410), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_410), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_394), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_511), .B(n_383), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_502), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g516 ( .A1(n_446), .A2(n_428), .B1(n_432), .B2(n_397), .C1(n_390), .C2(n_383), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_505), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_512), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_480), .B(n_376), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_480), .B(n_376), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_433), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_469), .B(n_427), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_503), .B(n_392), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_469), .B(n_427), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_442), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_488), .A2(n_378), .B1(n_432), .B2(n_429), .Y(n_526) );
INVx2_ASAP7_75t_SL g527 ( .A(n_438), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_466), .A2(n_392), .B(n_393), .C(n_401), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_449), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_436), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_463), .B(n_429), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_470), .Y(n_532) );
OR4x1_ASAP7_75t_L g533 ( .A(n_437), .B(n_417), .C(n_425), .D(n_424), .Y(n_533) );
INVxp67_ASAP7_75t_SL g534 ( .A(n_459), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_439), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_452), .B(n_456), .Y(n_536) );
NOR2xp67_ASAP7_75t_SL g537 ( .A(n_500), .B(n_430), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_443), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_503), .B(n_389), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_507), .B(n_389), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_463), .B(n_402), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_507), .B(n_393), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_464), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_458), .B(n_405), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_434), .B(n_401), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_441), .B(n_391), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_465), .B(n_402), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_444), .Y(n_548) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_464), .B(n_430), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_461), .B(n_391), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_459), .B(n_399), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_445), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_447), .Y(n_553) );
AOI32xp33_ASAP7_75t_L g554 ( .A1(n_488), .A2(n_403), .A3(n_409), .B1(n_396), .B2(n_418), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_495), .B(n_399), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_494), .Y(n_556) );
OR2x6_ASAP7_75t_L g557 ( .A(n_451), .B(n_394), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_465), .B(n_403), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_457), .B(n_417), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_455), .Y(n_560) );
AOI31xp33_ASAP7_75t_L g561 ( .A1(n_451), .A2(n_418), .A3(n_425), .B(n_424), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_464), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_467), .B(n_396), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_460), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_478), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_482), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_SL g567 ( .A1(n_437), .A2(n_494), .B(n_510), .C(n_509), .Y(n_567) );
NOR2xp67_ASAP7_75t_SL g568 ( .A(n_471), .B(n_394), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_474), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_486), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_450), .B(n_426), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_487), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_454), .B(n_407), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_473), .B(n_396), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_468), .B(n_426), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_467), .B(n_396), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_491), .B(n_407), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_499), .B(n_407), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_477), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_477), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_479), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_462), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_490), .B(n_415), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_483), .B(n_415), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_479), .Y(n_585) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_508), .B(n_415), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_471), .A2(n_409), .B1(n_419), .B2(n_426), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_435), .B(n_409), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_519), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_516), .A2(n_472), .B1(n_493), .B2(n_489), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_536), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_549), .A2(n_476), .B1(n_484), .B2(n_485), .Y(n_592) );
OAI22xp33_ASAP7_75t_SL g593 ( .A1(n_527), .A2(n_498), .B1(n_475), .B2(n_473), .Y(n_593) );
A2O1A1Ixp33_ASAP7_75t_L g594 ( .A1(n_537), .A2(n_472), .B(n_435), .C(n_473), .Y(n_594) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_554), .A2(n_489), .B1(n_493), .B2(n_506), .C(n_497), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_532), .B(n_496), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_532), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_516), .A2(n_481), .B1(n_409), .B2(n_501), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_559), .B(n_513), .Y(n_599) );
OAI21xp5_ASAP7_75t_L g600 ( .A1(n_561), .A2(n_513), .B(n_504), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_533), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_545), .B(n_440), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_561), .B(n_440), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_528), .A2(n_504), .B(n_501), .Y(n_604) );
AOI211x1_ASAP7_75t_L g605 ( .A1(n_568), .A2(n_9), .B(n_10), .C(n_11), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_567), .A2(n_164), .B1(n_453), .B2(n_448), .C(n_492), .Y(n_606) );
OAI21xp5_ASAP7_75t_L g607 ( .A1(n_586), .A2(n_492), .B(n_453), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_587), .B(n_448), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_520), .Y(n_609) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_526), .A2(n_10), .B(n_11), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_518), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_546), .B(n_419), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_534), .A2(n_419), .B(n_138), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_526), .A2(n_162), .B1(n_122), .B2(n_138), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g615 ( .A1(n_543), .A2(n_141), .B1(n_147), .B2(n_143), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_557), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_543), .A2(n_162), .B1(n_110), .B2(n_123), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_557), .A2(n_162), .B1(n_113), .B2(n_121), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_515), .Y(n_619) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_562), .A2(n_162), .B1(n_191), .B2(n_167), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g621 ( .A1(n_557), .A2(n_241), .B(n_162), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_517), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_525), .B(n_12), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_562), .A2(n_162), .B1(n_14), .B2(n_15), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_521), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_563), .B(n_162), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_551), .B(n_267), .C(n_14), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_576), .B(n_13), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_514), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_556), .A2(n_167), .B1(n_191), .B2(n_17), .C(n_18), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_551), .A2(n_167), .B1(n_191), .B2(n_19), .C(n_20), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_529), .B(n_13), .Y(n_632) );
AO22x2_ASAP7_75t_L g633 ( .A1(n_569), .A2(n_16), .B1(n_21), .B2(n_23), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_587), .A2(n_16), .B1(n_21), .B2(n_23), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g636 ( .A1(n_582), .A2(n_24), .B1(n_25), .B2(n_191), .Y(n_636) );
OR2x2_ASAP7_75t_L g637 ( .A(n_555), .B(n_24), .Y(n_637) );
AOI21xp5_ASAP7_75t_SL g638 ( .A1(n_600), .A2(n_574), .B(n_523), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_616), .B(n_588), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_590), .A2(n_574), .B1(n_581), .B2(n_580), .Y(n_640) );
AOI322xp5_ASAP7_75t_L g641 ( .A1(n_595), .A2(n_585), .A3(n_579), .B1(n_531), .B2(n_522), .C1(n_524), .C2(n_558), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_611), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_600), .B(n_530), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_629), .B(n_514), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_603), .A2(n_571), .B(n_575), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_598), .A2(n_566), .B1(n_535), .B2(n_538), .C(n_548), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_609), .B(n_552), .Y(n_647) );
AOI222xp33_ASAP7_75t_L g648 ( .A1(n_601), .A2(n_560), .B1(n_553), .B2(n_564), .C1(n_572), .C2(n_570), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_591), .B(n_565), .Y(n_649) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_594), .A2(n_542), .B(n_578), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_593), .A2(n_584), .B1(n_550), .B2(n_573), .C(n_539), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_592), .A2(n_540), .B1(n_547), .B2(n_541), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_597), .A2(n_544), .B1(n_577), .B2(n_25), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_596), .A2(n_191), .B1(n_167), .B2(n_241), .Y(n_654) );
AOI21xp33_ASAP7_75t_SL g655 ( .A1(n_633), .A2(n_28), .B(n_31), .Y(n_655) );
AOI221x1_ASAP7_75t_L g656 ( .A1(n_633), .A2(n_191), .B1(n_167), .B2(n_241), .C(n_44), .Y(n_656) );
XOR2x2_ASAP7_75t_L g657 ( .A(n_605), .B(n_39), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_597), .A2(n_191), .B1(n_167), .B2(n_45), .C(n_46), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_626), .A2(n_167), .B(n_43), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_606), .A2(n_41), .B(n_47), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_589), .B(n_48), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_619), .B(n_49), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_622), .B(n_50), .Y(n_663) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_627), .A2(n_51), .B(n_54), .C(n_56), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g665 ( .A1(n_635), .A2(n_57), .B(n_58), .Y(n_665) );
OAI211xp5_ASAP7_75t_L g666 ( .A1(n_610), .A2(n_59), .B(n_60), .C(n_61), .Y(n_666) );
AO21x1_ASAP7_75t_L g667 ( .A1(n_637), .A2(n_62), .B(n_63), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_634), .A2(n_64), .B1(n_66), .B2(n_67), .C(n_68), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_602), .A2(n_69), .B(n_71), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_625), .Y(n_670) );
NAND3xp33_ASAP7_75t_SL g671 ( .A(n_636), .B(n_73), .C(n_75), .Y(n_671) );
AOI211x1_ASAP7_75t_L g672 ( .A1(n_632), .A2(n_76), .B(n_77), .C(n_79), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_623), .A2(n_80), .B1(n_86), .B2(n_87), .Y(n_673) );
AO221x1_ASAP7_75t_L g674 ( .A1(n_618), .A2(n_88), .B1(n_90), .B2(n_93), .C(n_94), .Y(n_674) );
OAI22xp33_ASAP7_75t_L g675 ( .A1(n_604), .A2(n_96), .B1(n_99), .B2(n_101), .Y(n_675) );
NAND3xp33_ASAP7_75t_SL g676 ( .A(n_613), .B(n_102), .C(n_614), .Y(n_676) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_608), .A2(n_624), .B1(n_628), .B2(n_630), .C(n_599), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_631), .B(n_617), .C(n_615), .D(n_620), .Y(n_678) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_657), .B(n_653), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_641), .A2(n_677), .B(n_638), .C(n_648), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_655), .B(n_667), .C(n_664), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_648), .B(n_645), .Y(n_682) );
OAI211xp5_ASAP7_75t_SL g683 ( .A1(n_643), .A2(n_651), .B(n_640), .C(n_646), .Y(n_683) );
INVxp33_ASAP7_75t_L g684 ( .A(n_678), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_676), .B(n_671), .C(n_675), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_684), .B(n_650), .Y(n_686) );
AND5x1_ASAP7_75t_L g687 ( .A(n_685), .B(n_662), .C(n_668), .D(n_673), .E(n_652), .Y(n_687) );
NAND2x1p5_ASAP7_75t_L g688 ( .A(n_682), .B(n_660), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g689 ( .A(n_680), .B(n_666), .C(n_658), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_686), .B(n_679), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_689), .A2(n_683), .B1(n_681), .B2(n_674), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_688), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_691), .B(n_642), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_692), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g695 ( .A1(n_694), .A2(n_690), .B1(n_687), .B2(n_649), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_693), .A2(n_661), .B1(n_670), .B2(n_644), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_695), .A2(n_647), .B1(n_665), .B2(n_639), .Y(n_697) );
AOI21xp33_ASAP7_75t_SL g698 ( .A1(n_696), .A2(n_663), .B(n_669), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_697), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_698), .B(n_659), .Y(n_700) );
AO221x2_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_607), .B1(n_672), .B2(n_612), .C(n_656), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_607), .B1(n_654), .B2(n_621), .Y(n_702) );
endmodule