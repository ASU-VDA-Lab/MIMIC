module fake_jpeg_32039_n_530 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_530);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g143 ( 
.A(n_52),
.Y(n_143)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_60),
.B(n_61),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_10),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_49),
.B(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_62),
.B(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_29),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_64),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_48),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_9),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_22),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_83),
.Y(n_141)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_27),
.B(n_11),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_84),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_27),
.B(n_11),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_88),
.B(n_91),
.Y(n_151)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_30),
.B(n_11),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_8),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_96),
.B(n_97),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_35),
.Y(n_131)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_99),
.B(n_100),
.Y(n_155)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_35),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_24),
.B(n_28),
.C(n_23),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_106),
.B(n_156),
.Y(n_170)
);

HAxp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_50),
.CON(n_108),
.SN(n_108)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_108),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_50),
.B1(n_37),
.B2(n_24),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_112),
.A2(n_132),
.B1(n_154),
.B2(n_54),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_56),
.A2(n_47),
.B1(n_44),
.B2(n_31),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_115),
.A2(n_127),
.B1(n_159),
.B2(n_75),
.Y(n_179)
);

NAND3xp33_ASAP7_75t_L g121 ( 
.A(n_67),
.B(n_47),
.C(n_44),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_124),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_52),
.B(n_41),
.Y(n_124)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_41),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_126),
.B(n_131),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_19),
.B1(n_26),
.B2(n_40),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_31),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_148),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_96),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_161),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_59),
.A2(n_43),
.B1(n_38),
.B2(n_28),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_52),
.B(n_40),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_57),
.A2(n_26),
.B1(n_19),
.B2(n_36),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_157),
.A2(n_162),
.B1(n_138),
.B2(n_51),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_85),
.A2(n_36),
.B1(n_20),
.B2(n_35),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_79),
.B(n_36),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_63),
.A2(n_36),
.B1(n_20),
.B2(n_35),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_167),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_168),
.Y(n_269)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_139),
.A2(n_65),
.B1(n_68),
.B2(n_71),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_173),
.A2(n_186),
.B1(n_218),
.B2(n_223),
.Y(n_248)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_174),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_95),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_175),
.B(n_185),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_176),
.B(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_134),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_177),
.Y(n_266)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_178),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_104),
.B(n_81),
.C(n_92),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_180),
.B(n_184),
.Y(n_252)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_181),
.Y(n_240)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_190),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_101),
.B(n_86),
.C(n_35),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_84),
.B1(n_87),
.B2(n_101),
.Y(n_186)
);

AO22x1_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_90),
.B1(n_82),
.B2(n_77),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_187),
.B(n_191),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_120),
.A2(n_66),
.B1(n_36),
.B2(n_20),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_199),
.B1(n_207),
.B2(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_36),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_192),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_144),
.A2(n_20),
.B1(n_1),
.B2(n_0),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_193),
.A2(n_198),
.B1(n_136),
.B2(n_113),
.Y(n_241)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_194),
.Y(n_274)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_196),
.Y(n_239)
);

INVx11_ASAP7_75t_L g197 ( 
.A(n_102),
.Y(n_197)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_109),
.A2(n_20),
.B1(n_12),
.B2(n_2),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_141),
.A2(n_12),
.B1(n_17),
.B2(n_3),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_105),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_160),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_209),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_108),
.A2(n_12),
.B1(n_17),
.B2(n_4),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_13),
.B(n_14),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_128),
.A2(n_13),
.B1(n_16),
.B2(n_5),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_122),
.Y(n_208)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_143),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_210),
.B(n_211),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_143),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_217),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_106),
.B(n_8),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_213),
.B(n_222),
.Y(n_267)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_151),
.A2(n_8),
.B1(n_15),
.B2(n_5),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_18),
.B1(n_6),
.B2(n_13),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_163),
.B1(n_146),
.B2(n_116),
.Y(n_245)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_129),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_122),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_103),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_221),
.Y(n_264)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_103),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_6),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_110),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_213),
.A2(n_116),
.B(n_158),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_224),
.A2(n_256),
.B(n_210),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_187),
.A2(n_146),
.B1(n_147),
.B2(n_163),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_231),
.A2(n_270),
.B1(n_259),
.B2(n_249),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_170),
.B(n_114),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_233),
.B(n_234),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_164),
.B(n_114),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_188),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_263),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_243),
.B1(n_245),
.B2(n_255),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_137),
.B1(n_152),
.B2(n_147),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_176),
.A2(n_107),
.B1(n_102),
.B2(n_110),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_251),
.A2(n_253),
.B1(n_260),
.B2(n_271),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_166),
.A2(n_107),
.B1(n_113),
.B2(n_140),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_191),
.A2(n_140),
.B1(n_136),
.B2(n_1),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_193),
.A2(n_14),
.B1(n_18),
.B2(n_0),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_200),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_222),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_273),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_187),
.A2(n_0),
.B1(n_18),
.B2(n_193),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_182),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_169),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_211),
.Y(n_273)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_193),
.B1(n_197),
.B2(n_208),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_277),
.A2(n_285),
.B1(n_300),
.B2(n_317),
.Y(n_331)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

OAI21xp33_ASAP7_75t_SL g279 ( 
.A1(n_256),
.A2(n_175),
.B(n_185),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_279),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_244),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_280),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_290),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_246),
.B1(n_271),
.B2(n_252),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_282),
.A2(n_284),
.B1(n_301),
.B2(n_304),
.Y(n_324)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_246),
.A2(n_205),
.B1(n_206),
.B2(n_171),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_216),
.B1(n_212),
.B2(n_196),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_287),
.Y(n_342)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_254),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_288),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_229),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_291),
.Y(n_357)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_292),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_252),
.B(n_180),
.C(n_221),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_293),
.B(n_318),
.C(n_300),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_229),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_294),
.B(n_298),
.Y(n_330)
);

XOR2x2_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_219),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_297),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_296),
.B(n_307),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_178),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_226),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_252),
.A2(n_218),
.B1(n_168),
.B2(n_165),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_247),
.A2(n_201),
.B1(n_192),
.B2(n_194),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_237),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_306),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_195),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_303),
.B(n_296),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_247),
.A2(n_174),
.B1(n_181),
.B2(n_204),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_241),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_315),
.B(n_270),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_248),
.A2(n_209),
.B1(n_214),
.B2(n_273),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_309),
.A2(n_313),
.B1(n_269),
.B2(n_232),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_264),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_310),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_224),
.A2(n_233),
.B(n_225),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_240),
.B(n_235),
.Y(n_333)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_235),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_314),
.Y(n_329)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_238),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_255),
.A2(n_251),
.B(n_224),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_234),
.A2(n_272),
.B(n_236),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_316),
.A2(n_228),
.B(n_230),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_243),
.A2(n_245),
.B1(n_225),
.B2(n_236),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_253),
.B(n_240),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_250),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_319),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_321),
.A2(n_230),
.B1(n_232),
.B2(n_269),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_305),
.A2(n_249),
.B1(n_266),
.B2(n_250),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_332),
.A2(n_333),
.B(n_341),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_305),
.A2(n_258),
.B1(n_266),
.B2(n_242),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_336),
.B(n_351),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_282),
.A2(n_258),
.B1(n_242),
.B2(n_232),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_339),
.A2(n_359),
.B1(n_275),
.B2(n_310),
.Y(n_373)
);

AO22x1_ASAP7_75t_L g340 ( 
.A1(n_315),
.A2(n_268),
.B1(n_262),
.B2(n_274),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_340),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_311),
.A2(n_262),
.B(n_274),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_343),
.A2(n_346),
.B1(n_340),
.B2(n_344),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_289),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_345),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_346),
.A2(n_299),
.B1(n_301),
.B2(n_298),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_297),
.B(n_269),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_350),
.C(n_355),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_303),
.B(n_293),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_280),
.A2(n_281),
.B(n_308),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_318),
.B(n_304),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_341),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_295),
.B(n_314),
.C(n_283),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_288),
.C(n_290),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_319),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_358),
.B(n_362),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_299),
.A2(n_275),
.B1(n_317),
.B2(n_285),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_278),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_320),
.B(n_294),
.Y(n_362)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_329),
.Y(n_365)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_329),
.Y(n_366)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_330),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_367),
.B(n_385),
.Y(n_420)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_330),
.Y(n_368)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_353),
.Y(n_371)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_371),
.Y(n_419)
);

AOI322xp5_ASAP7_75t_L g372 ( 
.A1(n_351),
.A2(n_335),
.A3(n_323),
.B1(n_345),
.B2(n_327),
.C1(n_340),
.C2(n_326),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_SL g411 ( 
.A(n_372),
.B(n_348),
.C(n_325),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_382),
.B1(n_397),
.B2(n_352),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_350),
.B(n_307),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_393),
.C(n_349),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_376),
.A2(n_380),
.B1(n_387),
.B2(n_392),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_378),
.B(n_379),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_331),
.A2(n_291),
.B1(n_312),
.B2(n_286),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_381),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_313),
.B1(n_287),
.B2(n_292),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_383),
.A2(n_334),
.B(n_352),
.Y(n_407)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_342),
.Y(n_384)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_326),
.Y(n_385)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_386),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_331),
.A2(n_276),
.B1(n_306),
.B2(n_354),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_388),
.A2(n_357),
.B(n_343),
.Y(n_422)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_389),
.Y(n_403)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_344),
.Y(n_390)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_390),
.Y(n_410)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_332),
.A2(n_340),
.B1(n_327),
.B2(n_324),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_355),
.C(n_347),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_322),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_394),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_324),
.A2(n_356),
.B1(n_333),
.B2(n_339),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_408),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_328),
.Y(n_404)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_405),
.A2(n_409),
.B1(n_411),
.B2(n_424),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_407),
.A2(n_374),
.B1(n_369),
.B2(n_364),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_347),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_373),
.A2(n_328),
.B1(n_361),
.B2(n_322),
.Y(n_409)
);

XOR2x2_ASAP7_75t_SL g413 ( 
.A(n_388),
.B(n_348),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_415),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_336),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_338),
.B(n_358),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_418),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_357),
.C(n_338),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_375),
.C(n_379),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_422),
.B(n_425),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_337),
.Y(n_423)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_423),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_374),
.A2(n_369),
.B1(n_397),
.B2(n_395),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_395),
.B(n_337),
.C(n_360),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_365),
.B(n_366),
.Y(n_427)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_427),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_431),
.C(n_432),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_378),
.C(n_363),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_400),
.B(n_396),
.C(n_392),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_415),
.C(n_414),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_433),
.B(n_434),
.C(n_452),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_409),
.C(n_411),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_399),
.B(n_371),
.Y(n_435)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_435),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g460 ( 
.A1(n_436),
.A2(n_407),
.B(n_422),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_412),
.A2(n_364),
.B1(n_382),
.B2(n_383),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_451),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_424),
.B(n_387),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_398),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_380),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_442),
.B(n_443),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_404),
.B(n_381),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_384),
.Y(n_444)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_444),
.Y(n_457)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_446),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_401),
.B(n_386),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_450),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_418),
.B(n_389),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_412),
.A2(n_376),
.B1(n_391),
.B2(n_390),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_423),
.C(n_402),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_419),
.B(n_426),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_453),
.B(n_398),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_SL g459 ( 
.A(n_447),
.B(n_413),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_L g483 ( 
.A(n_459),
.B(n_462),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_465),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_442),
.A2(n_441),
.B1(n_439),
.B2(n_445),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_460),
.B1(n_438),
.B2(n_459),
.Y(n_488)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_463),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_428),
.B(n_403),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_430),
.Y(n_466)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_SL g468 ( 
.A(n_437),
.B(n_403),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_469),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_428),
.B(n_416),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_416),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_470),
.B(n_436),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_474),
.Y(n_477)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_440),
.Y(n_473)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_473),
.Y(n_486)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_478),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_429),
.C(n_433),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_482),
.C(n_458),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_481),
.B(n_489),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_471),
.C(n_465),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_448),
.Y(n_485)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_471),
.B(n_467),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_490),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_488),
.A2(n_481),
.B1(n_476),
.B2(n_464),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_454),
.A2(n_448),
.B(n_434),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_456),
.B(n_431),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_462),
.A2(n_437),
.B1(n_451),
.B2(n_406),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_491),
.B(n_464),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_475),
.B(n_461),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_494),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_480),
.B(n_469),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_497),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_485),
.A2(n_454),
.B(n_468),
.Y(n_499)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_499),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_501),
.B(n_482),
.C(n_476),
.Y(n_509)
);

INVx11_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_502),
.Y(n_510)
);

OR2x2_ASAP7_75t_SL g503 ( 
.A(n_489),
.B(n_406),
.Y(n_503)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_503),
.Y(n_512)
);

XNOR2x1_ASAP7_75t_SL g504 ( 
.A(n_483),
.B(n_491),
.Y(n_504)
);

NOR2xp67_ASAP7_75t_SL g507 ( 
.A(n_504),
.B(n_483),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_498),
.A2(n_500),
.B1(n_486),
.B2(n_494),
.Y(n_505)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_505),
.Y(n_515)
);

AO21x1_ASAP7_75t_L g516 ( 
.A1(n_507),
.A2(n_504),
.B(n_503),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_509),
.B(n_513),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_477),
.C(n_479),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_511),
.A2(n_496),
.B(n_499),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_514),
.A2(n_518),
.B(n_519),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_508),
.Y(n_523)
);

OAI211xp5_ASAP7_75t_L g518 ( 
.A1(n_512),
.A2(n_484),
.B(n_500),
.C(n_492),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g519 ( 
.A1(n_506),
.A2(n_410),
.B(n_502),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_510),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_521),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_515),
.B(n_509),
.C(n_513),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_522),
.Y(n_525)
);

XNOR2x1_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_518),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_526),
.A2(n_520),
.B(n_524),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_527),
.B(n_523),
.C(n_505),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_410),
.Y(n_529)
);

NAND2x1_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_479),
.Y(n_530)
);


endmodule