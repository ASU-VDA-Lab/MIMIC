module fake_jpeg_14373_n_574 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_574);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_574;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx3_ASAP7_75t_SL g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_20),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_62),
.B(n_80),
.Y(n_127)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_69),
.Y(n_161)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_0),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_22),
.B(n_0),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_82),
.B(n_99),
.Y(n_167)
);

BUFx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_85),
.Y(n_172)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_89),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_91),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g117 ( 
.A(n_92),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_103),
.Y(n_114)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_101),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_102),
.B(n_49),
.Y(n_158)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_49),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_106),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_35),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_48),
.B(n_0),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_22),
.B(n_1),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_26),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_83),
.A2(n_35),
.B1(n_48),
.B2(n_21),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_111),
.A2(n_116),
.B1(n_132),
.B2(n_140),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_61),
.A2(n_35),
.B1(n_48),
.B2(n_21),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_51),
.C(n_46),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_119),
.B(n_46),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_125),
.B(n_153),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_57),
.A2(n_35),
.B1(n_45),
.B2(n_43),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_158),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_92),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_62),
.A2(n_44),
.B1(n_42),
.B2(n_45),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_150),
.B1(n_24),
.B2(n_27),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_50),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_145),
.B(n_47),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_88),
.A2(n_44),
.B1(n_42),
.B2(n_34),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_146),
.A2(n_156),
.B1(n_49),
.B2(n_76),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_82),
.A2(n_38),
.B1(n_50),
.B2(n_26),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_38),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_32),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_157),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_105),
.A2(n_34),
.B1(n_49),
.B2(n_27),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_32),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_101),
.A2(n_47),
.B1(n_39),
.B2(n_51),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_168),
.A2(n_49),
.B1(n_72),
.B2(n_68),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_53),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_77),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_87),
.B1(n_85),
.B2(n_84),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_173),
.A2(n_196),
.B1(n_225),
.B2(n_146),
.Y(n_253)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_162),
.Y(n_174)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_175),
.Y(n_240)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_114),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_177),
.B(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_178),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_134),
.Y(n_180)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_181),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_113),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_183),
.B(n_214),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_184),
.B(n_218),
.Y(n_245)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_131),
.Y(n_186)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_188),
.A2(n_202),
.B1(n_228),
.B2(n_232),
.Y(n_238)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_189),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_190),
.B(n_203),
.Y(n_260)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

INVx11_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_192),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_39),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_201),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_194),
.Y(n_283)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_195),
.Y(n_279)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_126),
.Y(n_197)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_115),
.Y(n_198)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_198),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_142),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_200),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_24),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_127),
.A2(n_34),
.B1(n_49),
.B2(n_69),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_205),
.B(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_207),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_208),
.A2(n_224),
.B1(n_130),
.B2(n_113),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_112),
.Y(n_210)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_210),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_120),
.A2(n_71),
.A3(n_67),
.B1(n_66),
.B2(n_49),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_132),
.B(n_156),
.Y(n_255)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_212),
.Y(n_287)
);

INVx13_ASAP7_75t_L g213 ( 
.A(n_136),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_135),
.Y(n_215)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_217),
.B(n_222),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_159),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_147),
.B(n_163),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_129),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_220),
.B(n_229),
.Y(n_266)
);

INVx3_ASAP7_75t_SL g221 ( 
.A(n_163),
.Y(n_221)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_223),
.B(n_233),
.Y(n_286)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_116),
.A2(n_34),
.B1(n_36),
.B2(n_4),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_169),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_129),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_121),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_227),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_109),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_130),
.B(n_4),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_133),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_231),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_109),
.Y(n_232)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_133),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_234),
.B(n_235),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_154),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_190),
.B(n_124),
.C(n_111),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_244),
.B(n_262),
.C(n_223),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_251),
.A2(n_261),
.B1(n_269),
.B2(n_175),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_253),
.B(n_255),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_196),
.A2(n_140),
.B1(n_149),
.B2(n_152),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_256),
.A2(n_280),
.B1(n_183),
.B2(n_184),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_199),
.A2(n_201),
.B1(n_221),
.B2(n_222),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_182),
.A2(n_164),
.B1(n_154),
.B2(n_160),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_182),
.B(n_152),
.C(n_122),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_208),
.A2(n_128),
.B1(n_160),
.B2(n_164),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_264),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_182),
.B(n_161),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_277),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_211),
.A2(n_161),
.B1(n_110),
.B2(n_7),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_206),
.B(n_110),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_179),
.B(n_5),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_278),
.B(n_210),
.Y(n_309)
);

OA22x2_ASAP7_75t_L g281 ( 
.A1(n_227),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g308 ( 
.A(n_281),
.B(n_8),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_252),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_297),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_191),
.B(n_176),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_290),
.A2(n_294),
.B(n_279),
.Y(n_347)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_237),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_248),
.B(n_187),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_293),
.B(n_323),
.Y(n_341)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_252),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_296),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_250),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_308),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_181),
.B1(n_185),
.B2(n_197),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_299),
.A2(n_311),
.B1(n_317),
.B2(n_328),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_248),
.B(n_219),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_313),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_305),
.B1(n_314),
.B2(n_315),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_238),
.A2(n_251),
.B1(n_244),
.B2(n_268),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_306),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_260),
.A2(n_193),
.B(n_216),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_319),
.B(n_306),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g358 ( 
.A(n_309),
.B(n_325),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_267),
.Y(n_310)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_310),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_277),
.A2(n_262),
.B1(n_280),
.B2(n_245),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_326),
.C(n_242),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_243),
.B(n_246),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_261),
.A2(n_204),
.B1(n_186),
.B2(n_189),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_266),
.A2(n_174),
.B1(n_214),
.B2(n_192),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_246),
.B(n_198),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_324),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_276),
.A2(n_230),
.B1(n_226),
.B2(n_228),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_281),
.A2(n_232),
.B1(n_233),
.B2(n_231),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_318),
.A2(n_285),
.B1(n_267),
.B2(n_275),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_241),
.A2(n_209),
.B(n_213),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_288),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_322),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_236),
.A2(n_212),
.B1(n_195),
.B2(n_10),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g355 ( 
.A(n_321),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_288),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_270),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_288),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_270),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_8),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_272),
.Y(n_327)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_327),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_236),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_329),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_281),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_330),
.A2(n_281),
.B1(n_274),
.B2(n_242),
.Y(n_353)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_284),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_274),
.B(n_11),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_275),
.B(n_17),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_336),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_249),
.B(n_12),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g375 ( 
.A(n_335),
.Y(n_375)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_303),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_339),
.B(n_370),
.C(n_371),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_340),
.A2(n_366),
.B1(n_367),
.B2(n_310),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_347),
.A2(n_310),
.B(n_332),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_290),
.A2(n_273),
.B(n_274),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_348),
.A2(n_376),
.B(n_378),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_353),
.A2(n_359),
.B1(n_373),
.B2(n_294),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_298),
.A2(n_265),
.B1(n_240),
.B2(n_247),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_360),
.B(n_372),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_315),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_364),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_334),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_300),
.A2(n_285),
.B1(n_239),
.B2(n_249),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_305),
.A2(n_265),
.B1(n_258),
.B2(n_254),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_293),
.B(n_302),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_313),
.B(n_284),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_291),
.C(n_316),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_291),
.A2(n_247),
.B1(n_273),
.B2(n_258),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_295),
.A2(n_291),
.B(n_311),
.Y(n_376)
);

OAI32xp33_ASAP7_75t_L g377 ( 
.A1(n_308),
.A2(n_279),
.A3(n_239),
.B1(n_263),
.B2(n_271),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_377),
.B(n_331),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_307),
.B(n_254),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_263),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_317),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_380),
.B(n_314),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_339),
.B(n_326),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_395),
.C(n_416),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_383),
.A2(n_392),
.B1(n_404),
.B2(n_415),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_338),
.A2(n_304),
.B1(n_297),
.B2(n_330),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_388),
.B1(n_390),
.B2(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_385),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_348),
.A2(n_376),
.B(n_378),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_397),
.B(n_413),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_338),
.A2(n_299),
.B1(n_308),
.B2(n_318),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_354),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_389),
.B(n_399),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_367),
.A2(n_308),
.B1(n_296),
.B2(n_292),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_346),
.Y(n_391)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_391),
.Y(n_432)
);

AOI32xp33_ASAP7_75t_L g392 ( 
.A1(n_341),
.A2(n_319),
.A3(n_289),
.B1(n_324),
.B2(n_322),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_365),
.Y(n_393)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_309),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_347),
.A2(n_333),
.B(n_320),
.Y(n_397)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_398),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_356),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_400),
.A2(n_408),
.B(n_407),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_352),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_401),
.B(n_410),
.Y(n_435)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_405),
.Y(n_420)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_407),
.Y(n_426)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_343),
.A2(n_327),
.B(n_336),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_409),
.B(n_379),
.Y(n_424)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_362),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_411),
.Y(n_429)
);

O2A1O1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_343),
.A2(n_335),
.B(n_328),
.C(n_287),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_358),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_414),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_351),
.A2(n_301),
.B1(n_329),
.B2(n_282),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_344),
.B(n_271),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_372),
.A2(n_301),
.B1(n_287),
.B2(n_282),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_417),
.A2(n_363),
.B1(n_349),
.B2(n_374),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_404),
.A2(n_361),
.B1(n_344),
.B2(n_380),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_418),
.B(n_422),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_386),
.B(n_360),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_421),
.B(n_427),
.C(n_430),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_396),
.A2(n_340),
.B1(n_343),
.B2(n_350),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_433),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_386),
.B(n_371),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_350),
.C(n_373),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g431 ( 
.A(n_385),
.B(n_375),
.C(n_365),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_416),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_412),
.B(n_351),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_395),
.B(n_362),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_437),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_383),
.A2(n_394),
.B1(n_381),
.B2(n_387),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_443),
.Y(n_461)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_441),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_381),
.A2(n_400),
.B(n_397),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_442),
.A2(n_355),
.B(n_393),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_402),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_405),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_445),
.B(n_393),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_446),
.A2(n_413),
.B(n_406),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_349),
.B1(n_353),
.B2(n_359),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_384),
.A2(n_345),
.B1(n_363),
.B2(n_377),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_382),
.B(n_369),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_450),
.B(n_12),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_452),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_446),
.A2(n_408),
.B(n_410),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_453),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_423),
.A2(n_444),
.B1(n_436),
.B2(n_439),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_454),
.A2(n_458),
.B1(n_428),
.B2(n_422),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g457 ( 
.A1(n_442),
.A2(n_436),
.B(n_438),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_423),
.A2(n_388),
.B1(n_390),
.B2(n_417),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_435),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_464),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_462),
.B(n_425),
.Y(n_493)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_435),
.Y(n_463)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_463),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_SL g464 ( 
.A1(n_444),
.A2(n_391),
.B(n_409),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_369),
.Y(n_465)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_465),
.Y(n_482)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_420),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_466),
.B(n_469),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_467),
.A2(n_477),
.B(n_434),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_420),
.Y(n_469)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_346),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_475),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_426),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_474),
.A2(n_476),
.B1(n_479),
.B2(n_429),
.Y(n_490)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

INVx13_ASAP7_75t_L g477 ( 
.A(n_432),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_440),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_421),
.C(n_433),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_485),
.B(n_503),
.C(n_492),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_427),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_487),
.B(n_495),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_490),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_491),
.A2(n_498),
.B1(n_456),
.B2(n_455),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_460),
.B(n_419),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_492),
.B(n_497),
.Y(n_518)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_493),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_494),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_478),
.B(n_430),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_439),
.B1(n_418),
.B2(n_443),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_496),
.A2(n_499),
.B1(n_500),
.B2(n_501),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_460),
.B(n_419),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_458),
.A2(n_434),
.B1(n_445),
.B2(n_424),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_471),
.A2(n_450),
.B1(n_437),
.B2(n_16),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_461),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_461),
.A2(n_15),
.B1(n_16),
.B2(n_455),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_460),
.B(n_457),
.C(n_468),
.Y(n_503)
);

INVx11_ASAP7_75t_L g504 ( 
.A(n_481),
.Y(n_504)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_489),
.A2(n_457),
.B(n_451),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_507),
.A2(n_465),
.B(n_472),
.Y(n_538)
);

MAJx2_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_462),
.C(n_454),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_510),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_512),
.B(n_499),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_495),
.B(n_456),
.C(n_452),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_520),
.C(n_488),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_484),
.B(n_463),
.Y(n_515)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_515),
.Y(n_534)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_516),
.Y(n_536)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_502),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_522),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_497),
.B(n_464),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_519),
.B(n_498),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_467),
.C(n_476),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_482),
.B(n_459),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g526 ( 
.A(n_521),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_480),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_SL g523 ( 
.A(n_507),
.B(n_486),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_523),
.B(n_533),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_524),
.B(n_525),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_487),
.C(n_488),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_506),
.B(n_479),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_527),
.B(n_531),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_513),
.A2(n_491),
.B1(n_466),
.B2(n_469),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_528),
.B(n_535),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_520),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_489),
.C(n_474),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_483),
.C(n_470),
.Y(n_535)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_537),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_547),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_543),
.B(n_525),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_536),
.A2(n_505),
.B1(n_521),
.B2(n_508),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_545),
.A2(n_546),
.B1(n_501),
.B2(n_523),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_526),
.A2(n_505),
.B1(n_515),
.B2(n_514),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_L g547 ( 
.A1(n_534),
.A2(n_504),
.B1(n_509),
.B2(n_512),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_532),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_548),
.B(n_549),
.Y(n_552)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_531),
.Y(n_549)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_541),
.A2(n_535),
.B(n_529),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_551),
.B(n_555),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_554),
.B(n_558),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_539),
.A2(n_524),
.B(n_529),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_544),
.B(n_518),
.C(n_530),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_557),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_543),
.B(n_533),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_556),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_560),
.B(n_550),
.Y(n_566)
);

NOR2x1_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_545),
.Y(n_561)
);

NAND4xp25_ASAP7_75t_L g564 ( 
.A(n_561),
.B(n_540),
.C(n_552),
.D(n_546),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_566),
.Y(n_567)
);

AOI21xp33_ASAP7_75t_L g565 ( 
.A1(n_562),
.A2(n_540),
.B(n_558),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_565),
.B(n_559),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_563),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_569),
.B(n_567),
.C(n_550),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_561),
.B(n_453),
.Y(n_571)
);

OAI321xp33_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_477),
.A3(n_522),
.B1(n_475),
.B2(n_500),
.C(n_518),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_483),
.C(n_477),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_573),
.B(n_519),
.Y(n_574)
);


endmodule