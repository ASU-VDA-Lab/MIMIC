module fake_ibex_307_n_1455 (n_151, n_147, n_85, n_167, n_128, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_8, n_118, n_224, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_27, n_165, n_242, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_14, n_0, n_239, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_80, n_172, n_215, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_92, n_144, n_170, n_213, n_101, n_190, n_113, n_138, n_230, n_96, n_185, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_132, n_174, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1455);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_8;
input n_118;
input n_224;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_242;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_80;
input n_172;
input n_215;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_213;
input n_101;
input n_190;
input n_113;
input n_138;
input n_230;
input n_96;
input n_185;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_132;
input n_174;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1455;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_1382;
wire n_273;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_280;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_279;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1412;
wire n_262;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1301;
wire n_257;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_1434;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_639;
wire n_1332;
wire n_482;
wire n_282;
wire n_1424;
wire n_870;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_252;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_256;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1152;
wire n_371;
wire n_1036;
wire n_974;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_258;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1452;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1364;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_267;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_1420;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_272;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_268;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_303;
wire n_717;
wire n_1357;
wire n_668;
wire n_871;
wire n_266;
wire n_1339;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_260;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_281;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_255;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_317;
wire n_326;
wire n_270;
wire n_1340;
wire n_259;
wire n_276;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_251;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_278;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1188;
wire n_261;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_490;
wire n_407;
wire n_595;
wire n_1001;
wire n_269;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_246;
wire n_922;
wire n_851;
wire n_993;
wire n_253;
wire n_300;
wire n_1135;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_1337;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_1406;
wire n_804;
wire n_484;
wire n_480;
wire n_354;
wire n_1057;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_248;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_277;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_247;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1221;
wire n_284;
wire n_1047;
wire n_1374;
wire n_1435;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1257;
wire n_274;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1362;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_1330;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_249;
wire n_1443;
wire n_478;
wire n_336;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1187;
wire n_1361;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_265;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1369;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1381;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1419;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_263;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_305;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_264;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_254;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_271;
wire n_1393;
wire n_984;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g246 ( 
.A(n_78),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_235),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_54),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_94),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_101),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_214),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_76),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_30),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_181),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_144),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_131),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_103),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_34),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_224),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_191),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_158),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_195),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_139),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_219),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_170),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_190),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_178),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_187),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_65),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_188),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_133),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_59),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_155),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_55),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_154),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_236),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_40),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_48),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_171),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_57),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_243),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_152),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_98),
.Y(n_289)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_143),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_223),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_228),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_194),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

BUFx2_ASAP7_75t_SL g298 ( 
.A(n_160),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_46),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_212),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_28),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_162),
.Y(n_302)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_126),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_11),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_25),
.Y(n_305)
);

NOR2xp67_ASAP7_75t_L g306 ( 
.A(n_95),
.B(n_172),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_230),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_113),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_76),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_38),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_117),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_65),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_186),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_17),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_132),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_161),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_34),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_83),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_179),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_53),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_30),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_112),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_180),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_88),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_89),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_106),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_0),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_101),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_67),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_64),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_98),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_220),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_15),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_107),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_196),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_111),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_164),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_33),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_35),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_3),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_198),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_100),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_226),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_83),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_244),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_169),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_189),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_231),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_221),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_176),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_128),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_233),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_15),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_46),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_205),
.Y(n_356)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_211),
.B(n_67),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_234),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_163),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_33),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_206),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_108),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_23),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_237),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_22),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_66),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_185),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_177),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_36),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_102),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_134),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_26),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_96),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_63),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_99),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_203),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_215),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_51),
.Y(n_378)
);

BUFx10_ASAP7_75t_L g379 ( 
.A(n_209),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_42),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_202),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_217),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_142),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_225),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_122),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_140),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_149),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_110),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_165),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_201),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_166),
.Y(n_391)
);

CKINVDCx6p67_ASAP7_75t_R g392 ( 
.A(n_104),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_135),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_112),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_138),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_174),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_218),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_240),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_222),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_22),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_153),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_199),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_216),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_200),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_110),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_17),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_204),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_52),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_85),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_68),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_192),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_238),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_82),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_102),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_1),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_49),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_141),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_232),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_93),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_90),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_81),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_167),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_118),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_106),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_91),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_184),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_114),
.Y(n_427)
);

BUFx10_ASAP7_75t_L g428 ( 
.A(n_119),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_207),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_159),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_197),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_157),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_87),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_61),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_148),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_173),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_70),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_229),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_156),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_150),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_182),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_74),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_175),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_81),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_213),
.Y(n_445)
);

BUFx8_ASAP7_75t_SL g446 ( 
.A(n_254),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_253),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_303),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_248),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_285),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_440),
.B(n_1),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_305),
.Y(n_452)
);

AND2x6_ASAP7_75t_L g453 ( 
.A(n_303),
.B(n_115),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_372),
.B(n_2),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_408),
.B(n_290),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g456 ( 
.A(n_303),
.B(n_116),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_253),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_247),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_247),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_290),
.B(n_2),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

OAI22x1_ASAP7_75t_SL g463 ( 
.A1(n_254),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_253),
.Y(n_464)
);

BUFx12f_ASAP7_75t_L g465 ( 
.A(n_316),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_378),
.B(n_4),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_361),
.B(n_5),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_316),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_426),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_416),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_265),
.A2(n_121),
.B(n_120),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_426),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_265),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_273),
.A2(n_124),
.B(n_123),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_302),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_270),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_273),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_272),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_425),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_270),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_327),
.B(n_6),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_314),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_437),
.B(n_6),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_275),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_314),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_272),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_333),
.Y(n_490)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_316),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_277),
.B(n_7),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_439),
.B(n_7),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_277),
.B(n_315),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_333),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_325),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_345),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_340),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_340),
.B(n_8),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_379),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_281),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_281),
.Y(n_503)
);

BUFx8_ASAP7_75t_SL g504 ( 
.A(n_331),
.Y(n_504)
);

BUFx12f_ASAP7_75t_L g505 ( 
.A(n_379),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_389),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_439),
.B(n_8),
.Y(n_507)
);

INVx2_ASAP7_75t_SL g508 ( 
.A(n_398),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_345),
.B(n_9),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_389),
.B(n_10),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_392),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_511)
);

OA21x2_ASAP7_75t_L g512 ( 
.A1(n_390),
.A2(n_127),
.B(n_125),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_390),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_402),
.Y(n_515)
);

INVx4_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

BUFx8_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_432),
.B(n_12),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_331),
.B(n_13),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_288),
.B(n_14),
.Y(n_522)
);

INVx5_ASAP7_75t_L g523 ( 
.A(n_428),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_420),
.B(n_14),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_432),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_435),
.A2(n_130),
.B(n_129),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_435),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_497),
.B(n_516),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_506),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_506),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_492),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_506),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_506),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_525),
.Y(n_534)
);

INVx8_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_513),
.B(n_246),
.Y(n_536)
);

AO22x2_ASAP7_75t_L g537 ( 
.A1(n_520),
.A2(n_255),
.B1(n_260),
.B2(n_251),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_525),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_449),
.B(n_261),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_525),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_492),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_492),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_497),
.B(n_516),
.Y(n_543)
);

AND3x2_ASAP7_75t_L g544 ( 
.A(n_484),
.B(n_489),
.C(n_481),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_500),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_478),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_525),
.Y(n_547)
);

BUFx10_ASAP7_75t_L g548 ( 
.A(n_499),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_479),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_500),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_479),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_499),
.Y(n_553)
);

BUFx16f_ASAP7_75t_R g554 ( 
.A(n_449),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_479),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_453),
.B(n_256),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_479),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

AO21x2_ASAP7_75t_L g560 ( 
.A1(n_477),
.A2(n_268),
.B(n_267),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_510),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_518),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_518),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_513),
.B(n_269),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_485),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_466),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_447),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_485),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_485),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_517),
.B(n_427),
.C(n_424),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_448),
.B(n_274),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_495),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_522),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_513),
.B(n_276),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_466),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_448),
.B(n_278),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_519),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_495),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_478),
.Y(n_581)
);

INVx8_ASAP7_75t_L g582 ( 
.A(n_501),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_448),
.B(n_486),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_447),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_SL g586 ( 
.A(n_522),
.B(n_261),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_448),
.B(n_486),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_447),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_453),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_461),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_501),
.Y(n_591)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_446),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_461),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_501),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_468),
.B(n_294),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_446),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_461),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_471),
.Y(n_599)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_508),
.B(n_297),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_448),
.B(n_311),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_521),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_457),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_471),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_482),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_482),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_453),
.B(n_256),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_452),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_465),
.B(n_344),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_521),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_453),
.B(n_257),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_514),
.Y(n_615)
);

AND2x6_ASAP7_75t_L g616 ( 
.A(n_451),
.B(n_313),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_454),
.A2(n_511),
.B1(n_524),
.B2(n_509),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_456),
.B(n_451),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_L g619 ( 
.A(n_456),
.B(n_257),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_521),
.B(n_280),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_521),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_523),
.B(n_346),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_456),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_464),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_472),
.Y(n_625)
);

CKINVDCx6p67_ASAP7_75t_R g626 ( 
.A(n_465),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_464),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_523),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_494),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_494),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_491),
.B(n_322),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_460),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_469),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_470),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_493),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_523),
.B(n_350),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_450),
.B(n_351),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_459),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_470),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_475),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_475),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_517),
.B(n_353),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_480),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_480),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_470),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_L g647 ( 
.A(n_456),
.B(n_258),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_470),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_470),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_474),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_487),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_502),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_474),
.Y(n_653)
);

INVx5_ASAP7_75t_L g654 ( 
.A(n_456),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_491),
.B(n_359),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_474),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_503),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_528),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g659 ( 
.A(n_579),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_462),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_543),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_635),
.B(n_462),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_600),
.B(n_462),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_589),
.B(n_505),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_600),
.B(n_574),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_539),
.Y(n_668)
);

BUFx12f_ASAP7_75t_SL g669 ( 
.A(n_631),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_611),
.B(n_456),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_554),
.Y(n_672)
);

NAND2x1p5_ASAP7_75t_L g673 ( 
.A(n_643),
.B(n_507),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_SL g674 ( 
.A(n_589),
.B(n_282),
.Y(n_674)
);

BUFx6f_ASAP7_75t_SL g675 ( 
.A(n_536),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_629),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_654),
.B(n_262),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_626),
.B(n_322),
.Y(n_678)
);

NOR2xp67_ASAP7_75t_L g679 ( 
.A(n_592),
.B(n_467),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_R g680 ( 
.A(n_546),
.B(n_282),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_567),
.B(n_483),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_630),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_586),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_654),
.B(n_263),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_576),
.B(n_488),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_590),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_594),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_598),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_654),
.B(n_263),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_599),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_536),
.B(n_488),
.Y(n_691)
);

INVxp67_ASAP7_75t_SL g692 ( 
.A(n_618),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_536),
.B(n_490),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_596),
.B(n_601),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_620),
.B(n_264),
.Y(n_696)
);

AND2x2_ASAP7_75t_SL g697 ( 
.A(n_612),
.B(n_504),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_620),
.B(n_266),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_565),
.B(n_271),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_654),
.B(n_271),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_626),
.B(n_581),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_655),
.B(n_496),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_575),
.B(n_422),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_605),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_571),
.B(n_498),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_551),
.B(n_423),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_623),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_623),
.Y(n_708)
);

OAI221xp5_ASAP7_75t_L g709 ( 
.A1(n_638),
.A2(n_433),
.B1(n_354),
.B2(n_332),
.C(n_286),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_537),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_616),
.B(n_431),
.Y(n_711)
);

AO221x1_ASAP7_75t_L g712 ( 
.A1(n_537),
.A2(n_504),
.B1(n_520),
.B2(n_463),
.C(n_387),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_577),
.B(n_503),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_531),
.B(n_515),
.Y(n_714)
);

INVx4_ASAP7_75t_L g715 ( 
.A(n_535),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_606),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_541),
.B(n_436),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_542),
.B(n_515),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_545),
.B(n_527),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_550),
.B(n_527),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_555),
.B(n_436),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_607),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_559),
.B(n_561),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_586),
.Y(n_724)
);

OAI22xp33_ASAP7_75t_L g725 ( 
.A1(n_546),
.A2(n_406),
.B1(n_367),
.B2(n_387),
.Y(n_725)
);

OAI22x1_ASAP7_75t_SL g726 ( 
.A1(n_597),
.A2(n_406),
.B1(n_367),
.B2(n_391),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_608),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_548),
.B(n_553),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_553),
.B(n_438),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_564),
.B(n_441),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_553),
.B(n_441),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_617),
.A2(n_391),
.B1(n_395),
.B2(n_287),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_616),
.B(n_443),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_537),
.B(n_249),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_593),
.B(n_610),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_616),
.A2(n_283),
.B1(n_289),
.B2(n_284),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_618),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_562),
.B(n_445),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_593),
.B(n_252),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_562),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_636),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_535),
.B(n_582),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_582),
.B(n_250),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_557),
.B(n_287),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_557),
.A2(n_291),
.B1(n_309),
.B2(n_304),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_544),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_639),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_625),
.B(n_279),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_641),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_642),
.Y(n_750)
);

XNOR2xp5_ASAP7_75t_L g751 ( 
.A(n_597),
.B(n_395),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_644),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_583),
.B(n_526),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_645),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_587),
.B(n_473),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_609),
.A2(n_619),
.B1(n_647),
.B2(n_614),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_587),
.B(n_473),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_591),
.B(n_292),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_651),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_652),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_657),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_560),
.B(n_512),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_595),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_560),
.B(n_512),
.Y(n_764)
);

XOR2xp5_ASAP7_75t_L g765 ( 
.A(n_622),
.B(n_299),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_603),
.B(n_384),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_549),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_613),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_609),
.B(n_308),
.C(n_301),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_637),
.B(n_310),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_613),
.B(n_16),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_621),
.B(n_364),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_628),
.B(n_293),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_572),
.B(n_312),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_572),
.B(n_386),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_552),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_578),
.B(n_295),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_552),
.Y(n_778)
);

OR2x2_ASAP7_75t_L g779 ( 
.A(n_578),
.B(n_318),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_602),
.B(n_296),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_602),
.B(n_300),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_556),
.B(n_326),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_SL g783 ( 
.A(n_556),
.B(n_330),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_558),
.B(n_307),
.Y(n_784)
);

OR2x6_ASAP7_75t_L g785 ( 
.A(n_563),
.B(n_298),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_566),
.Y(n_786)
);

AO221x1_ASAP7_75t_L g787 ( 
.A1(n_566),
.A2(n_321),
.B1(n_319),
.B2(n_259),
.C(n_323),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_569),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_569),
.B(n_381),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_570),
.B(n_382),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_570),
.B(n_383),
.Y(n_791)
);

NAND2x1_ASAP7_75t_L g792 ( 
.A(n_573),
.B(n_385),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_580),
.A2(n_334),
.B1(n_341),
.B2(n_329),
.C(n_328),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_584),
.B(n_397),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_529),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_529),
.B(n_317),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_530),
.B(n_320),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_530),
.B(n_399),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_532),
.B(n_324),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_533),
.B(n_336),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_533),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_534),
.B(n_338),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_538),
.B(n_342),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_540),
.B(n_403),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_547),
.B(n_404),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_585),
.B(n_407),
.Y(n_806)
);

INVx8_ASAP7_75t_L g807 ( 
.A(n_568),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_666),
.B(n_335),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_666),
.Y(n_809)
);

O2A1O1Ixp33_ASAP7_75t_SL g810 ( 
.A1(n_670),
.A2(n_429),
.B(n_430),
.C(n_411),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_740),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_753),
.A2(n_757),
.B(n_755),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_674),
.A2(n_744),
.B1(n_683),
.B2(n_662),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_691),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_693),
.Y(n_815)
);

AOI222xp33_ASAP7_75t_L g816 ( 
.A1(n_726),
.A2(n_380),
.B1(n_388),
.B2(n_394),
.C1(n_370),
.C2(n_405),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_686),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_664),
.B(n_735),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_680),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_660),
.B(n_337),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_660),
.B(n_339),
.Y(n_821)
);

O2A1O1Ixp5_ASAP7_75t_L g822 ( 
.A1(n_694),
.A2(n_355),
.B(n_363),
.C(n_343),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_715),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_663),
.B(n_360),
.Y(n_824)
);

AO21x1_ASAP7_75t_L g825 ( 
.A1(n_764),
.A2(n_419),
.B(n_415),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_663),
.B(n_362),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_750),
.B(n_658),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_701),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_675),
.B(n_365),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_721),
.B(n_366),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_734),
.B(n_369),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_687),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_732),
.B(n_373),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_707),
.B(n_347),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_721),
.B(n_374),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_756),
.A2(n_434),
.B1(n_442),
.B2(n_421),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_714),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_730),
.B(n_375),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_714),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_688),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_692),
.A2(n_444),
.B1(n_306),
.B2(n_357),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_738),
.B(n_400),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_675),
.B(n_409),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_679),
.B(n_259),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_718),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_718),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_751),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_672),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_707),
.B(n_348),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_725),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_690),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_672),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_678),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_746),
.B(n_16),
.Y(n_854)
);

NOR2x2_ASAP7_75t_L g855 ( 
.A(n_712),
.B(n_410),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_738),
.B(n_413),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_723),
.A2(n_627),
.B(n_624),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_676),
.B(n_414),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_716),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_682),
.B(n_349),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_739),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_741),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_669),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_724),
.B(n_352),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_702),
.B(n_356),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_717),
.B(n_358),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_708),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_705),
.B(n_368),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_745),
.B(n_371),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_728),
.B(n_376),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_736),
.B(n_377),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_737),
.A2(n_319),
.B(n_321),
.C(n_259),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_681),
.A2(n_634),
.B(n_633),
.Y(n_873)
);

INVx1_ASAP7_75t_SL g874 ( 
.A(n_696),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_733),
.B(n_393),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_685),
.A2(n_634),
.B(n_633),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_747),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_699),
.B(n_396),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_710),
.B(n_319),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_703),
.B(n_401),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_754),
.B(n_759),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_713),
.A2(n_646),
.B(n_640),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_709),
.B(n_417),
.C(n_412),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_761),
.B(n_418),
.Y(n_884)
);

AOI21xp33_ASAP7_75t_L g885 ( 
.A1(n_769),
.A2(n_476),
.B(n_474),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_719),
.A2(n_476),
.B1(n_653),
.B2(n_650),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_720),
.A2(n_476),
.B1(n_648),
.B2(n_656),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_720),
.A2(n_476),
.B1(n_648),
.B2(n_604),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_704),
.B(n_722),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_727),
.B(n_673),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_749),
.B(n_18),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_752),
.B(n_19),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_697),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_782),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_760),
.B(n_19),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_768),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_661),
.A2(n_649),
.B(n_604),
.C(n_588),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_765),
.B(n_20),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_792),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_698),
.B(n_20),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_774),
.B(n_21),
.Y(n_901)
);

INVxp67_ASAP7_75t_L g902 ( 
.A(n_770),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_779),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_772),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_711),
.A2(n_649),
.B1(n_25),
.B2(n_26),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_785),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_667),
.B(n_671),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_798),
.A2(n_137),
.B(n_136),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_665),
.B(n_24),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_783),
.B(n_27),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_793),
.B(n_29),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_775),
.B(n_31),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_798),
.A2(n_146),
.B(n_145),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_768),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_804),
.A2(n_151),
.B(n_147),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_763),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_748),
.B(n_32),
.Y(n_917)
);

BUFx8_ASAP7_75t_SL g918 ( 
.A(n_785),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_668),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_729),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_731),
.A2(n_37),
.B(n_39),
.C(n_40),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_766),
.B(n_41),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_771),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_743),
.Y(n_924)
);

NOR2x1_ASAP7_75t_L g925 ( 
.A(n_758),
.B(n_43),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_773),
.B(n_44),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_706),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_927)
);

AND2x2_ASAP7_75t_SL g928 ( 
.A(n_742),
.B(n_50),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_777),
.B(n_56),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_695),
.B(n_56),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_789),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_L g932 ( 
.A(n_780),
.B(n_58),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_789),
.A2(n_60),
.B(n_61),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_L g934 ( 
.A1(n_790),
.A2(n_60),
.B(n_62),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_781),
.B(n_62),
.Y(n_935)
);

NOR2xp67_ASAP7_75t_L g936 ( 
.A(n_790),
.B(n_63),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_791),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_695),
.B(n_70),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_787),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_806),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_803),
.A2(n_784),
.B1(n_797),
.B2(n_684),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_794),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_807),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_807),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_794),
.B(n_71),
.Y(n_945)
);

NOR3xp33_ASAP7_75t_L g946 ( 
.A(n_677),
.B(n_72),
.C(n_73),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_805),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_689),
.B(n_72),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_700),
.B(n_74),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_800),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_786),
.B(n_75),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_788),
.B(n_75),
.Y(n_952)
);

BUFx2_ASAP7_75t_L g953 ( 
.A(n_802),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_796),
.B(n_799),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_767),
.B(n_77),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_776),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_778),
.A2(n_79),
.B(n_84),
.C(n_85),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_862),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_861),
.B(n_850),
.Y(n_959)
);

AO31x2_ASAP7_75t_L g960 ( 
.A1(n_825),
.A2(n_801),
.A3(n_795),
.B(n_88),
.Y(n_960)
);

INVxp67_ASAP7_75t_L g961 ( 
.A(n_828),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_827),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_831),
.B(n_86),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_889),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_889),
.Y(n_965)
);

INVx6_ASAP7_75t_SL g966 ( 
.A(n_929),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_903),
.B(n_92),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_863),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_918),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_943),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_881),
.A2(n_97),
.B1(n_103),
.B2(n_104),
.Y(n_971)
);

OAI22x1_ASAP7_75t_L g972 ( 
.A1(n_813),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_902),
.B(n_105),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_833),
.B(n_109),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_904),
.B(n_111),
.Y(n_975)
);

AND2x2_ASAP7_75t_SL g976 ( 
.A(n_928),
.B(n_113),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_817),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_848),
.B(n_114),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_832),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_840),
.Y(n_980)
);

OAI22xp33_ASAP7_75t_L g981 ( 
.A1(n_808),
.A2(n_947),
.B1(n_819),
.B2(n_911),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_877),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_851),
.Y(n_983)
);

AO21x1_ASAP7_75t_L g984 ( 
.A1(n_908),
.A2(n_915),
.B(n_913),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_874),
.B(n_894),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_901),
.A2(n_942),
.B(n_912),
.C(n_900),
.Y(n_986)
);

BUFx2_ASAP7_75t_SL g987 ( 
.A(n_848),
.Y(n_987)
);

AOI21x1_ASAP7_75t_L g988 ( 
.A1(n_888),
.A2(n_939),
.B(n_954),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_859),
.Y(n_989)
);

NOR2x1_ASAP7_75t_R g990 ( 
.A(n_852),
.B(n_893),
.Y(n_990)
);

CKINVDCx6p67_ASAP7_75t_R g991 ( 
.A(n_852),
.Y(n_991)
);

BUFx3_ASAP7_75t_L g992 ( 
.A(n_853),
.Y(n_992)
);

NAND3xp33_ASAP7_75t_SL g993 ( 
.A(n_816),
.B(n_883),
.C(n_919),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_814),
.B(n_815),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_836),
.B(n_820),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_924),
.B(n_898),
.Y(n_996)
);

OAI21xp5_ASAP7_75t_L g997 ( 
.A1(n_940),
.A2(n_857),
.B(n_907),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_906),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_909),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_821),
.B(n_824),
.Y(n_1000)
);

OAI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_907),
.A2(n_872),
.B(n_882),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_826),
.B(n_842),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_909),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_856),
.B(n_830),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_900),
.A2(n_945),
.B(n_811),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_835),
.B(n_838),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_929),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_884),
.A2(n_860),
.B(n_876),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_896),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_858),
.B(n_911),
.Y(n_1010)
);

OAI21xp33_ASAP7_75t_L g1011 ( 
.A1(n_933),
.A2(n_934),
.B(n_922),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_953),
.B(n_950),
.Y(n_1012)
);

AO31x2_ASAP7_75t_L g1013 ( 
.A1(n_841),
.A2(n_897),
.A3(n_887),
.B(n_886),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_873),
.A2(n_916),
.B(n_875),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_879),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_868),
.B(n_865),
.Y(n_1016)
);

OAI22x1_ASAP7_75t_L g1017 ( 
.A1(n_923),
.A2(n_847),
.B1(n_956),
.B2(n_925),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_936),
.Y(n_1018)
);

AO21x2_ASAP7_75t_L g1019 ( 
.A1(n_885),
.A2(n_930),
.B(n_938),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_917),
.B(n_844),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_926),
.B(n_869),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_810),
.A2(n_878),
.B(n_880),
.Y(n_1022)
);

OAI22x1_ASAP7_75t_L g1023 ( 
.A1(n_829),
.A2(n_843),
.B1(n_927),
.B2(n_932),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_914),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_891),
.A2(n_895),
.B(n_892),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_892),
.A2(n_895),
.B(n_951),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_866),
.B(n_935),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_951),
.A2(n_952),
.B(n_905),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_914),
.Y(n_1029)
);

AOI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_864),
.A2(n_871),
.B(n_870),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_885),
.A2(n_949),
.B(n_948),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_899),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_931),
.A2(n_937),
.B1(n_955),
.B2(n_957),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_841),
.B(n_946),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_867),
.Y(n_1035)
);

NOR2x1_ASAP7_75t_R g1036 ( 
.A(n_910),
.B(n_855),
.Y(n_1036)
);

AO21x1_ASAP7_75t_L g1037 ( 
.A1(n_941),
.A2(n_834),
.B(n_849),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_854),
.B(n_867),
.Y(n_1038)
);

INVxp67_ASAP7_75t_L g1039 ( 
.A(n_809),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_809),
.B(n_903),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_809),
.B(n_666),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_848),
.B(n_852),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_809),
.B(n_666),
.Y(n_1043)
);

OAI22x1_ASAP7_75t_L g1044 ( 
.A1(n_850),
.A2(n_520),
.B1(n_732),
.B2(n_659),
.Y(n_1044)
);

NAND3xp33_ASAP7_75t_L g1045 ( 
.A(n_822),
.B(n_921),
.C(n_920),
.Y(n_1045)
);

OR2x6_ASAP7_75t_L g1046 ( 
.A(n_848),
.B(n_852),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_837),
.A2(n_845),
.B1(n_846),
.B2(n_839),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_809),
.B(n_666),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_862),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_837),
.A2(n_845),
.B1(n_846),
.B2(n_839),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_809),
.B(n_666),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_918),
.B(n_589),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_809),
.B(n_666),
.Y(n_1053)
);

AOI21xp33_ASAP7_75t_L g1054 ( 
.A1(n_818),
.A2(n_659),
.B(n_660),
.Y(n_1054)
);

AOI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_818),
.A2(n_809),
.B1(n_674),
.B2(n_744),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_848),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_SL g1057 ( 
.A1(n_809),
.A2(n_710),
.B(n_732),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_809),
.B(n_600),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_809),
.B(n_666),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_862),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_837),
.A2(n_845),
.B1(n_846),
.B2(n_839),
.Y(n_1061)
);

NAND2x1p5_ASAP7_75t_L g1062 ( 
.A(n_943),
.B(n_944),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_809),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_809),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_861),
.B(n_659),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_809),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_809),
.B(n_666),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_809),
.B(n_903),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_809),
.B(n_666),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_918),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_818),
.B(n_659),
.Y(n_1071)
);

NOR2xp67_ASAP7_75t_L g1072 ( 
.A(n_809),
.B(n_660),
.Y(n_1072)
);

AND2x2_ASAP7_75t_SL g1073 ( 
.A(n_928),
.B(n_674),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_809),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_809),
.B(n_666),
.Y(n_1075)
);

NAND3xp33_ASAP7_75t_L g1076 ( 
.A(n_822),
.B(n_921),
.C(n_920),
.Y(n_1076)
);

AO221x2_ASAP7_75t_L g1077 ( 
.A1(n_931),
.A2(n_520),
.B1(n_725),
.B2(n_937),
.C(n_511),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_837),
.A2(n_845),
.B1(n_846),
.B2(n_839),
.Y(n_1078)
);

AOI21xp33_ASAP7_75t_L g1079 ( 
.A1(n_818),
.A2(n_659),
.B(n_660),
.Y(n_1079)
);

AND2x6_ASAP7_75t_SL g1080 ( 
.A(n_898),
.B(n_554),
.Y(n_1080)
);

AND2x4_ASAP7_75t_L g1081 ( 
.A(n_809),
.B(n_903),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_SL g1082 ( 
.A1(n_881),
.A2(n_890),
.B(n_889),
.Y(n_1082)
);

NAND2x1_ASAP7_75t_L g1083 ( 
.A(n_823),
.B(n_715),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_861),
.B(n_659),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_809),
.B(n_666),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_809),
.B(n_903),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_825),
.A2(n_812),
.A3(n_764),
.B(n_762),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_809),
.B(n_666),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_809),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_818),
.B(n_659),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_809),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1058),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1057),
.B(n_959),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_SL g1094 ( 
.A1(n_1082),
.A2(n_1050),
.B(n_1047),
.Y(n_1094)
);

AOI22x1_ASAP7_75t_L g1095 ( 
.A1(n_1017),
.A2(n_1023),
.B1(n_1022),
.B2(n_1008),
.Y(n_1095)
);

AO21x2_ASAP7_75t_L g1096 ( 
.A1(n_984),
.A2(n_988),
.B(n_1028),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_970),
.Y(n_1097)
);

BUFx2_ASAP7_75t_SL g1098 ( 
.A(n_970),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_964),
.B(n_965),
.Y(n_1099)
);

AOI221xp5_ASAP7_75t_L g1100 ( 
.A1(n_1071),
.A2(n_1090),
.B1(n_1079),
.B2(n_1054),
.C(n_1044),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1072),
.B(n_1039),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_1077),
.A2(n_1050),
.B1(n_1061),
.B2(n_1047),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_962),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1061),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1057),
.B(n_993),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1041),
.B(n_1043),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_986),
.A2(n_1072),
.B(n_1000),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1063),
.B(n_1064),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_1078),
.Y(n_1109)
);

OR3x4_ASAP7_75t_SL g1110 ( 
.A(n_1036),
.B(n_1080),
.C(n_1077),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1078),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_987),
.B(n_978),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_976),
.A2(n_1073),
.B1(n_1040),
.B2(n_1068),
.Y(n_1113)
);

BUFx2_ASAP7_75t_R g1114 ( 
.A(n_1070),
.Y(n_1114)
);

INVx4_ASAP7_75t_SL g1115 ( 
.A(n_978),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_978),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1048),
.B(n_1051),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_1056),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1053),
.B(n_1059),
.Y(n_1119)
);

AO21x2_ASAP7_75t_L g1120 ( 
.A1(n_1028),
.A2(n_1026),
.B(n_1025),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_1066),
.B(n_1074),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_1011),
.A2(n_1001),
.B(n_1031),
.Y(n_1122)
);

BUFx2_ASAP7_75t_R g1123 ( 
.A(n_1065),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1067),
.B(n_1069),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1089),
.B(n_1091),
.Y(n_1125)
);

AND2x4_ASAP7_75t_L g1126 ( 
.A(n_1040),
.B(n_1068),
.Y(n_1126)
);

BUFx8_ASAP7_75t_L g1127 ( 
.A(n_999),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_995),
.A2(n_1010),
.B1(n_1033),
.B2(n_1034),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1007),
.B(n_1081),
.Y(n_1129)
);

OA21x2_ASAP7_75t_L g1130 ( 
.A1(n_1005),
.A2(n_997),
.B(n_1014),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1084),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1081),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1086),
.B(n_1075),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1086),
.B(n_1002),
.Y(n_1134)
);

CKINVDCx14_ASAP7_75t_R g1135 ( 
.A(n_969),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_1006),
.B(n_1003),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_1019),
.A2(n_1076),
.B(n_1045),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1042),
.B(n_1046),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_985),
.B(n_1012),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_977),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1004),
.A2(n_1016),
.B(n_1027),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_979),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_1012),
.B(n_961),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_980),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_996),
.B(n_981),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_983),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_989),
.Y(n_1148)
);

AO31x2_ASAP7_75t_L g1149 ( 
.A1(n_1037),
.A2(n_971),
.A3(n_972),
.B(n_975),
.Y(n_1149)
);

BUFx2_ASAP7_75t_L g1150 ( 
.A(n_966),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_994),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_992),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1038),
.A2(n_1018),
.B(n_1020),
.Y(n_1153)
);

INVx2_ASAP7_75t_SL g1154 ( 
.A(n_991),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1055),
.A2(n_967),
.B1(n_974),
.B2(n_1052),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1052),
.B(n_990),
.Y(n_1157)
);

OR3x4_ASAP7_75t_SL g1158 ( 
.A(n_1036),
.B(n_1080),
.C(n_990),
.Y(n_1158)
);

CKINVDCx11_ASAP7_75t_R g1159 ( 
.A(n_1042),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1021),
.B(n_973),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1042),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_958),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1030),
.A2(n_1013),
.B(n_963),
.Y(n_1163)
);

OA21x2_ASAP7_75t_L g1164 ( 
.A1(n_982),
.A2(n_1060),
.B(n_1049),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_1062),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1046),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_967),
.B(n_998),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_1009),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1083),
.A2(n_1035),
.B(n_1013),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_968),
.B(n_1015),
.Y(n_1170)
);

AO22x2_ASAP7_75t_L g1171 ( 
.A1(n_1015),
.A2(n_960),
.B1(n_1013),
.B2(n_1032),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1024),
.A2(n_1029),
.B(n_1087),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1087),
.A2(n_960),
.B(n_1046),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_964),
.B(n_965),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1058),
.B(n_600),
.Y(n_1175)
);

AND2x6_ASAP7_75t_L g1176 ( 
.A(n_964),
.B(n_965),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_1047),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1058),
.B(n_600),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_1047),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1058),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1058),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1058),
.B(n_600),
.Y(n_1182)
);

BUFx2_ASAP7_75t_SL g1183 ( 
.A(n_970),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_964),
.B(n_965),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1058),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1047),
.A2(n_1061),
.B1(n_1078),
.B2(n_1050),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1065),
.Y(n_1187)
);

INVx6_ASAP7_75t_L g1188 ( 
.A(n_970),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_970),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_970),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1058),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1151),
.B(n_1106),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1105),
.A2(n_1093),
.B1(n_1146),
.B2(n_1100),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1131),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1175),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1094),
.Y(n_1196)
);

AOI222xp33_ASAP7_75t_L g1197 ( 
.A1(n_1142),
.A2(n_1105),
.B1(n_1160),
.B2(n_1134),
.C1(n_1146),
.C2(n_1093),
.Y(n_1197)
);

HB1xp67_ASAP7_75t_L g1198 ( 
.A(n_1187),
.Y(n_1198)
);

CKINVDCx6p67_ASAP7_75t_R g1199 ( 
.A(n_1118),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1152),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1102),
.A2(n_1186),
.B1(n_1112),
.B2(n_1134),
.Y(n_1201)
);

BUFx12f_ASAP7_75t_L g1202 ( 
.A(n_1118),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1099),
.B(n_1128),
.Y(n_1203)
);

CKINVDCx14_ASAP7_75t_R g1204 ( 
.A(n_1135),
.Y(n_1204)
);

BUFx2_ASAP7_75t_SL g1205 ( 
.A(n_1176),
.Y(n_1205)
);

HB1xp67_ASAP7_75t_L g1206 ( 
.A(n_1133),
.Y(n_1206)
);

INVx2_ASAP7_75t_SL g1207 ( 
.A(n_1188),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1115),
.B(n_1176),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1176),
.Y(n_1209)
);

BUFx2_ASAP7_75t_R g1210 ( 
.A(n_1098),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1133),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1135),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1112),
.A2(n_1156),
.B1(n_1104),
.B2(n_1111),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1112),
.A2(n_1128),
.B1(n_1133),
.B2(n_1107),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1117),
.B(n_1119),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1159),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1176),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1115),
.A2(n_1160),
.B1(n_1101),
.B2(n_1176),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1168),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1168),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1104),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1103),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1092),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1140),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1189),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1099),
.B(n_1108),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1168),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1116),
.A2(n_1157),
.B1(n_1177),
.B2(n_1111),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1115),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1095),
.B(n_1113),
.C(n_1136),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1099),
.B(n_1108),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1120),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1108),
.B(n_1121),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1173),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1109),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1109),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1177),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1179),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1121),
.B(n_1125),
.Y(n_1239)
);

BUFx3_ASAP7_75t_L g1240 ( 
.A(n_1189),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_1190),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1159),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1124),
.A2(n_1139),
.B1(n_1138),
.B2(n_1166),
.Y(n_1243)
);

BUFx12f_ASAP7_75t_L g1244 ( 
.A(n_1116),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1164),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1164),
.Y(n_1246)
);

OR2x6_ASAP7_75t_L g1247 ( 
.A(n_1138),
.B(n_1183),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1168),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1180),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1121),
.B(n_1125),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1174),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1184),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1213),
.B(n_1163),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1245),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1245),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1203),
.B(n_1163),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1225),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1246),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1208),
.B(n_1169),
.Y(n_1259)
);

INVxp67_ASAP7_75t_SL g1260 ( 
.A(n_1251),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1208),
.B(n_1172),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1203),
.B(n_1171),
.Y(n_1262)
);

OR2x2_ASAP7_75t_L g1263 ( 
.A(n_1221),
.B(n_1137),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1233),
.B(n_1171),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1233),
.B(n_1171),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1251),
.B(n_1181),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1239),
.B(n_1137),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1239),
.B(n_1250),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1252),
.B(n_1185),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1219),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1194),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1205),
.B(n_1138),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1250),
.B(n_1096),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1198),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1208),
.B(n_1096),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_1252),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1226),
.B(n_1122),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1226),
.B(n_1122),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1231),
.B(n_1122),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1231),
.B(n_1130),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1197),
.A2(n_1101),
.B1(n_1126),
.B2(n_1136),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1217),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1217),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1215),
.B(n_1191),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1192),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1221),
.B(n_1149),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1224),
.B(n_1125),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1205),
.A2(n_1217),
.B1(n_1204),
.B2(n_1229),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1225),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1235),
.B(n_1149),
.Y(n_1290)
);

OR2x2_ASAP7_75t_L g1291 ( 
.A(n_1236),
.B(n_1149),
.Y(n_1291)
);

BUFx3_ASAP7_75t_L g1292 ( 
.A(n_1240),
.Y(n_1292)
);

BUFx4f_ASAP7_75t_SL g1293 ( 
.A(n_1202),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1218),
.A2(n_1101),
.B1(n_1123),
.B2(n_1166),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1219),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1193),
.A2(n_1126),
.B1(n_1129),
.B2(n_1144),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1209),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1202),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1296),
.A2(n_1214),
.B1(n_1281),
.B2(n_1201),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1254),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1257),
.Y(n_1301)
);

OAI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1260),
.A2(n_1228),
.B(n_1230),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1254),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1255),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1280),
.B(n_1232),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1296),
.A2(n_1243),
.B1(n_1216),
.B2(n_1206),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1261),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1267),
.B(n_1237),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1258),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1276),
.Y(n_1310)
);

BUFx3_ASAP7_75t_L g1311 ( 
.A(n_1257),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1275),
.B(n_1234),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1294),
.A2(n_1216),
.B1(n_1211),
.B2(n_1196),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1293),
.B(n_1199),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1273),
.A2(n_1196),
.B1(n_1195),
.B2(n_1229),
.Y(n_1315)
);

INVxp67_ASAP7_75t_SL g1316 ( 
.A(n_1289),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1298),
.B(n_1199),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1285),
.B(n_1222),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1271),
.B(n_1223),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1267),
.B(n_1238),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1280),
.B(n_1232),
.Y(n_1321)
);

AND2x4_ASAP7_75t_SL g1322 ( 
.A(n_1272),
.B(n_1229),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1274),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1292),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1266),
.B(n_1249),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1272),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_SL g1327 ( 
.A(n_1326),
.B(n_1310),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1305),
.B(n_1277),
.Y(n_1328)
);

INVxp33_ASAP7_75t_L g1329 ( 
.A(n_1317),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1300),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1305),
.B(n_1256),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1300),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1303),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1321),
.B(n_1277),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1321),
.B(n_1256),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1307),
.B(n_1278),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1308),
.B(n_1263),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1304),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1307),
.B(n_1278),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1299),
.A2(n_1262),
.B1(n_1273),
.B2(n_1264),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1307),
.B(n_1279),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1307),
.B(n_1279),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1311),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1312),
.B(n_1262),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1309),
.B(n_1290),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1310),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1330),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1328),
.B(n_1264),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1337),
.B(n_1308),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1330),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1327),
.A2(n_1302),
.B(n_1272),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1338),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1340),
.B(n_1323),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1337),
.B(n_1331),
.Y(n_1354)
);

NOR2x1p5_ASAP7_75t_SL g1355 ( 
.A(n_1338),
.B(n_1286),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1327),
.A2(n_1306),
.B1(n_1313),
.B2(n_1302),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1332),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1346),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1332),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1333),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1343),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1331),
.B(n_1320),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1328),
.B(n_1316),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1333),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1338),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1328),
.B(n_1319),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1334),
.B(n_1265),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1354),
.B(n_1334),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1351),
.B(n_1298),
.Y(n_1369)
);

AOI321xp33_ASAP7_75t_L g1370 ( 
.A1(n_1353),
.A2(n_1346),
.A3(n_1315),
.B1(n_1336),
.B2(n_1342),
.C(n_1339),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1349),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1349),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1354),
.B(n_1334),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1361),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1356),
.A2(n_1326),
.B1(n_1272),
.B2(n_1343),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1348),
.B(n_1335),
.Y(n_1376)
);

OAI32xp33_ASAP7_75t_L g1377 ( 
.A1(n_1363),
.A2(n_1329),
.A3(n_1212),
.B1(n_1324),
.B2(n_1326),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1347),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1358),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1362),
.A2(n_1326),
.B1(n_1288),
.B2(n_1272),
.Y(n_1380)
);

OAI222xp33_ASAP7_75t_L g1381 ( 
.A1(n_1361),
.A2(n_1301),
.B1(n_1282),
.B2(n_1247),
.C1(n_1335),
.C2(n_1344),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1352),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1348),
.B(n_1367),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1366),
.A2(n_1336),
.B1(n_1342),
.B2(n_1339),
.Y(n_1384)
);

NAND2x2_ASAP7_75t_L g1385 ( 
.A(n_1362),
.B(n_1158),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1347),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_SL g1387 ( 
.A1(n_1367),
.A2(n_1314),
.B1(n_1242),
.B2(n_1311),
.Y(n_1387)
);

AOI21xp33_ASAP7_75t_L g1388 ( 
.A1(n_1375),
.A2(n_1301),
.B(n_1318),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1387),
.A2(n_1322),
.B1(n_1311),
.B2(n_1282),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1380),
.A2(n_1344),
.B1(n_1341),
.B2(n_1336),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1382),
.Y(n_1391)
);

OAI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1369),
.A2(n_1283),
.B1(n_1247),
.B2(n_1209),
.Y(n_1392)
);

AOI21xp33_ASAP7_75t_L g1393 ( 
.A1(n_1375),
.A2(n_1200),
.B(n_1242),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1377),
.A2(n_1342),
.B1(n_1339),
.B2(n_1341),
.C(n_1110),
.Y(n_1394)
);

OAI322xp33_ASAP7_75t_L g1395 ( 
.A1(n_1379),
.A2(n_1350),
.A3(n_1364),
.B1(n_1360),
.B2(n_1357),
.C1(n_1359),
.C2(n_1253),
.Y(n_1395)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1396 ( 
.A1(n_1370),
.A2(n_1110),
.B(n_1158),
.C(n_1325),
.D(n_1287),
.Y(n_1396)
);

XNOR2xp5_ASAP7_75t_L g1397 ( 
.A(n_1371),
.B(n_1154),
.Y(n_1397)
);

OA21x2_ASAP7_75t_L g1398 ( 
.A1(n_1379),
.A2(n_1365),
.B(n_1352),
.Y(n_1398)
);

AOI31xp33_ASAP7_75t_L g1399 ( 
.A1(n_1394),
.A2(n_1385),
.A3(n_1210),
.B(n_1114),
.Y(n_1399)
);

NOR3xp33_ASAP7_75t_L g1400 ( 
.A(n_1393),
.B(n_1381),
.C(n_1155),
.Y(n_1400)
);

AOI211xp5_ASAP7_75t_L g1401 ( 
.A1(n_1388),
.A2(n_1381),
.B(n_1374),
.C(n_1372),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1390),
.A2(n_1384),
.B1(n_1368),
.B2(n_1385),
.C(n_1373),
.Y(n_1402)
);

AOI21xp33_ASAP7_75t_L g1403 ( 
.A1(n_1397),
.A2(n_1284),
.B(n_1150),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1391),
.B(n_1376),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1398),
.A2(n_1247),
.B(n_1292),
.Y(n_1405)
);

OAI22x1_ASAP7_75t_L g1406 ( 
.A1(n_1398),
.A2(n_1396),
.B1(n_1389),
.B2(n_1283),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1395),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1396),
.A2(n_1392),
.B1(n_1244),
.B2(n_1268),
.Y(n_1408)
);

AOI21xp33_ASAP7_75t_L g1409 ( 
.A1(n_1394),
.A2(n_1244),
.B(n_1161),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1396),
.A2(n_1378),
.B(n_1386),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1397),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1397),
.B(n_1383),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1399),
.B(n_1322),
.Y(n_1413)
);

NOR3xp33_ASAP7_75t_L g1414 ( 
.A(n_1402),
.B(n_1097),
.C(n_1153),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1404),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1401),
.B(n_1127),
.C(n_1170),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_1411),
.B(n_1345),
.Y(n_1417)
);

NOR3xp33_ASAP7_75t_L g1418 ( 
.A(n_1400),
.B(n_1097),
.C(n_1167),
.Y(n_1418)
);

AND3x1_ASAP7_75t_L g1419 ( 
.A(n_1408),
.B(n_1283),
.C(n_1297),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_SL g1420 ( 
.A(n_1406),
.B(n_1365),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1408),
.A2(n_1312),
.B1(n_1275),
.B2(n_1247),
.Y(n_1421)
);

NAND3xp33_ASAP7_75t_L g1422 ( 
.A(n_1407),
.B(n_1127),
.C(n_1170),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1415),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1422),
.B(n_1416),
.C(n_1414),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_L g1425 ( 
.A(n_1418),
.B(n_1409),
.C(n_1410),
.Y(n_1425)
);

NOR2x1_ASAP7_75t_L g1426 ( 
.A(n_1413),
.B(n_1405),
.Y(n_1426)
);

INVxp67_ASAP7_75t_SL g1427 ( 
.A(n_1417),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1421),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1420),
.B(n_1412),
.Y(n_1429)
);

NOR2x1_ASAP7_75t_L g1430 ( 
.A(n_1419),
.B(n_1190),
.Y(n_1430)
);

AOI211xp5_ASAP7_75t_L g1431 ( 
.A1(n_1422),
.A2(n_1403),
.B(n_1129),
.C(n_1269),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1422),
.B(n_1127),
.C(n_1240),
.Y(n_1432)
);

NOR3xp33_ASAP7_75t_L g1433 ( 
.A(n_1424),
.B(n_1182),
.C(n_1178),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1426),
.B(n_1241),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1423),
.Y(n_1435)
);

NOR3xp33_ASAP7_75t_L g1436 ( 
.A(n_1425),
.B(n_1207),
.C(n_1219),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1427),
.B(n_1355),
.Y(n_1437)
);

OAI322xp33_ASAP7_75t_L g1438 ( 
.A1(n_1429),
.A2(n_1286),
.A3(n_1132),
.B1(n_1253),
.B2(n_1291),
.C1(n_1290),
.C2(n_1345),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1432),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1430),
.B(n_1241),
.Y(n_1440)
);

NAND2x1p5_ASAP7_75t_L g1441 ( 
.A(n_1439),
.B(n_1220),
.Y(n_1441)
);

NAND4xp75_ASAP7_75t_L g1442 ( 
.A(n_1435),
.B(n_1428),
.C(n_1431),
.D(n_1207),
.Y(n_1442)
);

OAI322xp33_ASAP7_75t_L g1443 ( 
.A1(n_1437),
.A2(n_1145),
.A3(n_1143),
.B1(n_1147),
.B2(n_1148),
.C1(n_1141),
.C2(n_1291),
.Y(n_1443)
);

NOR2xp67_ASAP7_75t_L g1444 ( 
.A(n_1434),
.B(n_1220),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1436),
.A2(n_1275),
.B1(n_1259),
.B2(n_1312),
.Y(n_1445)
);

OA22x2_ASAP7_75t_L g1446 ( 
.A1(n_1445),
.A2(n_1433),
.B1(n_1440),
.B2(n_1438),
.Y(n_1446)
);

AOI22x1_ASAP7_75t_SL g1447 ( 
.A1(n_1442),
.A2(n_1227),
.B1(n_1248),
.B2(n_1220),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1446),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1448),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1449),
.A2(n_1441),
.B1(n_1444),
.B2(n_1447),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1450),
.A2(n_1443),
.B1(n_1188),
.B2(n_1270),
.Y(n_1451)
);

AOI221xp5_ASAP7_75t_L g1452 ( 
.A1(n_1451),
.A2(n_1165),
.B1(n_1248),
.B2(n_1227),
.C(n_1162),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1452),
.B(n_1268),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1453),
.B(n_1188),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1454),
.A2(n_1227),
.B1(n_1248),
.B2(n_1295),
.Y(n_1455)
);


endmodule