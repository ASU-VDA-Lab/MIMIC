module fake_jpeg_15205_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_12),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_41),
.Y(n_50)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_48),
.B1(n_53),
.B2(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_47),
.B(n_64),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_31),
.B1(n_22),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_36),
.B1(n_26),
.B2(n_37),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_33),
.C(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_35),
.B1(n_29),
.B2(n_27),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_54),
.B(n_20),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_35),
.B1(n_29),
.B2(n_27),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_21),
.Y(n_61)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_25),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_46),
.B1(n_48),
.B2(n_47),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_72),
.A2(n_86),
.B1(n_106),
.B2(n_36),
.Y(n_122)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_88),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_20),
.B1(n_34),
.B2(n_17),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_62),
.A2(n_20),
.B1(n_34),
.B2(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_85),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_36),
.B1(n_32),
.B2(n_30),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_32),
.B(n_30),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_36),
.B1(n_44),
.B2(n_42),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_91),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_33),
.B(n_24),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_100),
.Y(n_114)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_45),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_53),
.A2(n_36),
.B1(n_28),
.B2(n_42),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_45),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_66),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_50),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_110),
.B(n_113),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_50),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_69),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_117),
.B(n_131),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_125),
.C(n_45),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_128),
.B(n_84),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_122),
.A2(n_126),
.B1(n_134),
.B2(n_102),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_45),
.C(n_39),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_26),
.A3(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_87),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_72),
.A2(n_42),
.B1(n_44),
.B2(n_39),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_73),
.B1(n_94),
.B2(n_100),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_75),
.A2(n_42),
.B1(n_44),
.B2(n_39),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_33),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_137),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_128),
.B(n_110),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_157),
.B(n_165),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_24),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_140),
.B(n_141),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_112),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_155),
.B1(n_161),
.B2(n_37),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_112),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_145),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_151),
.B1(n_120),
.B2(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_102),
.B(n_75),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_139),
.B(n_165),
.Y(n_179)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_124),
.A2(n_99),
.B1(n_89),
.B2(n_88),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_2),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_122),
.A2(n_86),
.B1(n_44),
.B2(n_101),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_123),
.B1(n_133),
.B2(n_125),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_78),
.B1(n_98),
.B2(n_16),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_0),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_78),
.Y(n_160)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_166),
.C(n_6),
.Y(n_199)
);

AO21x1_ASAP7_75t_SL g161 ( 
.A1(n_109),
.A2(n_37),
.B(n_33),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_164),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_113),
.A2(n_33),
.B(n_24),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_104),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_108),
.B(n_96),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_90),
.Y(n_182)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_115),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_168),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_169),
.A2(n_171),
.B1(n_190),
.B2(n_151),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_173),
.B(n_175),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_129),
.B(n_126),
.C(n_136),
.D(n_120),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_142),
.A2(n_111),
.B1(n_132),
.B2(n_116),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_177),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_179),
.A2(n_186),
.B(n_143),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_111),
.B1(n_116),
.B2(n_37),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_129),
.C(n_121),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_185),
.C(n_196),
.Y(n_201)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_121),
.C(n_90),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_158),
.A2(n_83),
.B1(n_70),
.B2(n_43),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_8),
.B1(n_13),
.B2(n_12),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_190)
);

NOR2x1_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_7),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_9),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_6),
.C(n_11),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_200),
.C(n_145),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_137),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_210),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_195),
.A2(n_162),
.B(n_163),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_203),
.A2(n_217),
.B(n_8),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_144),
.C(n_157),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_206),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_215),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_196),
.C(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_144),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_175),
.B(n_146),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_216),
.B(n_224),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_149),
.B(n_147),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_197),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_159),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_222),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_194),
.B(n_164),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_5),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_198),
.B(n_192),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_141),
.C(n_140),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_156),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_187),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_169),
.A2(n_150),
.B1(n_3),
.B2(n_4),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_226),
.A2(n_186),
.B1(n_188),
.B2(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_222),
.A2(n_177),
.B1(n_183),
.B2(n_173),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_231),
.A2(n_233),
.B1(n_236),
.B2(n_237),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_208),
.A2(n_179),
.B1(n_189),
.B2(n_182),
.Y(n_233)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_207),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_212),
.A2(n_180),
.B1(n_3),
.B2(n_4),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_2),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_217),
.B(n_5),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_214),
.B1(n_213),
.B2(n_9),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_245),
.A2(n_237),
.B(n_230),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_227),
.A2(n_223),
.B(n_211),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_254),
.B(n_263),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_211),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_251),
.Y(n_273)
);

OA21x2_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_202),
.B(n_206),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_247),
.A2(n_224),
.B1(n_219),
.B2(n_226),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_201),
.B1(n_239),
.B2(n_245),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_231),
.A2(n_220),
.B1(n_225),
.B2(n_209),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_228),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_201),
.C(n_204),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_238),
.C(n_242),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_229),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_210),
.B(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_2),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_248),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_235),
.B1(n_233),
.B2(n_232),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_271),
.B1(n_272),
.B2(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_277),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_240),
.C(n_216),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_274),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_245),
.B1(n_236),
.B2(n_209),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_240),
.C(n_203),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_203),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_275),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_250),
.B(n_3),
.C(n_16),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_260),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_288),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_276),
.A2(n_249),
.B(n_263),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_259),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_264),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_287),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_251),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_252),
.B(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_264),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_255),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_291),
.B(n_253),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_281),
.A2(n_274),
.B1(n_253),
.B2(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_298),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_270),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_289),
.B1(n_283),
.B2(n_287),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_266),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_298),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_305),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_280),
.B(n_286),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_304),
.A2(n_296),
.B(n_297),
.Y(n_308)
);

NAND4xp25_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_11),
.C(n_16),
.D(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_306),
.B(n_301),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_309),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_303),
.Y(n_310)
);

FAx1_ASAP7_75t_SL g311 ( 
.A(n_310),
.B(n_305),
.CI(n_307),
.CON(n_311),
.SN(n_311)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_311),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_311),
.Y(n_315)
);


endmodule