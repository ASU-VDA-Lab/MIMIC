module fake_jpeg_27909_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_8),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_27),
.Y(n_43)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_41),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_21),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_16),
.B1(n_30),
.B2(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_53),
.B1(n_56),
.B2(n_20),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_49),
.Y(n_66)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_22),
.Y(n_60)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_34),
.A2(n_41),
.B(n_24),
.C(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_16),
.B1(n_29),
.B2(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_33),
.A2(n_16),
.B1(n_28),
.B2(n_18),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_20),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_22),
.Y(n_75)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_73),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_21),
.A3(n_24),
.B1(n_19),
.B2(n_31),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_47),
.CI(n_49),
.CON(n_77),
.SN(n_77)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_50),
.A2(n_20),
.B(n_25),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_43),
.C(n_31),
.Y(n_82)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_76),
.B(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_50),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_79),
.A2(n_23),
.B1(n_62),
.B2(n_22),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_15),
.B(n_73),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_84),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_57),
.C(n_54),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_72),
.C(n_66),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_86),
.Y(n_104)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_52),
.B1(n_45),
.B2(n_46),
.Y(n_90)
);

AO21x2_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_63),
.B(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_52),
.B1(n_45),
.B2(n_48),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_52),
.B1(n_61),
.B2(n_74),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_61),
.B(n_19),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_21),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_95),
.B(n_98),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_109),
.B1(n_83),
.B2(n_91),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_15),
.B1(n_25),
.B2(n_23),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_82),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_81),
.B(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_108),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_59),
.B1(n_62),
.B2(n_63),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_91),
.B1(n_83),
.B2(n_89),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_80),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_84),
.C(n_85),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_105),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_77),
.B(n_80),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_100),
.B(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_121),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_124),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_112),
.B1(n_123),
.B2(n_120),
.C(n_122),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_124),
.A2(n_109),
.B(n_110),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_77),
.C(n_13),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_132),
.B(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_116),
.B(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_136),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_109),
.A3(n_103),
.B1(n_97),
.B2(n_102),
.C1(n_101),
.C2(n_9),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_134),
.B(n_119),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_113),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_144),
.B(n_131),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_130),
.B1(n_121),
.B2(n_128),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_112),
.B1(n_123),
.B2(n_64),
.Y(n_145)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_146),
.B(n_150),
.Y(n_156)
);

AOI321xp33_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_131),
.A3(n_126),
.B1(n_129),
.B2(n_12),
.C(n_14),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_64),
.B1(n_3),
.B2(n_4),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_13),
.B(n_12),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_147),
.B(n_11),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_144),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_153),
.A2(n_154),
.B(n_156),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_143),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_157),
.B1(n_0),
.B2(n_3),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_149),
.B(n_143),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_11),
.B(n_3),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_158),
.A2(n_153),
.B1(n_6),
.B2(n_7),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_159),
.B(n_160),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_0),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_165),
.A2(n_161),
.B(n_6),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_164),
.C(n_6),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_166),
.Y(n_169)
);


endmodule