module real_aes_2212_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_153;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_210;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_0), .B(n_131), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g139 ( .A1(n_1), .A2(n_140), .B(n_145), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_2), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_3), .B(n_131), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_4), .B(n_147), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_5), .B(n_147), .Y(n_185) );
INVx1_ASAP7_75t_L g138 ( .A(n_6), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_7), .B(n_147), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g762 ( .A(n_8), .Y(n_762) );
NAND2xp33_ASAP7_75t_L g174 ( .A(n_9), .B(n_149), .Y(n_174) );
AND2x2_ASAP7_75t_L g484 ( .A(n_10), .B(n_168), .Y(n_484) );
AND2x2_ASAP7_75t_L g492 ( .A(n_11), .B(n_125), .Y(n_492) );
INVx2_ASAP7_75t_L g128 ( .A(n_12), .Y(n_128) );
AOI221x1_ASAP7_75t_L g220 ( .A1(n_13), .A2(n_24), .B1(n_131), .B2(n_140), .C(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_14), .B(n_147), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_15), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_16), .B(n_131), .Y(n_170) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_17), .A2(n_168), .B(n_169), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_18), .B(n_151), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_19), .B(n_147), .Y(n_161) );
AO21x1_ASAP7_75t_L g180 ( .A1(n_20), .A2(n_131), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_21), .B(n_131), .Y(n_465) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_23), .A2(n_89), .B1(n_131), .B2(n_500), .Y(n_499) );
NAND2x1_ASAP7_75t_L g193 ( .A(n_25), .B(n_147), .Y(n_193) );
NAND2x1_ASAP7_75t_L g212 ( .A(n_26), .B(n_149), .Y(n_212) );
AOI222xp33_ASAP7_75t_L g100 ( .A1(n_27), .A2(n_101), .B1(n_755), .B2(n_766), .C1(n_781), .C2(n_785), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_27), .A2(n_62), .B1(n_771), .B2(n_772), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_27), .Y(n_771) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_28), .A2(n_86), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g153 ( .A(n_28), .B(n_86), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_29), .B(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_30), .B(n_147), .Y(n_173) );
AO21x2_ASAP7_75t_L g439 ( .A1(n_31), .A2(n_125), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_32), .B(n_149), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_33), .A2(n_140), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_34), .B(n_147), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_35), .A2(n_140), .B(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g137 ( .A(n_36), .B(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g141 ( .A(n_36), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g508 ( .A(n_36), .Y(n_508) );
OR2x6_ASAP7_75t_L g112 ( .A(n_37), .B(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_38), .B(n_131), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_39), .B(n_131), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_40), .B(n_147), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_41), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_42), .B(n_149), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_43), .B(n_131), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_44), .A2(n_140), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_45), .A2(n_140), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_46), .B(n_149), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g102 ( .A1(n_47), .A2(n_50), .B1(n_103), .B2(n_104), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_47), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_48), .B(n_149), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g441 ( .A(n_49), .B(n_131), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_50), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_51), .Y(n_780) );
INVx1_ASAP7_75t_L g134 ( .A(n_52), .Y(n_134) );
INVx1_ASAP7_75t_L g144 ( .A(n_52), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_53), .B(n_147), .Y(n_490) );
AND2x2_ASAP7_75t_L g456 ( .A(n_54), .B(n_151), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_55), .B(n_149), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_56), .B(n_147), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_57), .B(n_149), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_58), .A2(n_140), .B(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_59), .B(n_131), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_60), .B(n_131), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_61), .A2(n_140), .B(n_449), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_62), .Y(n_772) );
AO21x1_ASAP7_75t_L g182 ( .A1(n_63), .A2(n_140), .B(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g471 ( .A(n_64), .B(n_152), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_65), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_66), .B(n_149), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_67), .B(n_131), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_68), .B(n_149), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_69), .A2(n_94), .B1(n_140), .B2(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g205 ( .A(n_70), .B(n_152), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_71), .B(n_147), .Y(n_468) );
INVx1_ASAP7_75t_L g136 ( .A(n_72), .Y(n_136) );
INVx1_ASAP7_75t_L g142 ( .A(n_72), .Y(n_142) );
AND2x2_ASAP7_75t_L g216 ( .A(n_73), .B(n_125), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_74), .B(n_149), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_75), .A2(n_140), .B(n_460), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_76), .A2(n_140), .B(n_529), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_77), .A2(n_140), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g453 ( .A(n_78), .B(n_152), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_79), .B(n_151), .Y(n_497) );
INVx1_ASAP7_75t_L g115 ( .A(n_80), .Y(n_115) );
AND2x2_ASAP7_75t_L g124 ( .A(n_81), .B(n_125), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_82), .B(n_131), .Y(n_163) );
AND2x2_ASAP7_75t_L g532 ( .A(n_83), .B(n_168), .Y(n_532) );
AND2x2_ASAP7_75t_L g181 ( .A(n_84), .B(n_157), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_85), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_87), .B(n_149), .Y(n_162) );
AND2x2_ASAP7_75t_L g197 ( .A(n_88), .B(n_125), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_90), .B(n_147), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_91), .A2(n_140), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_92), .B(n_149), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_93), .A2(n_140), .B(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_95), .B(n_147), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_96), .B(n_147), .Y(n_146) );
BUFx2_ASAP7_75t_L g470 ( .A(n_97), .Y(n_470) );
BUFx2_ASAP7_75t_L g763 ( .A(n_98), .Y(n_763) );
BUFx2_ASAP7_75t_SL g789 ( .A(n_98), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_99), .A2(n_140), .B(n_172), .Y(n_171) );
OAI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_105), .B(n_746), .Y(n_101) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_102), .A2(n_747), .B(n_751), .Y(n_746) );
INVxp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI22xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_116), .B1(n_433), .B2(n_742), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g750 ( .A(n_108), .Y(n_750) );
CKINVDCx11_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
OR2x6_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x6_ASAP7_75t_SL g745 ( .A(n_110), .B(n_112), .Y(n_745) );
OR2x2_ASAP7_75t_L g754 ( .A(n_110), .B(n_112), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_110), .B(n_111), .Y(n_765) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx3_ASAP7_75t_L g749 ( .A(n_116), .Y(n_749) );
AND2x4_ASAP7_75t_L g116 ( .A(n_117), .B(n_342), .Y(n_116) );
NOR4xp25_ASAP7_75t_L g117 ( .A(n_118), .B(n_260), .C(n_286), .D(n_326), .Y(n_117) );
OAI211xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_175), .B(n_206), .C(n_246), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_154), .Y(n_120) );
AND2x2_ASAP7_75t_L g413 ( .A(n_121), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_122), .B(n_154), .Y(n_280) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g207 ( .A(n_123), .B(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_123), .B(n_233), .Y(n_232) );
INVx5_ASAP7_75t_L g266 ( .A(n_123), .Y(n_266) );
NOR2x1_ASAP7_75t_SL g308 ( .A(n_123), .B(n_155), .Y(n_308) );
AND2x2_ASAP7_75t_L g364 ( .A(n_123), .B(n_167), .Y(n_364) );
OR2x6_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
INVx3_ASAP7_75t_L g196 ( .A(n_125), .Y(n_196) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AO21x2_ASAP7_75t_L g485 ( .A1(n_126), .A2(n_486), .B(n_492), .Y(n_485) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
BUFx4f_ASAP7_75t_L g168 ( .A(n_127), .Y(n_168) );
AND2x2_ASAP7_75t_SL g152 ( .A(n_128), .B(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g157 ( .A(n_128), .B(n_153), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_139), .B(n_151), .Y(n_129) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
AND2x6_ASAP7_75t_L g149 ( .A(n_133), .B(n_142), .Y(n_149) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x4_ASAP7_75t_L g147 ( .A(n_135), .B(n_144), .Y(n_147) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx5_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
AND2x2_ASAP7_75t_L g143 ( .A(n_138), .B(n_144), .Y(n_143) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_138), .Y(n_503) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx3_ASAP7_75t_L g504 ( .A(n_141), .Y(n_504) );
INVx2_ASAP7_75t_L g510 ( .A(n_142), .Y(n_510) );
AND2x4_ASAP7_75t_L g506 ( .A(n_143), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g502 ( .A(n_144), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_148), .B(n_150), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_149), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_150), .A2(n_161), .B(n_162), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_150), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_150), .A2(n_184), .B(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_150), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_150), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_150), .A2(n_212), .B(n_213), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_150), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_150), .A2(n_444), .B(n_445), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g449 ( .A1(n_150), .A2(n_450), .B(n_451), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_150), .A2(n_461), .B(n_462), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_150), .A2(n_468), .B(n_469), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_150), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_150), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_150), .A2(n_530), .B(n_531), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_151), .Y(n_215) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_151), .A2(n_220), .B(n_224), .Y(n_219) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_151), .A2(n_220), .B(n_224), .Y(n_259) );
AO21x2_ASAP7_75t_L g498 ( .A1(n_151), .A2(n_499), .B(n_505), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_151), .A2(n_527), .B(n_528), .Y(n_526) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_166), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_155), .B(n_167), .Y(n_236) );
AND2x2_ASAP7_75t_L g297 ( .A(n_155), .B(n_266), .Y(n_297) );
AO21x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_164), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_156), .B(n_165), .Y(n_164) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_156), .A2(n_158), .B(n_164), .Y(n_250) );
INVx1_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_157), .A2(n_170), .B(n_171), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_157), .B(n_187), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_157), .A2(n_441), .B(n_442), .Y(n_440) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_157), .A2(n_458), .B(n_459), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_163), .Y(n_158) );
AND2x2_ASAP7_75t_L g309 ( .A(n_166), .B(n_233), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_166), .B(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g353 ( .A(n_166), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g386 ( .A(n_166), .B(n_207), .Y(n_386) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g230 ( .A(n_167), .Y(n_230) );
AND2x2_ASAP7_75t_L g263 ( .A(n_167), .B(n_264), .Y(n_263) );
BUFx3_ASAP7_75t_L g298 ( .A(n_167), .Y(n_298) );
OR2x2_ASAP7_75t_L g374 ( .A(n_167), .B(n_233), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_168), .A2(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_SL g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_188), .Y(n_176) );
AOI211x1_ASAP7_75t_SL g303 ( .A1(n_177), .A2(n_295), .B(n_304), .C(n_306), .Y(n_303) );
AND2x2_ASAP7_75t_SL g348 ( .A(n_177), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_177), .B(n_346), .Y(n_393) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g218 ( .A(n_179), .Y(n_218) );
OAI21x1_ASAP7_75t_SL g179 ( .A1(n_180), .A2(n_182), .B(n_186), .Y(n_179) );
INVx1_ASAP7_75t_L g187 ( .A(n_181), .Y(n_187) );
AOI322xp5_ASAP7_75t_L g206 ( .A1(n_188), .A2(n_207), .A3(n_217), .B1(n_225), .B2(n_228), .C1(n_234), .C2(n_237), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_188), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_198), .Y(n_188) );
INVx2_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
INVxp67_ASAP7_75t_L g283 ( .A(n_189), .Y(n_283) );
BUFx3_ASAP7_75t_L g347 ( .A(n_189), .Y(n_347) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_196), .B(n_197), .Y(n_189) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_190), .A2(n_196), .B(n_197), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_195), .Y(n_190) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_196), .A2(n_199), .B(n_205), .Y(n_198) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_196), .A2(n_199), .B(n_205), .Y(n_245) );
AO21x1_ASAP7_75t_SL g446 ( .A1(n_196), .A2(n_447), .B(n_453), .Y(n_446) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_196), .A2(n_447), .B(n_453), .Y(n_522) );
INVx2_ASAP7_75t_L g256 ( .A(n_198), .Y(n_256) );
AND2x2_ASAP7_75t_L g305 ( .A(n_198), .B(n_219), .Y(n_305) );
AND2x2_ASAP7_75t_L g349 ( .A(n_198), .B(n_258), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_200), .B(n_204), .Y(n_199) );
AND2x2_ASAP7_75t_L g234 ( .A(n_207), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_207), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_SL g428 ( .A(n_207), .B(n_263), .Y(n_428) );
INVx4_ASAP7_75t_L g233 ( .A(n_208), .Y(n_233) );
AND2x2_ASAP7_75t_L g265 ( .A(n_208), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_208), .Y(n_318) );
AO21x2_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_215), .B(n_216), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_214), .Y(n_209) );
AOI21x1_ASAP7_75t_L g477 ( .A1(n_215), .A2(n_478), .B(n_484), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_217), .B(n_302), .Y(n_327) );
INVx1_ASAP7_75t_SL g366 ( .A(n_217), .Y(n_366) );
AND2x4_ASAP7_75t_L g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x4_ASAP7_75t_L g257 ( .A(n_218), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_218), .B(n_256), .Y(n_325) );
AND2x2_ASAP7_75t_L g377 ( .A(n_218), .B(n_227), .Y(n_377) );
OR2x2_ASAP7_75t_L g401 ( .A(n_218), .B(n_219), .Y(n_401) );
AND2x2_ASAP7_75t_L g225 ( .A(n_219), .B(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g275 ( .A(n_219), .B(n_256), .Y(n_275) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_219), .B(n_243), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_225), .B(n_338), .Y(n_355) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx2_ASAP7_75t_L g290 ( .A(n_227), .Y(n_290) );
AND2x4_ASAP7_75t_SL g330 ( .A(n_227), .B(n_244), .Y(n_330) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
OR2x2_ASAP7_75t_L g278 ( .A(n_229), .B(n_232), .Y(n_278) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g247 ( .A(n_230), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g395 ( .A(n_230), .B(n_308), .Y(n_395) );
AND2x2_ASAP7_75t_L g411 ( .A(n_230), .B(n_265), .Y(n_411) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AOI311xp33_ASAP7_75t_L g381 ( .A1(n_232), .A2(n_320), .A3(n_382), .B(n_384), .C(n_391), .Y(n_381) );
AND2x4_ASAP7_75t_L g248 ( .A(n_233), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g252 ( .A(n_233), .Y(n_252) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_233), .B(n_266), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_233), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g365 ( .A(n_233), .B(n_352), .Y(n_365) );
AND2x2_ASAP7_75t_L g251 ( .A(n_235), .B(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_236), .Y(n_269) );
OR2x2_ASAP7_75t_L g358 ( .A(n_236), .B(n_322), .Y(n_358) );
INVx1_ASAP7_75t_L g414 ( .A(n_236), .Y(n_414) );
INVx1_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_242), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g323 ( .A(n_240), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g337 ( .A(n_240), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g412 ( .A(n_240), .B(n_285), .Y(n_412) );
BUFx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
AND2x2_ASAP7_75t_L g255 ( .A(n_241), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g274 ( .A(n_241), .B(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g336 ( .A(n_242), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_242), .A2(n_392), .B1(n_393), .B2(n_394), .Y(n_391) );
OR2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g285 ( .A(n_243), .B(n_256), .Y(n_285) );
AND2x4_ASAP7_75t_L g338 ( .A(n_243), .B(n_245), .Y(n_338) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
OAI21xp33_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_251), .B(n_253), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_247), .A2(n_333), .B1(n_337), .B2(n_339), .Y(n_332) );
AND2x2_ASAP7_75t_SL g292 ( .A(n_248), .B(n_266), .Y(n_292) );
INVx2_ASAP7_75t_L g354 ( .A(n_248), .Y(n_354) );
AND2x2_ASAP7_75t_L g368 ( .A(n_248), .B(n_364), .Y(n_368) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g264 ( .A(n_250), .Y(n_264) );
INVx1_ASAP7_75t_L g317 ( .A(n_250), .Y(n_317) );
INVx1_ASAP7_75t_L g268 ( .A(n_252), .Y(n_268) );
AND3x2_ASAP7_75t_L g296 ( .A(n_252), .B(n_297), .C(n_298), .Y(n_296) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g360 ( .A(n_255), .Y(n_360) );
AND2x2_ASAP7_75t_L g288 ( .A(n_257), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g359 ( .A(n_257), .B(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_257), .A2(n_371), .B1(n_375), .B2(n_378), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_257), .B(n_405), .Y(n_409) );
BUFx2_ASAP7_75t_L g300 ( .A(n_258), .Y(n_300) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g271 ( .A(n_259), .Y(n_271) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_259), .Y(n_390) );
OAI221xp5_ASAP7_75t_SL g260 ( .A1(n_261), .A2(n_270), .B1(n_272), .B2(n_273), .C(n_276), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
INVx1_ASAP7_75t_L g352 ( .A(n_264), .Y(n_352) );
INVx2_ASAP7_75t_SL g341 ( .A(n_265), .Y(n_341) );
AND2x2_ASAP7_75t_L g423 ( .A(n_265), .B(n_290), .Y(n_423) );
INVx4_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
INVx1_ASAP7_75t_L g272 ( .A(n_267), .Y(n_272) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
AND2x4_ASAP7_75t_L g383 ( .A(n_271), .B(n_338), .Y(n_383) );
INVx1_ASAP7_75t_SL g422 ( .A(n_271), .Y(n_422) );
AND2x2_ASAP7_75t_L g427 ( .A(n_271), .B(n_330), .Y(n_427) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g369 ( .A(n_275), .Y(n_369) );
OAI21xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_279), .B(n_281), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g302 ( .A(n_283), .Y(n_302) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g299 ( .A(n_285), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g389 ( .A(n_285), .B(n_390), .Y(n_389) );
OAI211xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_291), .B(n_293), .C(n_310), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g382 ( .A(n_289), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_290), .B(n_305), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_290), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g415 ( .A(n_290), .B(n_338), .Y(n_415) );
OAI221xp5_ASAP7_75t_SL g326 ( .A1(n_291), .A2(n_315), .B1(n_327), .B2(n_328), .C(n_332), .Y(n_326) );
INVx3_ASAP7_75t_SL g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g397 ( .A(n_292), .B(n_298), .Y(n_397) );
OAI32xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .A3(n_301), .B1(n_303), .B2(n_307), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVxp67_ASAP7_75t_SL g387 ( .A(n_297), .Y(n_387) );
INVx2_ASAP7_75t_L g320 ( .A(n_298), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g429 ( .A1(n_298), .A2(n_350), .B(n_430), .C(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g335 ( .A(n_300), .Y(n_335) );
OR2x2_ASAP7_75t_L g431 ( .A(n_300), .B(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_304), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g392 ( .A(n_307), .Y(n_392) );
AND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_L g373 ( .A(n_308), .Y(n_373) );
OAI21xp33_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_319), .B(n_323), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
OR2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_314), .B(n_317), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_316), .A2(n_348), .B1(n_417), .B2(n_420), .C(n_424), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_316), .Y(n_419) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
OR2x2_ASAP7_75t_L g340 ( .A(n_320), .B(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g407 ( .A(n_320), .B(n_365), .Y(n_407) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g405 ( .A(n_330), .Y(n_405) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_338), .B(n_368), .Y(n_425) );
INVx2_ASAP7_75t_L g432 ( .A(n_338), .Y(n_432) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_340), .A2(n_403), .B1(n_406), .B2(n_408), .C(n_410), .Y(n_402) );
AND5x1_ASAP7_75t_L g342 ( .A(n_343), .B(n_381), .C(n_396), .D(n_416), .E(n_426), .Y(n_342) );
NOR2xp33_ASAP7_75t_SL g343 ( .A(n_344), .B(n_361), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_350), .B1(n_353), .B2(n_355), .C(n_356), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI221xp5_ASAP7_75t_SL g361 ( .A1(n_362), .A2(n_366), .B1(n_367), .B2(n_369), .C(n_370), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_366), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
OR2x2_ASAP7_75t_L g379 ( .A(n_374), .B(n_380), .Y(n_379) );
CKINVDCx16_ASAP7_75t_R g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B(n_388), .Y(n_384) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_402), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_413), .B2(n_415), .Y(n_410) );
O2A1O1Ixp33_ASAP7_75t_L g426 ( .A1(n_412), .A2(n_427), .B(n_428), .C(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g430 ( .A(n_423), .Y(n_430) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx4_ASAP7_75t_L g748 ( .A(n_433), .Y(n_748) );
OAI22xp5_ASAP7_75t_SL g768 ( .A1(n_433), .A2(n_748), .B1(n_769), .B2(n_770), .Y(n_768) );
AND3x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_620), .C(n_716), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_562), .C(n_589), .Y(n_434) );
OAI211xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_472), .B(n_511), .C(n_535), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_454), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_437), .A2(n_513), .B(n_517), .C(n_523), .Y(n_512) );
OR2x2_ASAP7_75t_L g635 ( .A(n_437), .B(n_572), .Y(n_635) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g602 ( .A(n_438), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_438), .B(n_573), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_438), .B(n_718), .Y(n_733) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_446), .Y(n_438) );
AND2x2_ASAP7_75t_L g519 ( .A(n_439), .B(n_455), .Y(n_519) );
INVx1_ASAP7_75t_L g539 ( .A(n_439), .Y(n_539) );
OR2x2_ASAP7_75t_L g554 ( .A(n_439), .B(n_463), .Y(n_554) );
INVx2_ASAP7_75t_L g560 ( .A(n_439), .Y(n_560) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_439), .Y(n_615) );
INVx1_ASAP7_75t_L g692 ( .A(n_439), .Y(n_692) );
NOR2x1_ASAP7_75t_SL g541 ( .A(n_446), .B(n_463), .Y(n_541) );
AND2x2_ASAP7_75t_L g571 ( .A(n_446), .B(n_560), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_452), .Y(n_447) );
OR2x2_ASAP7_75t_L g565 ( .A(n_454), .B(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_454), .B(n_672), .Y(n_671) );
INVx3_ASAP7_75t_L g693 ( .A(n_454), .Y(n_693) );
NAND2x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_463), .Y(n_454) );
OR2x2_ASAP7_75t_SL g553 ( .A(n_455), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g557 ( .A(n_455), .Y(n_557) );
INVx4_ASAP7_75t_L g573 ( .A(n_455), .Y(n_573) );
OR2x2_ASAP7_75t_L g588 ( .A(n_455), .B(n_521), .Y(n_588) );
AND2x2_ASAP7_75t_L g627 ( .A(n_455), .B(n_541), .Y(n_627) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_455), .Y(n_639) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
AND2x2_ASAP7_75t_L g520 ( .A(n_463), .B(n_521), .Y(n_520) );
OR2x2_ASAP7_75t_L g572 ( .A(n_463), .B(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_L g587 ( .A(n_463), .Y(n_587) );
AND2x2_ASAP7_75t_L g603 ( .A(n_463), .B(n_573), .Y(n_603) );
AND2x2_ASAP7_75t_L g616 ( .A(n_463), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g648 ( .A(n_463), .B(n_560), .Y(n_648) );
INVx2_ASAP7_75t_SL g718 ( .A(n_463), .Y(n_718) );
OR2x6_ASAP7_75t_L g463 ( .A(n_464), .B(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_474), .B(n_493), .Y(n_473) );
OAI211xp5_ASAP7_75t_L g589 ( .A1(n_474), .A2(n_590), .B(n_594), .C(n_610), .Y(n_589) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g685 ( .A(n_475), .B(n_524), .Y(n_685) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_485), .Y(n_475) );
INVx2_ASAP7_75t_L g534 ( .A(n_476), .Y(n_534) );
AND2x4_ASAP7_75t_SL g545 ( .A(n_476), .B(n_525), .Y(n_545) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_476), .Y(n_549) );
AND2x2_ASAP7_75t_L g607 ( .A(n_476), .B(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g681 ( .A(n_476), .Y(n_681) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_477), .Y(n_583) );
AND2x2_ASAP7_75t_L g626 ( .A(n_477), .B(n_485), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_483), .Y(n_478) );
INVx2_ASAP7_75t_L g516 ( .A(n_485), .Y(n_516) );
AND2x2_ASAP7_75t_L g576 ( .A(n_485), .B(n_525), .Y(n_576) );
INVx2_ASAP7_75t_L g608 ( .A(n_485), .Y(n_608) );
OR2x2_ASAP7_75t_L g631 ( .A(n_485), .B(n_496), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_493), .B(n_548), .Y(n_655) );
AND2x2_ASAP7_75t_L g689 ( .A(n_493), .B(n_625), .Y(n_689) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
OAI31xp33_ASAP7_75t_SL g610 ( .A1(n_494), .A2(n_591), .A3(n_611), .B(n_618), .Y(n_610) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_495), .B(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
AND2x2_ASAP7_75t_L g561 ( .A(n_496), .B(n_524), .Y(n_561) );
AND2x4_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AND2x4_ASAP7_75t_L g551 ( .A(n_497), .B(n_498), .Y(n_551) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
NOR2x1p5_ASAP7_75t_L g507 ( .A(n_508), .B(n_509), .Y(n_507) );
INVx3_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g696 ( .A(n_514), .Y(n_696) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_516), .B(n_525), .Y(n_578) );
AND2x2_ASAP7_75t_L g619 ( .A(n_516), .B(n_534), .Y(n_619) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
AND2x2_ASAP7_75t_L g599 ( .A(n_520), .B(n_557), .Y(n_599) );
AND2x2_ASAP7_75t_L g558 ( .A(n_521), .B(n_559), .Y(n_558) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_521), .Y(n_567) );
INVx2_ASAP7_75t_L g617 ( .A(n_521), .Y(n_617) );
AND2x2_ASAP7_75t_L g707 ( .A(n_521), .B(n_692), .Y(n_707) );
INVx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g713 ( .A(n_523), .Y(n_713) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_524), .B(n_533), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_524), .B(n_583), .Y(n_652) );
AND2x2_ASAP7_75t_L g700 ( .A(n_524), .B(n_626), .Y(n_700) );
INVx4_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g609 ( .A(n_525), .B(n_581), .Y(n_609) );
AND2x2_ASAP7_75t_L g618 ( .A(n_525), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g630 ( .A(n_525), .Y(n_630) );
BUFx2_ASAP7_75t_L g646 ( .A(n_525), .Y(n_646) );
AND2x4_ASAP7_75t_L g680 ( .A(n_525), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g725 ( .A(n_525), .B(n_626), .Y(n_725) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_532), .Y(n_525) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AOI222xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_542), .B1(n_546), .B2(n_552), .C1(n_555), .C2(n_561), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_537), .A2(n_601), .B1(n_604), .B2(n_609), .Y(n_600) );
OR2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
AND2x2_ASAP7_75t_L g584 ( .A(n_538), .B(n_585), .Y(n_584) );
AND2x4_ASAP7_75t_SL g598 ( .A(n_538), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_538), .B(n_603), .Y(n_736) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g697 ( .A(n_539), .B(n_603), .Y(n_697) );
OR2x2_ASAP7_75t_L g674 ( .A(n_540), .B(n_556), .Y(n_674) );
OR2x2_ASAP7_75t_L g682 ( .A(n_540), .B(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g666 ( .A(n_541), .B(n_559), .Y(n_666) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OR2x2_ASAP7_75t_L g574 ( .A(n_544), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g724 ( .A(n_544), .B(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g675 ( .A(n_545), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_545), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_SL g710 ( .A(n_545), .Y(n_710) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
INVx2_ASAP7_75t_L g695 ( .A(n_548), .Y(n_695) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g597 ( .A(n_549), .B(n_576), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_550), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g596 ( .A(n_550), .Y(n_596) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_550), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g699 ( .A(n_550), .B(n_571), .Y(n_699) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g633 ( .A(n_551), .B(n_619), .Y(n_633) );
AND2x2_ASAP7_75t_L g676 ( .A(n_551), .B(n_608), .Y(n_676) );
AND2x4_ASAP7_75t_L g591 ( .A(n_552), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g732 ( .A(n_554), .B(n_588), .Y(n_732) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_556), .B(n_571), .Y(n_715) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_557), .B(n_571), .Y(n_637) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_557), .A2(n_598), .B(n_699), .C(n_700), .Y(n_698) );
AND2x2_ASAP7_75t_L g729 ( .A(n_557), .B(n_707), .Y(n_729) );
INVx1_ASAP7_75t_L g640 ( .A(n_558), .Y(n_640) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_561), .B(n_625), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_574), .B(n_577), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_565), .A2(n_718), .B1(n_719), .B2(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g593 ( .A(n_567), .Y(n_593) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NOR2xp67_ASAP7_75t_L g614 ( .A(n_573), .B(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g665 ( .A(n_573), .Y(n_665) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_579), .B(n_584), .Y(n_577) );
INVx1_ASAP7_75t_L g656 ( .A(n_578), .Y(n_656) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_598), .B(n_600), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
OR2x2_ASAP7_75t_L g641 ( .A(n_596), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g678 ( .A(n_596), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_596), .B(n_626), .Y(n_714) );
INVx1_ASAP7_75t_L g734 ( .A(n_597), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_599), .A2(n_702), .B1(n_705), .B2(n_708), .C(n_711), .Y(n_701) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI321xp33_ASAP7_75t_L g722 ( .A1(n_604), .A2(n_639), .A3(n_723), .B1(n_726), .B2(n_728), .C(n_730), .Y(n_722) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g663 ( .A(n_608), .Y(n_663) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g657 ( .A(n_613), .Y(n_657) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx1_ASAP7_75t_L g683 ( .A(n_614), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_616), .A2(n_644), .B1(n_648), .B2(n_649), .C(n_654), .Y(n_643) );
INVxp67_ASAP7_75t_L g672 ( .A(n_617), .Y(n_672) );
INVx1_ASAP7_75t_L g642 ( .A(n_619), .Y(n_642) );
NOR2xp67_ASAP7_75t_L g620 ( .A(n_621), .B(n_667), .Y(n_620) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_643), .C(n_658), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_627), .B1(n_628), .B2(n_634), .C(n_636), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g741 ( .A(n_626), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_629), .B(n_632), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g721 ( .A(n_630), .B(n_676), .Y(n_721) );
INVx2_ASAP7_75t_SL g653 ( .A(n_631), .Y(n_653) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_632), .A2(n_637), .B1(n_638), .B2(n_641), .Y(n_636) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
HB1xp67_ASAP7_75t_L g727 ( .A(n_640), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_641), .B(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g647 ( .A(n_642), .Y(n_647) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_644), .A2(n_687), .B1(n_689), .B2(n_690), .C1(n_694), .C2(n_697), .Y(n_686) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_645), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g720 ( .A(n_645), .B(n_699), .Y(n_720) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_651), .B(n_653), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_653), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_653), .B(n_713), .Y(n_712) );
AOI21xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B(n_657), .Y(n_654) );
NAND2xp33_ASAP7_75t_SL g658 ( .A(n_659), .B(n_664), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_664), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND4xp25_ASAP7_75t_SL g667 ( .A(n_668), .B(n_686), .C(n_698), .D(n_701), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_673), .B(n_675), .C(n_677), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_674), .A2(n_678), .B1(n_682), .B2(n_684), .Y(n_677) );
INVx1_ASAP7_75t_L g704 ( .A(n_676), .Y(n_704) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_693), .Y(n_690) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_693), .B(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_710), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_715), .Y(n_711) );
NOR4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_722), .C(n_735), .D(n_737), .Y(n_716) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
HB1xp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx4_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx3_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
OAI22x1_ASAP7_75t_L g747 ( .A1(n_744), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
BUFx2_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AND2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_764), .Y(n_757) );
INVxp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_760), .B(n_763), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OR2x2_ASAP7_75t_SL g784 ( .A(n_761), .B(n_763), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_761), .A2(n_787), .B(n_790), .Y(n_786) );
INVx1_ASAP7_75t_SL g774 ( .A(n_764), .Y(n_774) );
BUFx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
BUFx3_ASAP7_75t_L g779 ( .A(n_765), .Y(n_779) );
BUFx2_ASAP7_75t_L g791 ( .A(n_765), .Y(n_791) );
INVxp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_773), .B(n_775), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx1_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
NOR2xp33_ASAP7_75t_SL g775 ( .A(n_776), .B(n_780), .Y(n_775) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
BUFx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_779), .Y(n_778) );
CKINVDCx9p33_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
CKINVDCx11_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx8_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
endmodule