module fake_jpeg_18635_n_159 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_159);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_159;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

INVx11_ASAP7_75t_SL g67 ( 
.A(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_7),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_40),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_69),
.Y(n_96)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_85),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_74),
.Y(n_92)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_50),
.B1(n_77),
.B2(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_93),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_54),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_73),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_75),
.B1(n_63),
.B2(n_65),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_94),
.A2(n_60),
.B1(n_62),
.B2(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_57),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_76),
.B1(n_60),
.B2(n_53),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_66),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_68),
.C(n_59),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_80),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_70),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_125),
.B(n_3),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_48),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_120),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_108),
.A2(n_51),
.B1(n_77),
.B2(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_122),
.B1(n_0),
.B2(n_2),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_126),
.C(n_28),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_106),
.B(n_71),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_123),
.B(n_5),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_80),
.B1(n_79),
.B2(n_84),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_105),
.A2(n_56),
.B1(n_55),
.B2(n_72),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_108),
.A2(n_79),
.B1(n_61),
.B2(n_21),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_106),
.B(n_20),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_13),
.C(n_44),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_127),
.B(n_131),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_116),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_26),
.C(n_43),
.Y(n_132)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_125),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_145),
.B(n_146),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_142),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_140),
.A2(n_112),
.B(n_128),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_147),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_144),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_150),
.B(n_144),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_151),
.A2(n_143),
.B1(n_128),
.B2(n_139),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_143),
.A3(n_114),
.B1(n_137),
.B2(n_141),
.C1(n_134),
.C2(n_115),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_136),
.B(n_141),
.C(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_155),
.A2(n_30),
.B(n_31),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_156),
.Y(n_157)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_33),
.B(n_37),
.Y(n_158)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_158),
.Y(n_159)
);


endmodule