module fake_jpeg_15487_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_96;

INVxp33_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_79),
.Y(n_87)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_56),
.B1(n_51),
.B2(n_72),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_57),
.B1(n_55),
.B2(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_68),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_47),
.B(n_63),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_54),
.B1(n_60),
.B2(n_48),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_56),
.B1(n_70),
.B2(n_58),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_70),
.B1(n_47),
.B2(n_67),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_94),
.Y(n_111)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_101),
.B1(n_104),
.B2(n_107),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_106),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_63),
.B1(n_53),
.B2(n_50),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_80),
.A2(n_53),
.B1(n_66),
.B2(n_52),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_93),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_112),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_85),
.B1(n_89),
.B2(n_97),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_109),
.Y(n_124)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_71),
.B1(n_65),
.B2(n_3),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_62),
.B1(n_49),
.B2(n_55),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_85),
.A2(n_20),
.B1(n_43),
.B2(n_41),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_85),
.A2(n_17),
.B1(n_39),
.B2(n_38),
.Y(n_119)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_0),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_127),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_132),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_98),
.B(n_104),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_140),
.B(n_122),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_101),
.B(n_100),
.C(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_118),
.B1(n_102),
.B2(n_113),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_141),
.A2(n_134),
.B1(n_128),
.B2(n_129),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_142),
.A2(n_144),
.B(n_145),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_141),
.B1(n_131),
.B2(n_137),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_125),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_131),
.B(n_103),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_146),
.A2(n_133),
.B(n_5),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_124),
.B1(n_139),
.B2(n_131),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_147),
.A2(n_149),
.B1(n_4),
.B2(n_5),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_138),
.B1(n_124),
.B2(n_111),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_4),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_153),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_23),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_150),
.CI(n_154),
.CON(n_158),
.SN(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_155),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_161),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_19),
.C(n_36),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_16),
.B(n_35),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_13),
.Y(n_166)
);

OAI321xp33_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_22),
.A3(n_31),
.B1(n_30),
.B2(n_29),
.C(n_27),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_11),
.B(n_26),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_44),
.C(n_25),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_24),
.Y(n_170)
);


endmodule