module fake_netlist_1_178_n_1086 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_225, n_39, n_1086);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1086;
wire n_663;
wire n_707;
wire n_791;
wire n_513;
wire n_361;
wire n_963;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_564;
wire n_353;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_975;
wire n_1042;
wire n_1060;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_937;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1025;
wire n_1011;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_771;
wire n_735;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_950;
wire n_427;
wire n_910;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_423;
wire n_420;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_1050;
wire n_370;
wire n_1058;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_899;
wire n_881;
wire n_806;
wire n_539;
wire n_1055;
wire n_1066;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_955;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_924;
wire n_912;
wire n_947;
wire n_1043;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1040;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
wire n_269;
INVx1_ASAP7_75t_L g266 ( .A(n_136), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_219), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_62), .Y(n_268) );
CKINVDCx14_ASAP7_75t_R g269 ( .A(n_197), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_53), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_211), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_166), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_142), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_259), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_141), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_143), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_174), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_125), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_84), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_50), .Y(n_280) );
BUFx2_ASAP7_75t_SL g281 ( .A(n_244), .Y(n_281) );
NOR2xp67_ASAP7_75t_L g282 ( .A(n_171), .B(n_231), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_189), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_217), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_193), .Y(n_285) );
CKINVDCx20_ASAP7_75t_R g286 ( .A(n_69), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_185), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_100), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_165), .Y(n_289) );
INVxp67_ASAP7_75t_L g290 ( .A(n_86), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_49), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_123), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_40), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_223), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_134), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_264), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_220), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_225), .Y(n_299) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_28), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_230), .Y(n_301) );
NOR2xp67_ASAP7_75t_L g302 ( .A(n_260), .B(n_168), .Y(n_302) );
CKINVDCx14_ASAP7_75t_R g303 ( .A(n_49), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_10), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_216), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_94), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g307 ( .A(n_48), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_24), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_154), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_18), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_239), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_51), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_35), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_215), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_252), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g316 ( .A(n_66), .Y(n_316) );
INVxp33_ASAP7_75t_L g317 ( .A(n_117), .Y(n_317) );
BUFx8_ASAP7_75t_SL g318 ( .A(n_4), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_241), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_32), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_21), .B(n_172), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_206), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_173), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_258), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_218), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_21), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_38), .Y(n_327) );
CKINVDCx16_ASAP7_75t_R g328 ( .A(n_176), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_59), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_192), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_207), .Y(n_331) );
INVx2_ASAP7_75t_SL g332 ( .A(n_203), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_13), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_194), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_118), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_78), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_127), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_163), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_233), .Y(n_339) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_65), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_153), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_235), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_175), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_157), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_181), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_243), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_29), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_145), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_135), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_257), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_164), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_139), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_238), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_101), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_248), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_29), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_95), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_74), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_263), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_242), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_1), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_209), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_47), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_101), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_167), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_72), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_195), .Y(n_367) );
CKINVDCx16_ASAP7_75t_R g368 ( .A(n_214), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_191), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_85), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_131), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_104), .Y(n_372) );
CKINVDCx14_ASAP7_75t_R g373 ( .A(n_234), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_76), .Y(n_374) );
INVxp33_ASAP7_75t_L g375 ( .A(n_169), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_13), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_170), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_45), .Y(n_378) );
BUFx2_ASAP7_75t_L g379 ( .A(n_202), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_232), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_158), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_254), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_208), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_129), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_137), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_57), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_196), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_183), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_16), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_67), .Y(n_390) );
BUFx2_ASAP7_75t_L g391 ( .A(n_261), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_47), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_245), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_224), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_109), .Y(n_395) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_14), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_59), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_182), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_55), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_148), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_71), .Y(n_401) );
CKINVDCx16_ASAP7_75t_R g402 ( .A(n_0), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g403 ( .A(n_204), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_184), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_200), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_186), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_222), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_57), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_308), .B(n_0), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_407), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_305), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_379), .B(n_1), .Y(n_412) );
INVx3_ASAP7_75t_L g413 ( .A(n_407), .Y(n_413) );
INVx5_ASAP7_75t_L g414 ( .A(n_407), .Y(n_414) );
OAI22xp5_ASAP7_75t_SL g415 ( .A1(n_286), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_278), .Y(n_416) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_355), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_305), .Y(n_418) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_355), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_278), .Y(n_420) );
INVx4_ASAP7_75t_L g421 ( .A(n_379), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_391), .B(n_5), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_289), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_289), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_308), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_309), .A2(n_311), .B(n_297), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_294), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_309), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_393), .Y(n_429) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_393), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_391), .B(n_6), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_303), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_371), .B(n_9), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_311), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_294), .Y(n_435) );
CKINVDCx8_ASAP7_75t_R g436 ( .A(n_328), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_297), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_313), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_313), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_329), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_298), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_382), .B(n_10), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_318), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_317), .B(n_11), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_310), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_310), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_320), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_298), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_332), .B(n_11), .Y(n_449) );
AND2x6_ASAP7_75t_L g450 ( .A(n_321), .B(n_116), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_318), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_421), .B(n_320), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_421), .B(n_326), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_435), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_425), .A2(n_288), .B1(n_402), .B2(n_366), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_443), .Y(n_456) );
XOR2xp5_ASAP7_75t_L g457 ( .A(n_451), .B(n_300), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_451), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_421), .B(n_368), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_435), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_421), .B(n_375), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_435), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_414), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_443), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_435), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_445), .B(n_326), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_435), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_445), .B(n_307), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_435), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_445), .B(n_307), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_414), .Y(n_472) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_435), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_422), .B(n_321), .Y(n_474) );
NAND2xp33_ASAP7_75t_SL g475 ( .A(n_444), .B(n_285), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_409), .A2(n_396), .B1(n_319), .B2(n_334), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_422), .B(n_395), .Y(n_477) );
BUFx4f_ASAP7_75t_L g478 ( .A(n_450), .Y(n_478) );
BUFx10_ASAP7_75t_L g479 ( .A(n_422), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_409), .A2(n_422), .B1(n_431), .B2(n_432), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_417), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_413), .B(n_316), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_414), .Y(n_483) );
OAI22xp5_ASAP7_75t_SL g484 ( .A1(n_415), .A2(n_300), .B1(n_401), .B2(n_340), .Y(n_484) );
BUFx10_ASAP7_75t_L g485 ( .A(n_422), .Y(n_485) );
INVx4_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_450), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_431), .A2(n_306), .B1(n_312), .B2(n_304), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_446), .Y(n_489) );
INVx2_ASAP7_75t_SL g490 ( .A(n_414), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_431), .B(n_271), .Y(n_491) );
OR2x6_ASAP7_75t_L g492 ( .A(n_431), .B(n_281), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_414), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_417), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_461), .B(n_444), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_474), .A2(n_450), .B1(n_411), .B2(n_428), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_452), .B(n_431), .Y(n_497) );
NOR2x1p5_ASAP7_75t_L g498 ( .A(n_456), .B(n_412), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_452), .B(n_412), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_452), .B(n_411), .Y(n_500) );
AND2x4_ASAP7_75t_L g501 ( .A(n_492), .B(n_433), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_452), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_453), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_489), .Y(n_505) );
INVx4_ASAP7_75t_L g506 ( .A(n_479), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_489), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_453), .B(n_418), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_453), .B(n_434), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_459), .B(n_434), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_466), .B(n_449), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_480), .A2(n_442), .B1(n_450), .B2(n_432), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_482), .B(n_413), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_454), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_477), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_468), .B(n_413), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_486), .B(n_414), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_486), .B(n_413), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_479), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_477), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_478), .A2(n_469), .B(n_463), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_471), .B(n_413), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_492), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_474), .B(n_436), .Y(n_524) );
AND2x6_ASAP7_75t_SL g525 ( .A(n_457), .B(n_442), .Y(n_525) );
OAI22xp33_ASAP7_75t_L g526 ( .A1(n_480), .A2(n_319), .B1(n_341), .B2(n_334), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_491), .A2(n_426), .B(n_410), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_458), .Y(n_528) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_479), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_492), .B(n_450), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_456), .Y(n_531) );
O2A1O1Ixp5_ASAP7_75t_L g532 ( .A1(n_478), .A2(n_446), .B(n_447), .C(n_410), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_488), .B(n_426), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_475), .A2(n_450), .B1(n_396), .B2(n_341), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_479), .B(n_426), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_485), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_487), .B(n_266), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_485), .B(n_446), .Y(n_538) );
INVx5_ASAP7_75t_L g539 ( .A(n_490), .Y(n_539) );
NAND3xp33_ASAP7_75t_SL g540 ( .A(n_464), .B(n_401), .C(n_340), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_485), .B(n_438), .Y(n_541) );
AND2x6_ASAP7_75t_L g542 ( .A(n_478), .B(n_410), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_476), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_487), .A2(n_450), .B1(n_416), .B2(n_423), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_454), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_455), .A2(n_416), .B(n_423), .C(n_420), .Y(n_546) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_484), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_472), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_472), .B(n_267), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_460), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_483), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_460), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_493), .B(n_439), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_462), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_465), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_484), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_462), .B(n_272), .Y(n_557) );
INVx8_ASAP7_75t_L g558 ( .A(n_462), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_481), .B(n_447), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_481), .B(n_447), .Y(n_560) );
INVx3_ASAP7_75t_L g561 ( .A(n_462), .Y(n_561) );
AND2x6_ASAP7_75t_SL g562 ( .A(n_462), .B(n_408), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_494), .B(n_271), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_470), .B(n_273), .Y(n_564) );
OR2x6_ASAP7_75t_L g565 ( .A(n_470), .B(n_281), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_470), .B(n_439), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_470), .B(n_275), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_465), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_467), .B(n_274), .Y(n_569) );
NAND2x1p5_ASAP7_75t_L g570 ( .A(n_506), .B(n_378), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_524), .B(n_327), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_535), .A2(n_467), .B(n_332), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_496), .A2(n_269), .B1(n_373), .B2(n_336), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_543), .B(n_333), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_504), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
BUFx4f_ASAP7_75t_L g577 ( .A(n_530), .Y(n_577) );
BUFx8_ASAP7_75t_L g578 ( .A(n_501), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_520), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_498), .B(n_268), .Y(n_580) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_546), .A2(n_290), .B(n_279), .C(n_280), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_519), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_511), .B(n_357), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_528), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_502), .Y(n_585) );
NOR3xp33_ASAP7_75t_SL g586 ( .A(n_526), .B(n_376), .C(n_370), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_519), .B(n_284), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_519), .B(n_284), .Y(n_588) );
O2A1O1Ixp33_ASAP7_75t_L g589 ( .A1(n_546), .A2(n_291), .B(n_293), .C(n_270), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_503), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_519), .B(n_287), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_540), .B(n_386), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_501), .A2(n_389), .B1(n_392), .B2(n_390), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_534), .A2(n_399), .B1(n_392), .B2(n_296), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_531), .B(n_399), .Y(n_595) );
NAND2xp33_ASAP7_75t_SL g596 ( .A(n_523), .B(n_287), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_499), .B(n_296), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_547), .B(n_556), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_500), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_510), .B(n_314), .Y(n_600) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_529), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_495), .B(n_347), .Y(n_602) );
CKINVDCx14_ASAP7_75t_R g603 ( .A(n_526), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_518), .A2(n_473), .B(n_277), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_508), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_509), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_541), .B(n_315), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_497), .A2(n_323), .B1(n_344), .B2(n_322), .Y(n_608) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_525), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_516), .A2(n_427), .B1(n_437), .B2(n_424), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_522), .B(n_440), .Y(n_611) );
BUFx3_ASAP7_75t_L g612 ( .A(n_539), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_529), .B(n_344), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_527), .A2(n_553), .B(n_533), .C(n_513), .Y(n_614) );
OAI21x1_ASAP7_75t_SL g615 ( .A1(n_544), .A2(n_337), .B(n_335), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_529), .B(n_346), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_536), .B(n_354), .Y(n_617) );
NOR2xp67_ASAP7_75t_L g618 ( .A(n_539), .B(n_437), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_553), .B(n_440), .Y(n_619) );
OR2x6_ASAP7_75t_L g620 ( .A(n_565), .B(n_329), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_551), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_544), .B(n_346), .Y(n_622) );
OAI22x1_ASAP7_75t_L g623 ( .A1(n_562), .A2(n_351), .B1(n_359), .B2(n_350), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_507), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_549), .Y(n_625) );
A2O1A1Ixp33_ASAP7_75t_L g626 ( .A1(n_532), .A2(n_448), .B(n_441), .C(n_358), .Y(n_626) );
INVx4_ASAP7_75t_L g627 ( .A(n_539), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_517), .A2(n_283), .B(n_276), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g629 ( .A1(n_537), .A2(n_361), .B(n_363), .C(n_356), .Y(n_629) );
OR2x6_ASAP7_75t_SL g630 ( .A(n_538), .B(n_365), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_537), .B(n_364), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_505), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_517), .A2(n_295), .B(n_292), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_521), .A2(n_301), .B(n_299), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_566), .A2(n_448), .B(n_441), .C(n_372), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_542), .A2(n_448), .B1(n_441), .B2(n_374), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_548), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_566), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_563), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_569), .A2(n_325), .B(n_324), .Y(n_641) );
AOI21x1_ASAP7_75t_L g642 ( .A1(n_557), .A2(n_302), .B(n_282), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_560), .A2(n_331), .B(n_330), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_558), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_557), .A2(n_387), .B1(n_403), .B2(n_385), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_542), .B(n_385), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_564), .A2(n_339), .B(n_338), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_564), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_567), .A2(n_403), .B1(n_387), .B2(n_397), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_567), .Y(n_650) );
OR2x6_ASAP7_75t_L g651 ( .A(n_558), .B(n_342), .Y(n_651) );
BUFx12f_ASAP7_75t_L g652 ( .A(n_554), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_514), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_568), .A2(n_343), .B(n_348), .C(n_345), .Y(n_654) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_545), .A2(n_352), .B(n_349), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_561), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_550), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_550), .Y(n_658) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_561), .Y(n_659) );
BUFx8_ASAP7_75t_L g660 ( .A(n_552), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_552), .A2(n_360), .B1(n_367), .B2(n_362), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_555), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_555), .B(n_12), .Y(n_663) );
BUFx12f_ASAP7_75t_L g664 ( .A(n_528), .Y(n_664) );
INVx3_ASAP7_75t_L g665 ( .A(n_506), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_524), .B(n_369), .Y(n_666) );
INVx3_ASAP7_75t_L g667 ( .A(n_506), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g668 ( .A(n_528), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_511), .B(n_377), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_512), .A2(n_380), .B1(n_383), .B2(n_381), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_511), .B(n_384), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_524), .B(n_388), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_511), .B(n_394), .Y(n_673) );
INVx8_ASAP7_75t_L g674 ( .A(n_519), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_504), .Y(n_675) );
AND2x4_ASAP7_75t_L g676 ( .A(n_506), .B(n_398), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_512), .A2(n_400), .B1(n_406), .B2(n_405), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_660), .Y(n_678) );
BUFx12f_ASAP7_75t_L g679 ( .A(n_660), .Y(n_679) );
CKINVDCx5p33_ASAP7_75t_R g680 ( .A(n_664), .Y(n_680) );
AO32x2_ASAP7_75t_L g681 ( .A1(n_573), .A2(n_430), .A3(n_429), .B1(n_419), .B2(n_417), .Y(n_681) );
OAI21xp33_ASAP7_75t_SL g682 ( .A1(n_670), .A2(n_404), .B(n_353), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_574), .B(n_12), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_603), .A2(n_430), .B1(n_429), .B2(n_419), .C(n_417), .Y(n_684) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_589), .A2(n_419), .B(n_429), .C(n_417), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_572), .A2(n_429), .B(n_419), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_662), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g688 ( .A1(n_578), .A2(n_430), .B1(n_429), .B2(n_419), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_578), .A2(n_429), .B1(n_430), .B2(n_419), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_586), .B(n_15), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_590), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_606), .B(n_17), .Y(n_692) );
INVx5_ASAP7_75t_L g693 ( .A(n_644), .Y(n_693) );
OAI21xp5_ASAP7_75t_L g694 ( .A1(n_626), .A2(n_430), .B(n_119), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_579), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_585), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_595), .A2(n_22), .B1(n_19), .B2(n_20), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_581), .A2(n_24), .B(n_22), .C(n_23), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_670), .A2(n_27), .B1(n_25), .B2(n_26), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_570), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_663), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_619), .Y(n_702) );
BUFx10_ASAP7_75t_L g703 ( .A(n_651), .Y(n_703) );
OAI22xp33_ASAP7_75t_L g704 ( .A1(n_592), .A2(n_630), .B1(n_593), .B2(n_651), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_576), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_658), .A2(n_121), .B(n_120), .Y(n_706) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_639), .A2(n_124), .B(n_122), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_651), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_583), .B(n_30), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_584), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_665), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_599), .B(n_31), .Y(n_712) );
BUFx10_ASAP7_75t_L g713 ( .A(n_676), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_605), .B(n_32), .Y(n_714) );
NAND2x1_ASAP7_75t_L g715 ( .A(n_627), .B(n_126), .Y(n_715) );
NOR2xp67_ASAP7_75t_L g716 ( .A(n_623), .B(n_33), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_653), .A2(n_130), .B(n_128), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_665), .B(n_33), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_637), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_620), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_720) );
OAI22x1_ASAP7_75t_L g721 ( .A1(n_609), .A2(n_34), .B1(n_36), .B2(n_37), .Y(n_721) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_600), .A2(n_39), .B1(n_40), .B2(n_41), .Y(n_722) );
INVx3_ASAP7_75t_SL g723 ( .A(n_668), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_580), .B(n_42), .Y(n_724) );
INVx1_ASAP7_75t_SL g725 ( .A(n_656), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_621), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_577), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g728 ( .A1(n_604), .A2(n_133), .B(n_132), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_580), .B(n_46), .Y(n_729) );
CKINVDCx6p67_ASAP7_75t_R g730 ( .A(n_652), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_666), .A2(n_50), .B(n_51), .C(n_52), .Y(n_731) );
CKINVDCx6p67_ASAP7_75t_R g732 ( .A(n_674), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_676), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_677), .B(n_54), .Y(n_734) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_607), .A2(n_56), .B1(n_58), .B2(n_60), .Y(n_735) );
AO31x2_ASAP7_75t_L g736 ( .A1(n_634), .A2(n_58), .A3(n_60), .B(n_61), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g737 ( .A1(n_641), .A2(n_140), .B(n_138), .Y(n_737) );
AO31x2_ASAP7_75t_L g738 ( .A1(n_635), .A2(n_61), .A3(n_62), .B(n_63), .Y(n_738) );
INVx1_ASAP7_75t_SL g739 ( .A(n_674), .Y(n_739) );
BUFx8_ASAP7_75t_L g740 ( .A(n_644), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_602), .A2(n_63), .B1(n_64), .B2(n_65), .C(n_67), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_611), .Y(n_742) );
CKINVDCx11_ASAP7_75t_R g743 ( .A(n_627), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_669), .B(n_68), .Y(n_744) );
AND2x4_ASAP7_75t_L g745 ( .A(n_667), .B(n_68), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g746 ( .A1(n_671), .A2(n_146), .B(n_144), .Y(n_746) );
BUFx2_ASAP7_75t_L g747 ( .A(n_577), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_617), .Y(n_748) );
INVx5_ASAP7_75t_L g749 ( .A(n_582), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_571), .B(n_70), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_673), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_751) );
OR2x2_ASAP7_75t_L g752 ( .A(n_608), .B(n_594), .Y(n_752) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_672), .A2(n_75), .B(n_76), .C(n_77), .Y(n_753) );
AND2x4_ASAP7_75t_L g754 ( .A(n_667), .B(n_77), .Y(n_754) );
OR2x6_ASAP7_75t_L g755 ( .A(n_612), .B(n_79), .Y(n_755) );
AOI221xp5_ASAP7_75t_SL g756 ( .A1(n_654), .A2(n_79), .B1(n_80), .B2(n_81), .C(n_82), .Y(n_756) );
OAI21xp5_ASAP7_75t_L g757 ( .A1(n_640), .A2(n_149), .B(n_147), .Y(n_757) );
AND2x4_ASAP7_75t_L g758 ( .A(n_618), .B(n_80), .Y(n_758) );
OAI21xp5_ASAP7_75t_L g759 ( .A1(n_638), .A2(n_629), .B(n_657), .Y(n_759) );
INVx4_ASAP7_75t_L g760 ( .A(n_582), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_SL g761 ( .A1(n_648), .A2(n_650), .B(n_661), .C(n_646), .Y(n_761) );
A2O1A1Ixp33_ASAP7_75t_L g762 ( .A1(n_631), .A2(n_81), .B(n_82), .C(n_83), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_575), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_675), .Y(n_764) );
A2O1A1Ixp33_ASAP7_75t_L g765 ( .A1(n_643), .A2(n_83), .B(n_84), .C(n_86), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_597), .B(n_87), .Y(n_766) );
AO32x2_ASAP7_75t_L g767 ( .A1(n_625), .A2(n_87), .A3(n_88), .B1(n_89), .B2(n_90), .Y(n_767) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_596), .B(n_88), .C(n_90), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g769 ( .A1(n_655), .A2(n_91), .B(n_92), .C(n_93), .Y(n_769) );
NOR2xp33_ASAP7_75t_SL g770 ( .A(n_582), .B(n_92), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g771 ( .A1(n_628), .A2(n_93), .B(n_94), .C(n_96), .Y(n_771) );
INVx4_ASAP7_75t_L g772 ( .A(n_601), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_645), .B(n_97), .Y(n_773) );
AO31x2_ASAP7_75t_L g774 ( .A1(n_647), .A2(n_98), .A3(n_99), .B(n_100), .Y(n_774) );
AOI221xp5_ASAP7_75t_L g775 ( .A1(n_649), .A2(n_99), .B1(n_102), .B2(n_103), .C(n_105), .Y(n_775) );
OR2x6_ASAP7_75t_L g776 ( .A(n_601), .B(n_102), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_613), .B(n_105), .Y(n_777) );
BUFx12f_ASAP7_75t_L g778 ( .A(n_659), .Y(n_778) );
O2A1O1Ixp33_ASAP7_75t_SL g779 ( .A1(n_622), .A2(n_190), .B(n_256), .C(n_255), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_633), .A2(n_106), .B(n_107), .C(n_108), .Y(n_780) );
BUFx3_ASAP7_75t_L g781 ( .A(n_624), .Y(n_781) );
A2O1A1Ixp33_ASAP7_75t_L g782 ( .A1(n_610), .A2(n_110), .B(n_111), .C(n_112), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g783 ( .A1(n_610), .A2(n_112), .B(n_113), .C(n_114), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_632), .A2(n_115), .B1(n_150), .B2(n_151), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_587), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g786 ( .A1(n_636), .A2(n_152), .B1(n_155), .B2(n_156), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_642), .Y(n_787) );
INVx1_ASAP7_75t_SL g788 ( .A(n_616), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_588), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_591), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g791 ( .A(n_664), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_660), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_660), .Y(n_793) );
AO32x2_ASAP7_75t_L g794 ( .A1(n_573), .A2(n_159), .A3(n_160), .B1(n_161), .B2(n_162), .Y(n_794) );
AND2x4_ASAP7_75t_L g795 ( .A(n_665), .B(n_265), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_574), .B(n_177), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_603), .A2(n_178), .B1(n_179), .B2(n_180), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_742), .B(n_693), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_693), .B(n_187), .Y(n_799) );
NOR2x1_ASAP7_75t_SL g800 ( .A(n_776), .B(n_188), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_683), .A2(n_198), .B1(n_199), .B2(n_201), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_719), .Y(n_802) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_748), .A2(n_205), .B1(n_210), .B2(n_212), .C(n_213), .Y(n_803) );
INVx2_ASAP7_75t_SL g804 ( .A(n_740), .Y(n_804) );
INVxp67_ASAP7_75t_L g805 ( .A(n_740), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_696), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_687), .B(n_221), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_705), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_776), .A2(n_226), .B1(n_227), .B2(n_228), .Y(n_809) );
AND2x4_ASAP7_75t_L g810 ( .A(n_693), .B(n_229), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_704), .A2(n_236), .B1(n_237), .B2(n_240), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_691), .Y(n_812) );
INVx2_ASAP7_75t_L g813 ( .A(n_726), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_752), .B(n_246), .Y(n_814) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_750), .A2(n_247), .B(n_249), .C(n_250), .Y(n_815) );
OR2x2_ASAP7_75t_L g816 ( .A(n_700), .B(n_251), .Y(n_816) );
OR2x6_ASAP7_75t_L g817 ( .A(n_679), .B(n_253), .Y(n_817) );
INVx3_ASAP7_75t_L g818 ( .A(n_778), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_695), .Y(n_819) );
AND2x4_ASAP7_75t_L g820 ( .A(n_708), .B(n_747), .Y(n_820) );
CKINVDCx6p67_ASAP7_75t_R g821 ( .A(n_678), .Y(n_821) );
AND2x4_ASAP7_75t_L g822 ( .A(n_749), .B(n_795), .Y(n_822) );
AND2x4_ASAP7_75t_L g823 ( .A(n_749), .B(n_795), .Y(n_823) );
OA21x2_ASAP7_75t_L g824 ( .A1(n_757), .A2(n_707), .B(n_756), .Y(n_824) );
AO21x2_ASAP7_75t_L g825 ( .A1(n_685), .A2(n_779), .B(n_777), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_766), .A2(n_745), .B1(n_718), .B2(n_754), .Y(n_826) );
INVx3_ASAP7_75t_L g827 ( .A(n_732), .Y(n_827) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_793), .Y(n_828) );
OAI21xp5_ASAP7_75t_L g829 ( .A1(n_759), .A2(n_712), .B(n_714), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_764), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_718), .A2(n_745), .B1(n_754), .B2(n_734), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_713), .B(n_724), .Y(n_832) );
INVx5_ASAP7_75t_L g833 ( .A(n_703), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_755), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_692), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g836 ( .A1(n_701), .A2(n_744), .B1(n_773), .B2(n_758), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g837 ( .A1(n_746), .A2(n_737), .B(n_728), .Y(n_837) );
NOR2xp67_ASAP7_75t_SL g838 ( .A(n_680), .B(n_791), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_709), .B(n_788), .Y(n_839) );
OAI21x1_ASAP7_75t_L g840 ( .A1(n_715), .A2(n_717), .B(n_706), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_713), .B(n_729), .Y(n_841) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_749), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_763), .Y(n_843) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_743), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_796), .B(n_781), .Y(n_845) );
AOI21xp5_ASAP7_75t_L g846 ( .A1(n_790), .A2(n_684), .B(n_789), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_730), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_703), .B(n_690), .Y(n_848) );
OAI21xp5_ASAP7_75t_L g849 ( .A1(n_698), .A2(n_783), .B(n_782), .Y(n_849) );
INVx3_ASAP7_75t_L g850 ( .A(n_760), .Y(n_850) );
AOI21xp5_ASAP7_75t_L g851 ( .A1(n_770), .A2(n_786), .B(n_785), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g852 ( .A1(n_765), .A2(n_722), .B(n_771), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_780), .A2(n_731), .B(n_753), .Y(n_853) );
AO21x2_ASAP7_75t_L g854 ( .A1(n_769), .A2(n_762), .B(n_768), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_751), .Y(n_855) );
AO31x2_ASAP7_75t_L g856 ( .A1(n_735), .A2(n_699), .A3(n_772), .B(n_720), .Y(n_856) );
NAND2x1p5_ASAP7_75t_L g857 ( .A(n_739), .B(n_710), .Y(n_857) );
BUFx4f_ASAP7_75t_L g858 ( .A(n_723), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_711), .A2(n_758), .B(n_689), .Y(n_859) );
OA21x2_ASAP7_75t_L g860 ( .A1(n_784), .A2(n_775), .B(n_741), .Y(n_860) );
OR2x2_ASAP7_75t_L g861 ( .A(n_697), .B(n_711), .Y(n_861) );
AO21x2_ASAP7_75t_L g862 ( .A1(n_681), .A2(n_727), .B(n_716), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_721), .B(n_738), .Y(n_863) );
AOI321xp33_ASAP7_75t_L g864 ( .A1(n_797), .A2(n_767), .A3(n_738), .B1(n_736), .B2(n_774), .C(n_794), .Y(n_864) );
AND2x2_ASAP7_75t_L g865 ( .A(n_767), .B(n_774), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_736), .B(n_774), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_736), .B(n_688), .Y(n_867) );
AND2x4_ASAP7_75t_L g868 ( .A(n_767), .B(n_742), .Y(n_868) );
INVx2_ASAP7_75t_SL g869 ( .A(n_740), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_702), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_702), .B(n_742), .Y(n_871) );
OR2x6_ASAP7_75t_L g872 ( .A(n_679), .B(n_792), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_678), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_702), .B(n_742), .Y(n_874) );
BUFx3_ASAP7_75t_L g875 ( .A(n_679), .Y(n_875) );
BUFx4f_ASAP7_75t_SL g876 ( .A(n_679), .Y(n_876) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_679), .Y(n_877) );
BUFx8_ASAP7_75t_L g878 ( .A(n_679), .Y(n_878) );
INVx2_ASAP7_75t_L g879 ( .A(n_719), .Y(n_879) );
OR2x6_ASAP7_75t_L g880 ( .A(n_679), .B(n_792), .Y(n_880) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_686), .A2(n_761), .B(n_572), .Y(n_881) );
OR2x2_ASAP7_75t_L g882 ( .A(n_725), .B(n_526), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_719), .Y(n_883) );
AO21x2_ASAP7_75t_L g884 ( .A1(n_694), .A2(n_787), .B(n_615), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_702), .B(n_742), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_682), .A2(n_614), .B(n_527), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g887 ( .A(n_702), .B(n_742), .Y(n_887) );
INVxp67_ASAP7_75t_SL g888 ( .A(n_740), .Y(n_888) );
INVx2_ASAP7_75t_L g889 ( .A(n_719), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_702), .B(n_742), .Y(n_890) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_740), .Y(n_891) );
OAI21xp5_ASAP7_75t_L g892 ( .A1(n_682), .A2(n_614), .B(n_527), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_702), .B(n_598), .Y(n_893) );
INVx1_ASAP7_75t_SL g894 ( .A(n_733), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_702), .Y(n_895) );
BUFx12f_ASAP7_75t_L g896 ( .A(n_679), .Y(n_896) );
INVx3_ASAP7_75t_L g897 ( .A(n_740), .Y(n_897) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_686), .A2(n_761), .B(n_572), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_686), .A2(n_761), .B(n_572), .Y(n_899) );
AO21x2_ASAP7_75t_L g900 ( .A1(n_866), .A2(n_867), .B(n_863), .Y(n_900) );
INVx2_ASAP7_75t_SL g901 ( .A(n_833), .Y(n_901) );
OR2x6_ASAP7_75t_L g902 ( .A(n_822), .B(n_823), .Y(n_902) );
OR2x2_ASAP7_75t_L g903 ( .A(n_836), .B(n_868), .Y(n_903) );
INVx1_ASAP7_75t_SL g904 ( .A(n_873), .Y(n_904) );
OR2x6_ASAP7_75t_L g905 ( .A(n_822), .B(n_823), .Y(n_905) );
AND2x2_ASAP7_75t_L g906 ( .A(n_879), .B(n_883), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_868), .Y(n_907) );
AND2x2_ASAP7_75t_L g908 ( .A(n_889), .B(n_819), .Y(n_908) );
BUFx3_ASAP7_75t_L g909 ( .A(n_878), .Y(n_909) );
OR2x6_ASAP7_75t_L g910 ( .A(n_817), .B(n_809), .Y(n_910) );
INVx3_ASAP7_75t_L g911 ( .A(n_842), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_893), .B(n_870), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_813), .B(n_802), .Y(n_913) );
OA21x2_ASAP7_75t_L g914 ( .A1(n_886), .A2(n_892), .B(n_899), .Y(n_914) );
OA21x2_ASAP7_75t_L g915 ( .A1(n_892), .A2(n_898), .B(n_881), .Y(n_915) );
OR2x6_ASAP7_75t_L g916 ( .A(n_817), .B(n_799), .Y(n_916) );
AND2x2_ASAP7_75t_L g917 ( .A(n_806), .B(n_808), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_812), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_830), .B(n_843), .Y(n_919) );
BUFx6f_ASAP7_75t_L g920 ( .A(n_842), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_865), .Y(n_921) );
OR2x6_ASAP7_75t_L g922 ( .A(n_817), .B(n_799), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_895), .B(n_871), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_855), .B(n_831), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_826), .B(n_894), .Y(n_925) );
INVx1_ASAP7_75t_L g926 ( .A(n_864), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_864), .Y(n_927) );
AND2x2_ASAP7_75t_L g928 ( .A(n_835), .B(n_798), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_798), .B(n_829), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_878), .Y(n_930) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_894), .Y(n_931) );
INVx2_ASAP7_75t_SL g932 ( .A(n_833), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_874), .Y(n_933) );
BUFx2_ASAP7_75t_L g934 ( .A(n_834), .Y(n_934) );
OR2x2_ASAP7_75t_L g935 ( .A(n_839), .B(n_882), .Y(n_935) );
CKINVDCx14_ASAP7_75t_R g936 ( .A(n_847), .Y(n_936) );
OR2x6_ASAP7_75t_L g937 ( .A(n_810), .B(n_859), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_885), .B(n_887), .Y(n_938) );
BUFx5_ASAP7_75t_L g939 ( .A(n_810), .Y(n_939) );
AOI221xp5_ASAP7_75t_SL g940 ( .A1(n_853), .A2(n_852), .B1(n_845), .B2(n_814), .C(n_846), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_861), .A2(n_854), .B1(n_860), .B2(n_848), .Y(n_941) );
OA21x2_ASAP7_75t_L g942 ( .A1(n_837), .A2(n_849), .B(n_840), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_890), .Y(n_943) );
BUFx2_ASAP7_75t_L g944 ( .A(n_850), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_854), .B(n_807), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_860), .A2(n_849), .B1(n_832), .B2(n_841), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_850), .B(n_800), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_816), .Y(n_948) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_801), .A2(n_811), .B1(n_851), .B2(n_857), .Y(n_949) );
INVxp67_ASAP7_75t_L g950 ( .A(n_888), .Y(n_950) );
AO21x2_ASAP7_75t_L g951 ( .A1(n_884), .A2(n_862), .B(n_825), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_820), .B(n_827), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g953 ( .A(n_827), .B(n_818), .Y(n_953) );
INVx4_ASAP7_75t_L g954 ( .A(n_897), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g955 ( .A1(n_891), .A2(n_805), .B1(n_804), .B2(n_869), .C(n_880), .Y(n_955) );
BUFx2_ASAP7_75t_L g956 ( .A(n_856), .Y(n_956) );
BUFx2_ASAP7_75t_SL g957 ( .A(n_897), .Y(n_957) );
OR2x2_ASAP7_75t_L g958 ( .A(n_856), .B(n_824), .Y(n_958) );
OA21x2_ASAP7_75t_L g959 ( .A1(n_815), .A2(n_803), .B(n_828), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_872), .Y(n_960) );
OR2x6_ASAP7_75t_L g961 ( .A(n_872), .B(n_880), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_872), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_880), .Y(n_963) );
AO21x2_ASAP7_75t_L g964 ( .A1(n_858), .A2(n_844), .B(n_821), .Y(n_964) );
OAI221xp5_ASAP7_75t_L g965 ( .A1(n_858), .A2(n_875), .B1(n_844), .B2(n_877), .C(n_838), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_844), .B(n_896), .Y(n_966) );
BUFx4f_ASAP7_75t_SL g967 ( .A(n_876), .Y(n_967) );
AO21x2_ASAP7_75t_L g968 ( .A1(n_866), .A2(n_867), .B(n_863), .Y(n_968) );
AO21x2_ASAP7_75t_L g969 ( .A1(n_866), .A2(n_867), .B(n_863), .Y(n_969) );
NOR2xp33_ASAP7_75t_L g970 ( .A(n_950), .B(n_904), .Y(n_970) );
INVx1_ASAP7_75t_SL g971 ( .A(n_957), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_921), .B(n_926), .Y(n_972) );
INVx5_ASAP7_75t_SL g973 ( .A(n_916), .Y(n_973) );
NAND2xp5_ASAP7_75t_L g974 ( .A(n_933), .B(n_943), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_927), .B(n_903), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_907), .B(n_924), .Y(n_976) );
BUFx2_ASAP7_75t_L g977 ( .A(n_910), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_924), .B(n_903), .Y(n_978) );
OR2x6_ASAP7_75t_L g979 ( .A(n_910), .B(n_937), .Y(n_979) );
HB1xp67_ASAP7_75t_L g980 ( .A(n_931), .Y(n_980) );
AND2x2_ASAP7_75t_L g981 ( .A(n_956), .B(n_917), .Y(n_981) );
OR2x2_ASAP7_75t_L g982 ( .A(n_935), .B(n_925), .Y(n_982) );
AND2x2_ASAP7_75t_L g983 ( .A(n_945), .B(n_918), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_900), .B(n_968), .Y(n_984) );
HB1xp67_ASAP7_75t_L g985 ( .A(n_908), .Y(n_985) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_916), .Y(n_986) );
BUFx2_ASAP7_75t_L g987 ( .A(n_937), .Y(n_987) );
OR2x2_ASAP7_75t_L g988 ( .A(n_925), .B(n_938), .Y(n_988) );
BUFx3_ASAP7_75t_L g989 ( .A(n_916), .Y(n_989) );
AND2x2_ASAP7_75t_L g990 ( .A(n_900), .B(n_968), .Y(n_990) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_922), .Y(n_991) );
OR2x6_ASAP7_75t_L g992 ( .A(n_937), .B(n_922), .Y(n_992) );
INVx4_ASAP7_75t_L g993 ( .A(n_939), .Y(n_993) );
AND2x2_ASAP7_75t_L g994 ( .A(n_969), .B(n_919), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_958), .B(n_941), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_958), .Y(n_996) );
BUFx2_ASAP7_75t_L g997 ( .A(n_939), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_913), .B(n_906), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_912), .B(n_923), .Y(n_999) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_944), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_929), .B(n_946), .Y(n_1001) );
OR2x2_ASAP7_75t_L g1002 ( .A(n_982), .B(n_914), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_983), .B(n_914), .Y(n_1003) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_982), .B(n_914), .Y(n_1004) );
INVx3_ASAP7_75t_L g1005 ( .A(n_993), .Y(n_1005) );
INVx1_ASAP7_75t_SL g1006 ( .A(n_971), .Y(n_1006) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_976), .B(n_929), .Y(n_1007) );
NAND2x1p5_ASAP7_75t_L g1008 ( .A(n_993), .B(n_947), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_993), .Y(n_1009) );
OR2x6_ASAP7_75t_L g1010 ( .A(n_979), .B(n_961), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_988), .B(n_934), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1012 ( .A(n_992), .Y(n_1012) );
OR2x2_ASAP7_75t_L g1013 ( .A(n_988), .B(n_934), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1014 ( .A(n_978), .B(n_951), .Y(n_1014) );
INVx5_ASAP7_75t_L g1015 ( .A(n_992), .Y(n_1015) );
CKINVDCx16_ASAP7_75t_R g1016 ( .A(n_998), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_978), .B(n_951), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1018 ( .A(n_994), .B(n_915), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_975), .B(n_960), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_972), .B(n_963), .Y(n_1020) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_985), .B(n_928), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g1022 ( .A(n_1000), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_981), .B(n_942), .Y(n_1023) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_972), .B(n_961), .Y(n_1024) );
NOR2xp33_ASAP7_75t_L g1025 ( .A(n_999), .B(n_955), .Y(n_1025) );
INVx3_ASAP7_75t_SL g1026 ( .A(n_1006), .Y(n_1026) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_1016), .B(n_995), .Y(n_1027) );
NAND3xp33_ASAP7_75t_L g1028 ( .A(n_1025), .B(n_980), .C(n_970), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_1005), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_1018), .B(n_984), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1018), .B(n_990), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_1002), .B(n_995), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_1002), .B(n_1001), .Y(n_1033) );
AND2x2_ASAP7_75t_SL g1034 ( .A(n_1012), .B(n_977), .Y(n_1034) );
OR2x2_ASAP7_75t_L g1035 ( .A(n_1004), .B(n_1001), .Y(n_1035) );
AND2x4_ASAP7_75t_L g1036 ( .A(n_1015), .B(n_1010), .Y(n_1036) );
INVx2_ASAP7_75t_SL g1037 ( .A(n_1005), .Y(n_1037) );
OAI32xp33_ASAP7_75t_L g1038 ( .A1(n_1011), .A2(n_986), .A3(n_991), .B1(n_989), .B2(n_909), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1003), .B(n_979), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_1003), .B(n_979), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_1010), .A2(n_979), .B1(n_992), .B2(n_989), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_1023), .B(n_996), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1020), .Y(n_1043) );
NAND2xp5_ASAP7_75t_L g1044 ( .A(n_1019), .B(n_974), .Y(n_1044) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1020), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_1007), .B(n_973), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_1029), .Y(n_1047) );
NOR2xp33_ASAP7_75t_L g1048 ( .A(n_1026), .B(n_964), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1033), .B(n_1004), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_1036), .B(n_1015), .Y(n_1050) );
NOR2x1_ASAP7_75t_L g1051 ( .A(n_1028), .B(n_1009), .Y(n_1051) );
INVx1_ASAP7_75t_SL g1052 ( .A(n_1026), .Y(n_1052) );
OAI22xp33_ASAP7_75t_L g1053 ( .A1(n_1027), .A2(n_1010), .B1(n_1015), .B2(n_1008), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1030), .B(n_1031), .Y(n_1054) );
OAI22xp5_ASAP7_75t_L g1055 ( .A1(n_1027), .A2(n_973), .B1(n_1034), .B2(n_1041), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1042), .B(n_1014), .Y(n_1056) );
INVxp67_ASAP7_75t_SL g1057 ( .A(n_1051), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1049), .Y(n_1058) );
AOI21xp33_ASAP7_75t_L g1059 ( .A1(n_1048), .A2(n_962), .B(n_1024), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1054), .B(n_1035), .Y(n_1060) );
INVx1_ASAP7_75t_SL g1061 ( .A(n_1052), .Y(n_1061) );
AOI211xp5_ASAP7_75t_SL g1062 ( .A1(n_1055), .A2(n_967), .B(n_965), .C(n_949), .Y(n_1062) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_1047), .A2(n_1032), .B1(n_1044), .B2(n_953), .C(n_1037), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_1053), .A2(n_973), .B1(n_1021), .B2(n_1013), .Y(n_1064) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_1056), .B(n_1043), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1056), .B(n_1045), .Y(n_1066) );
O2A1O1Ixp33_ASAP7_75t_L g1067 ( .A1(n_1057), .A2(n_936), .B(n_966), .C(n_1038), .Y(n_1067) );
AOI321xp33_ASAP7_75t_L g1068 ( .A1(n_1062), .A2(n_1050), .A3(n_1039), .B1(n_1040), .B2(n_1022), .C(n_1046), .Y(n_1068) );
A2O1A1Ixp33_ASAP7_75t_SL g1069 ( .A1(n_1063), .A2(n_911), .B(n_952), .C(n_948), .Y(n_1069) );
NOR3xp33_ASAP7_75t_L g1070 ( .A(n_1061), .B(n_930), .C(n_954), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1058), .Y(n_1071) );
NAND3xp33_ASAP7_75t_L g1072 ( .A(n_1068), .B(n_1059), .C(n_1064), .Y(n_1072) );
AOI321xp33_ASAP7_75t_L g1073 ( .A1(n_1067), .A2(n_1064), .A3(n_1060), .B1(n_1066), .B2(n_1065), .C(n_1017), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_1071), .Y(n_1074) );
NOR3xp33_ASAP7_75t_L g1075 ( .A(n_1072), .B(n_1070), .C(n_1069), .Y(n_1075) );
NAND3xp33_ASAP7_75t_SL g1076 ( .A(n_1073), .B(n_1069), .C(n_1008), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1075), .B(n_1074), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g1078 ( .A(n_1076), .Y(n_1078) );
NOR2xp67_ASAP7_75t_L g1079 ( .A(n_1078), .B(n_901), .Y(n_1079) );
AND2x4_ASAP7_75t_L g1080 ( .A(n_1077), .B(n_932), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1080), .Y(n_1081) );
NOR2xp33_ASAP7_75t_L g1082 ( .A(n_1081), .B(n_1079), .Y(n_1082) );
AOI222xp33_ASAP7_75t_SL g1083 ( .A1(n_1082), .A2(n_987), .B1(n_911), .B2(n_997), .C1(n_905), .C2(n_902), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1083), .Y(n_1084) );
AOI21xp33_ASAP7_75t_L g1085 ( .A1(n_1084), .A2(n_920), .B(n_940), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_1085), .A2(n_959), .B(n_920), .Y(n_1086) );
endmodule