module fake_jpeg_2734_n_47 (n_3, n_2, n_1, n_0, n_4, n_5, n_47);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_47;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_2),
.B(n_0),
.Y(n_6)
);

BUFx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_20),
.B1(n_12),
.B2(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_6),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_3),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AO22x1_ASAP7_75t_L g26 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_4),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.C(n_7),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_9),
.A2(n_1),
.B1(n_8),
.B2(n_12),
.Y(n_24)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_11),
.B(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_23),
.A2(n_11),
.B1(n_20),
.B2(n_24),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_15),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_26),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_25),
.A2(n_24),
.B1(n_17),
.B2(n_21),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_35),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_33),
.B(n_28),
.Y(n_37)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_26),
.B(n_25),
.Y(n_38)
);

OAI321xp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_25),
.A3(n_32),
.B1(n_27),
.B2(n_19),
.C(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_36),
.C(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

MAJx2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_38),
.C(n_31),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_41),
.B1(n_38),
.B2(n_44),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_41),
.Y(n_47)
);


endmodule