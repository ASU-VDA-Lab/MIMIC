module fake_jpeg_30687_n_375 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_375);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_375;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx11_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_51),
.Y(n_91)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_15),
.A2(n_14),
.B1(n_13),
.B2(n_2),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_15),
.B1(n_30),
.B2(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_54),
.Y(n_131)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_63),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_61),
.B(n_67),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_14),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g110 ( 
.A(n_66),
.Y(n_110)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_71),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_73),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_13),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_41),
.B(n_1),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_76),
.B(n_4),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_32),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_80),
.Y(n_118)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_40),
.B(n_22),
.Y(n_92)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_33),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_40),
.C(n_25),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_85),
.B(n_125),
.C(n_102),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_25),
.B1(n_23),
.B2(n_31),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_87),
.A2(n_106),
.B1(n_112),
.B2(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_41),
.B1(n_30),
.B2(n_15),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_93),
.B1(n_121),
.B2(n_123),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_92),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_23),
.B1(n_25),
.B2(n_31),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_96),
.A2(n_6),
.B1(n_7),
.B2(n_123),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_30),
.B1(n_27),
.B2(n_29),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_100),
.B1(n_113),
.B2(n_119),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_93),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_56),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_29),
.B1(n_27),
.B2(n_33),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_80),
.A2(n_26),
.B1(n_20),
.B2(n_22),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_38),
.B1(n_36),
.B2(n_21),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_26),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_69),
.Y(n_138)
);

OA22x2_ASAP7_75t_SL g117 ( 
.A1(n_50),
.A2(n_22),
.B1(n_20),
.B2(n_38),
.Y(n_117)
);

AO22x1_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_92),
.B1(n_103),
.B2(n_127),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_43),
.A2(n_47),
.B1(n_36),
.B2(n_21),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_70),
.B1(n_73),
.B2(n_61),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_46),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_124),
.A2(n_125),
.B1(n_129),
.B2(n_102),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_55),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_122),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_132),
.B(n_161),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_133),
.B(n_134),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_48),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_88),
.B(n_74),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_135),
.B(n_97),
.C(n_114),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_65),
.B1(n_44),
.B2(n_64),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_137),
.A2(n_146),
.B1(n_162),
.B2(n_131),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_154),
.Y(n_181)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g141 ( 
.A(n_117),
.B(n_75),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_156),
.Y(n_198)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_6),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_172),
.Y(n_186)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_147),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_91),
.B(n_7),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_149),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_7),
.Y(n_149)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_150),
.Y(n_207)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_151),
.B(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_104),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_85),
.B(n_96),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_155),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_156),
.B(n_167),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_157),
.B(n_158),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_84),
.B(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_160),
.B(n_165),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_101),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_117),
.B1(n_89),
.B2(n_83),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_144),
.B1(n_139),
.B2(n_164),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_101),
.B(n_102),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_109),
.Y(n_178)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_101),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_171),
.Y(n_208)
);

BUFx24_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

CKINVDCx11_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_103),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_170),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_127),
.B(n_126),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_105),
.B(n_83),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_94),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_174),
.B(n_171),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_105),
.B(n_94),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_109),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_R g177 ( 
.A(n_166),
.B(n_145),
.Y(n_177)
);

NOR2x1_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_178),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_189),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_97),
.B(n_114),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_169),
.B(n_197),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_206),
.B1(n_142),
.B2(n_150),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_132),
.B(n_131),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_190),
.B(n_185),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_158),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_194),
.C(n_215),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_138),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_199),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_164),
.B(n_157),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_198),
.A2(n_210),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_156),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_213),
.B1(n_193),
.B2(n_180),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_146),
.A2(n_141),
.B1(n_163),
.B2(n_161),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_144),
.B(n_172),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_135),
.A2(n_176),
.A3(n_154),
.B1(n_153),
.B2(n_167),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_135),
.A2(n_170),
.B1(n_165),
.B2(n_174),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_140),
.B(n_147),
.C(n_151),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_221),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_217),
.A2(n_219),
.B1(n_222),
.B2(n_189),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_218),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_210),
.A2(n_169),
.B1(n_192),
.B2(n_206),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_192),
.A2(n_169),
.B1(n_182),
.B2(n_205),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_229),
.B(n_237),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_200),
.B1(n_191),
.B2(n_177),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_234),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_233),
.Y(n_261)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_181),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_239),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_200),
.A2(n_197),
.B(n_181),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_184),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_196),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_244),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_181),
.B(n_208),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_241),
.A2(n_246),
.B(n_215),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_194),
.B(n_185),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_242),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_207),
.A2(n_201),
.B1(n_179),
.B2(n_198),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_207),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_247),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_274),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_240),
.B(n_183),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_250),
.B(n_252),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_195),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_218),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_221),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_258),
.A2(n_259),
.B1(n_270),
.B2(n_271),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_186),
.B1(n_204),
.B2(n_179),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_260),
.A2(n_266),
.B(n_255),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_201),
.C(n_220),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_264),
.B(n_273),
.C(n_242),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_228),
.A2(n_245),
.B(n_224),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_222),
.A2(n_243),
.B1(n_233),
.B2(n_227),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_217),
.B1(n_219),
.B2(n_216),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_220),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_229),
.A2(n_242),
.B1(n_237),
.B2(n_232),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_224),
.B(n_234),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_265),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_276),
.Y(n_310)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_282),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_267),
.A2(n_223),
.B(n_229),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_280),
.B(n_298),
.CI(n_249),
.CON(n_305),
.SN(n_305)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_291),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_265),
.B(n_266),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_230),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_284),
.B(n_287),
.Y(n_311)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_285),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_241),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_286),
.B(n_270),
.Y(n_299)
);

OA21x2_ASAP7_75t_L g287 ( 
.A1(n_257),
.A2(n_247),
.B(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_289),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_248),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_268),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_294),
.C(n_296),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_244),
.C(n_231),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_295),
.B(n_297),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_264),
.B(n_258),
.C(n_274),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_267),
.A2(n_255),
.B(n_263),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_308),
.B1(n_314),
.B2(n_283),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_278),
.A2(n_271),
.B1(n_257),
.B2(n_259),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_301),
.A2(n_293),
.B1(n_287),
.B2(n_294),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_260),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_302),
.B(n_305),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_276),
.A2(n_254),
.B1(n_256),
.B2(n_269),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_306),
.A2(n_279),
.B1(n_284),
.B2(n_277),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_252),
.B1(n_275),
.B2(n_269),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_285),
.A2(n_254),
.B(n_253),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_287),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_253),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_293),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_290),
.A3(n_282),
.B1(n_288),
.B2(n_289),
.C1(n_295),
.C2(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_318),
.B(n_323),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_302),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_320),
.B(n_321),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_304),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_307),
.Y(n_322)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_310),
.A2(n_286),
.B1(n_311),
.B2(n_278),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_324),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_325),
.A2(n_330),
.B1(n_311),
.B2(n_306),
.Y(n_334)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_327),
.B1(n_331),
.B2(n_333),
.Y(n_335)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_297),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_300),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_294),
.C(n_292),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_312),
.C(n_296),
.Y(n_338)
);

BUFx12_ASAP7_75t_L g331 ( 
.A(n_303),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_309),
.A2(n_277),
.B1(n_262),
.B2(n_248),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_334),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_338),
.B(n_315),
.C(n_319),
.Y(n_352)
);

AOI31xp67_ASAP7_75t_L g339 ( 
.A1(n_320),
.A2(n_287),
.A3(n_313),
.B(n_300),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_305),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_321),
.B(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_340),
.B(n_344),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_343),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_296),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_342),
.A2(n_332),
.B(n_322),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_349),
.A2(n_345),
.B(n_335),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_329),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_351),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_316),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_352),
.B(n_355),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_305),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_338),
.B(n_317),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_360),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_345),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_361),
.B(n_362),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_354),
.B(n_337),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_357),
.B(n_346),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_363),
.B(n_365),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_358),
.A2(n_348),
.B(n_326),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_347),
.C(n_348),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_366),
.B(n_361),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_369),
.A2(n_370),
.B(n_364),
.Y(n_371)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_367),
.A2(n_327),
.A3(n_336),
.B1(n_309),
.B2(n_359),
.C1(n_331),
.C2(n_344),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_371),
.A2(n_372),
.B(n_330),
.Y(n_373)
);

OAI221xp5_ASAP7_75t_SL g372 ( 
.A1(n_368),
.A2(n_328),
.B1(n_325),
.B2(n_313),
.C(n_280),
.Y(n_372)
);

NAND5xp2_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_301),
.C(n_331),
.D(n_341),
.E(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_374),
.Y(n_375)
);


endmodule