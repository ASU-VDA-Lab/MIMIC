module real_aes_416_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_927, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_926, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_927;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_926;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_555;
wire n_421;
wire n_852;
wire n_766;
wire n_919;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_865;
wire n_551;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_615;
wire n_550;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_909;
wire n_523;
wire n_860;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_885;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_880;
wire n_432;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_702;
wire n_912;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_569;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_649;
wire n_749;
wire n_358;
wire n_385;
wire n_397;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_831;
wire n_487;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_789;
wire n_544;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_922;
wire n_633;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_0), .A2(n_323), .B1(n_452), .B2(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_1), .A2(n_281), .B1(n_454), .B2(n_455), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_2), .A2(n_51), .B1(n_363), .B2(n_634), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_3), .A2(n_100), .B1(n_634), .B2(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_4), .A2(n_142), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_5), .A2(n_325), .B1(n_363), .B2(n_634), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_6), .A2(n_236), .B1(n_462), .B2(n_540), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_7), .A2(n_31), .B1(n_394), .B2(n_749), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_8), .A2(n_298), .B1(n_405), .B2(n_525), .Y(n_912) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_9), .A2(n_24), .B1(n_628), .B2(n_710), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_10), .A2(n_274), .B1(n_464), .B2(n_465), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_11), .A2(n_68), .B1(n_467), .B2(n_468), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_12), .Y(n_621) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_13), .A2(n_332), .B1(n_448), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_14), .A2(n_225), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_15), .A2(n_190), .B1(n_426), .B2(n_555), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_16), .A2(n_42), .B1(n_497), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_17), .A2(n_170), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_18), .A2(n_118), .B1(n_451), .B2(n_452), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_19), .A2(n_321), .B1(n_431), .B2(n_436), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_20), .A2(n_120), .B1(n_522), .B2(n_549), .Y(n_857) );
AO22x2_ASAP7_75t_L g813 ( .A1(n_21), .A2(n_814), .B1(n_826), .B2(n_827), .Y(n_813) );
INVx1_ASAP7_75t_L g826 ( .A(n_21), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_22), .A2(n_171), .B1(n_404), .B2(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_23), .A2(n_206), .B1(n_555), .B2(n_717), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_25), .A2(n_161), .B1(n_600), .B2(n_644), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_26), .A2(n_217), .B1(n_458), .B2(n_540), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_27), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g701 ( .A(n_28), .Y(n_701) );
INVx1_ASAP7_75t_SL g358 ( .A(n_29), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g882 ( .A(n_29), .B(n_38), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_30), .A2(n_45), .B1(n_522), .B2(n_595), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_32), .A2(n_287), .B1(n_629), .B2(n_677), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_33), .A2(n_178), .B1(n_452), .B2(n_516), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_34), .A2(n_77), .B1(n_454), .B2(n_455), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_35), .B(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_36), .A2(n_201), .B1(n_461), .B2(n_462), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_37), .B(n_446), .Y(n_533) );
AO22x2_ASAP7_75t_L g361 ( .A1(n_38), .A2(n_308), .B1(n_350), .B2(n_362), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_39), .A2(n_184), .B1(n_493), .B2(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_40), .B(n_446), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_41), .A2(n_265), .B1(n_555), .B2(n_556), .Y(n_554) );
XOR2xp5_ASAP7_75t_L g340 ( .A(n_43), .B(n_341), .Y(n_340) );
XOR2xp5_ASAP7_75t_L g499 ( .A(n_43), .B(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_44), .B(n_636), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_46), .A2(n_80), .B1(n_387), .B2(n_392), .Y(n_386) );
INVx1_ASAP7_75t_L g359 ( .A(n_47), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_48), .A2(n_93), .B1(n_459), .B2(n_465), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_49), .A2(n_191), .B1(n_378), .B2(n_483), .Y(n_816) );
AOI22xp33_ASAP7_75t_SL g903 ( .A1(n_50), .A2(n_289), .B1(n_479), .B2(n_818), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_52), .A2(n_172), .B1(n_599), .B2(n_600), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_53), .A2(n_318), .B1(n_640), .B2(n_757), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_54), .A2(n_128), .B1(n_431), .B2(n_436), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_55), .A2(n_254), .B1(n_489), .B2(n_548), .Y(n_718) );
XNOR2x1_ASAP7_75t_L g673 ( .A(n_56), .B(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_56), .A2(n_674), .B1(n_693), .B2(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_56), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_57), .A2(n_300), .B1(n_780), .B2(n_781), .Y(n_779) );
CKINVDCx20_ASAP7_75t_R g398 ( .A(n_58), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_59), .A2(n_212), .B1(n_467), .B2(n_468), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_60), .A2(n_159), .B1(n_454), .B2(n_582), .Y(n_581) );
AO22x2_ASAP7_75t_L g353 ( .A1(n_61), .A2(n_167), .B1(n_350), .B2(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g838 ( .A1(n_62), .A2(n_326), .B1(n_681), .B2(n_775), .Y(n_838) );
AO22x1_ASAP7_75t_L g851 ( .A1(n_63), .A2(n_247), .B1(n_556), .B2(n_852), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_64), .A2(n_304), .B1(n_496), .B2(n_497), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_65), .Y(n_413) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_66), .A2(n_127), .B1(n_468), .B2(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_67), .A2(n_145), .B1(n_597), .B2(n_647), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g434 ( .A(n_69), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g910 ( .A1(n_70), .A2(n_141), .B1(n_411), .B2(n_551), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_71), .A2(n_202), .B1(n_488), .B2(n_489), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_72), .A2(n_291), .B1(n_448), .B2(n_449), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g803 ( .A1(n_73), .A2(n_197), .B1(n_475), .B2(n_476), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g579 ( .A1(n_74), .A2(n_85), .B1(n_174), .B2(n_446), .C1(n_516), .C2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_75), .A2(n_245), .B1(n_464), .B2(n_465), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_76), .A2(n_176), .B1(n_462), .B2(n_464), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_78), .A2(n_333), .B1(n_516), .B2(n_580), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_79), .A2(n_316), .B1(n_516), .B2(n_580), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g612 ( .A1(n_81), .A2(n_207), .B1(n_613), .B2(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_82), .B(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_83), .A2(n_157), .B1(n_388), .B2(n_706), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_84), .A2(n_131), .B1(n_520), .B2(n_798), .Y(n_797) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_86), .A2(n_110), .B1(n_467), .B2(n_468), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_87), .A2(n_230), .B1(n_345), .B2(n_363), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_88), .A2(n_188), .B1(n_459), .B2(n_465), .Y(n_542) );
OA22x2_ASAP7_75t_L g574 ( .A1(n_89), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_89), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_90), .A2(n_186), .B1(n_600), .B2(n_783), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_91), .A2(n_97), .B1(n_459), .B2(n_462), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_92), .A2(n_257), .B1(n_462), .B2(n_464), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_94), .A2(n_124), .B1(n_436), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_95), .A2(n_195), .B1(n_525), .B2(n_647), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_96), .A2(n_310), .B1(n_467), .B2(n_468), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_98), .A2(n_271), .B1(n_642), .B2(n_757), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_99), .A2(n_203), .B1(n_464), .B2(n_465), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_101), .A2(n_177), .B1(n_628), .B2(n_629), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_102), .A2(n_224), .B1(n_482), .B2(n_630), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_103), .A2(n_223), .B1(n_908), .B2(n_909), .Y(n_907) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_104), .A2(n_135), .B1(n_604), .B2(n_605), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_105), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_106), .A2(n_312), .B1(n_437), .B2(n_464), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_107), .A2(n_192), .B1(n_448), .B2(n_449), .Y(n_659) );
AO22x2_ASAP7_75t_L g349 ( .A1(n_108), .A2(n_250), .B1(n_350), .B2(n_351), .Y(n_349) );
AOI222xp33_ASAP7_75t_SL g685 ( .A1(n_109), .A2(n_237), .B1(n_303), .B2(n_632), .C1(n_636), .C2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_111), .A2(n_204), .B1(n_405), .B2(n_553), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_112), .A2(n_137), .B1(n_364), .B2(n_563), .Y(n_562) );
XOR2x2_ASAP7_75t_L g830 ( .A(n_113), .B(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_114), .A2(n_252), .B1(n_431), .B2(n_551), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_115), .A2(n_329), .B1(n_411), .B2(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_116), .A2(n_290), .B1(n_760), .B2(n_762), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_117), .A2(n_295), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_119), .A2(n_133), .B1(n_620), .B2(n_632), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_121), .A2(n_153), .B1(n_458), .B2(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_122), .A2(n_278), .B1(n_465), .B2(n_642), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_123), .A2(n_185), .B1(n_600), .B2(n_644), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_125), .A2(n_315), .B1(n_620), .B2(n_632), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g892 ( .A1(n_126), .A2(n_893), .B1(n_915), .B2(n_917), .C1(n_921), .C2(n_922), .Y(n_892) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_126), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_129), .A2(n_239), .B1(n_493), .B2(n_522), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_130), .A2(n_156), .B1(n_455), .B2(n_628), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_132), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g514 ( .A1(n_134), .A2(n_160), .B1(n_454), .B2(n_455), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_136), .A2(n_266), .B1(n_458), .B2(n_461), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_138), .A2(n_263), .B1(n_378), .B2(n_772), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_139), .A2(n_211), .B1(n_629), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_140), .A2(n_296), .B1(n_467), .B2(n_468), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_143), .A2(n_282), .B1(n_364), .B2(n_475), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_144), .A2(n_269), .B1(n_480), .B2(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_146), .A2(n_297), .B1(n_467), .B2(n_468), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_147), .A2(n_233), .B1(n_448), .B2(n_584), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_148), .B(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_149), .A2(n_183), .B1(n_619), .B2(n_818), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_150), .A2(n_273), .B1(n_448), .B2(n_449), .Y(n_447) );
AO22x2_ASAP7_75t_L g721 ( .A1(n_151), .A2(n_722), .B1(n_734), .B2(n_735), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_151), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_152), .A2(n_214), .B1(n_437), .B2(n_496), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g758 ( .A1(n_154), .A2(n_168), .B1(n_600), .B2(n_644), .Y(n_758) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_155), .A2(n_327), .B1(n_548), .B2(n_549), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_158), .A2(n_264), .B1(n_448), .B2(n_449), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_162), .A2(n_240), .B1(n_451), .B2(n_580), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_163), .A2(n_280), .B1(n_475), .B2(n_681), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_164), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_165), .A2(n_244), .B1(n_403), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_166), .A2(n_205), .B1(n_451), .B2(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g881 ( .A(n_167), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_169), .A2(n_283), .B1(n_388), .B2(n_686), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_173), .A2(n_260), .B1(n_458), .B2(n_540), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_175), .A2(n_334), .B1(n_464), .B2(n_465), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_179), .A2(n_220), .B1(n_465), .B2(n_522), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_180), .A2(n_218), .B1(n_454), .B2(n_455), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_181), .A2(n_276), .B1(n_491), .B2(n_493), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_182), .B(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_187), .A2(n_246), .B1(n_751), .B2(n_753), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_189), .A2(n_248), .B1(n_404), .B2(n_553), .Y(n_552) );
XOR2x2_ASAP7_75t_L g442 ( .A(n_193), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g754 ( .A(n_194), .B(n_609), .Y(n_754) );
INVx2_ASAP7_75t_L g888 ( .A(n_196), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_198), .A2(n_267), .B1(n_482), .B2(n_483), .Y(n_481) );
XOR2x2_ASAP7_75t_L g768 ( .A(n_199), .B(n_769), .Y(n_768) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_200), .A2(n_259), .B1(n_617), .B2(n_620), .Y(n_616) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_208), .A2(n_314), .B1(n_565), .B2(n_710), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_209), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_210), .A2(n_294), .B1(n_493), .B2(n_640), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_213), .B(n_708), .Y(n_730) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_215), .A2(n_256), .B1(n_479), .B2(n_480), .Y(n_478) );
XNOR2x1_ASAP7_75t_L g530 ( .A(n_216), .B(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_219), .A2(n_249), .B1(n_467), .B2(n_468), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_221), .A2(n_258), .B1(n_410), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_222), .A2(n_272), .B1(n_378), .B2(n_382), .Y(n_377) );
XOR2x2_ASAP7_75t_L g744 ( .A(n_226), .B(n_745), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_227), .A2(n_330), .B1(n_475), .B2(n_476), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_228), .A2(n_286), .B1(n_628), .B2(n_629), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_229), .A2(n_322), .B1(n_403), .B2(n_597), .Y(n_596) );
XOR2xp5_ASAP7_75t_L g469 ( .A(n_231), .B(n_470), .Y(n_469) );
XNOR2x1_ASAP7_75t_L g498 ( .A(n_231), .B(n_470), .Y(n_498) );
INVx1_ASAP7_75t_L g527 ( .A(n_232), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_234), .A2(n_238), .B1(n_464), .B2(n_465), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_235), .A2(n_299), .B1(n_364), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_241), .A2(n_275), .B1(n_458), .B2(n_461), .Y(n_667) );
OA22x2_ASAP7_75t_L g790 ( .A1(n_242), .A2(n_791), .B1(n_792), .B2(n_805), .Y(n_790) );
INVx1_ASAP7_75t_L g805 ( .A(n_242), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_243), .B(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_250), .B(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g891 ( .A(n_251), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_253), .A2(n_302), .B1(n_382), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_255), .A2(n_306), .B1(n_488), .B2(n_715), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_261), .A2(n_285), .B1(n_458), .B2(n_728), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_262), .A2(n_293), .B1(n_364), .B2(n_752), .Y(n_901) );
INVx3_ASAP7_75t_L g350 ( .A(n_268), .Y(n_350) );
XOR2x1_ASAP7_75t_L g624 ( .A(n_270), .B(n_625), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_277), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_279), .A2(n_918), .B1(n_919), .B2(n_920), .Y(n_917) );
CKINVDCx20_ASAP7_75t_R g918 ( .A(n_279), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_284), .B(n_369), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_288), .B(n_636), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_292), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_301), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_305), .A2(n_313), .B1(n_454), .B2(n_582), .Y(n_662) );
INVx1_ASAP7_75t_L g671 ( .A(n_307), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_309), .B(n_708), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_311), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g876 ( .A(n_317), .Y(n_876) );
AND2x4_ASAP7_75t_L g890 ( .A(n_317), .B(n_877), .Y(n_890) );
AO21x1_ASAP7_75t_L g923 ( .A1(n_317), .A2(n_886), .B(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g877 ( .A(n_319), .Y(n_877) );
AND2x2_ASAP7_75t_R g921 ( .A(n_319), .B(n_876), .Y(n_921) );
INVx1_ASAP7_75t_L g850 ( .A(n_320), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_320), .A2(n_846), .B1(n_862), .B2(n_926), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_320), .A2(n_854), .B1(n_858), .B2(n_927), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_320), .B(n_851), .Y(n_864) );
INVxp67_ASAP7_75t_L g887 ( .A(n_324), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_328), .B(n_708), .Y(n_707) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_331), .B(n_545), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_336), .B(n_883), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_650), .B1(n_871), .B2(n_872), .C(n_873), .Y(n_336) );
INVx1_ASAP7_75t_L g871 ( .A(n_337), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_501), .B1(n_648), .B2(n_649), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx3_ASAP7_75t_SL g648 ( .A(n_339), .Y(n_648) );
OA22x2_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_438), .B1(n_439), .B2(n_499), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_396), .C(n_416), .Y(n_341) );
AND3x1_ASAP7_75t_L g500 ( .A(n_342), .B(n_396), .C(n_416), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_376), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_344), .B(n_368), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g613 ( .A(n_346), .Y(n_613) );
INVx2_ASAP7_75t_L g775 ( .A(n_346), .Y(n_775) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx3_ASAP7_75t_L g475 ( .A(n_347), .Y(n_475) );
BUFx5_ASAP7_75t_L g563 ( .A(n_347), .Y(n_563) );
BUFx3_ASAP7_75t_L g752 ( .A(n_347), .Y(n_752) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_355), .Y(n_347) );
AND2x4_ASAP7_75t_L g389 ( .A(n_348), .B(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g437 ( .A(n_348), .B(n_406), .Y(n_437) );
AND2x4_ASAP7_75t_L g448 ( .A(n_348), .B(n_355), .Y(n_448) );
AND2x2_ASAP7_75t_L g451 ( .A(n_348), .B(n_390), .Y(n_451) );
AND2x2_ASAP7_75t_L g462 ( .A(n_348), .B(n_406), .Y(n_462) );
AND2x2_ASAP7_75t_L g516 ( .A(n_348), .B(n_390), .Y(n_516) );
AND2x4_ASAP7_75t_L g348 ( .A(n_349), .B(n_352), .Y(n_348) );
AND2x2_ASAP7_75t_L g366 ( .A(n_349), .B(n_353), .Y(n_366) );
INVx1_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
INVx1_ASAP7_75t_L g381 ( .A(n_349), .Y(n_381) );
INVx2_ASAP7_75t_L g351 ( .A(n_350), .Y(n_351) );
INVx1_ASAP7_75t_L g354 ( .A(n_350), .Y(n_354) );
OAI22x1_ASAP7_75t_L g356 ( .A1(n_350), .A2(n_357), .B1(n_358), .B2(n_359), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_350), .Y(n_357) );
INVx1_ASAP7_75t_L g362 ( .A(n_350), .Y(n_362) );
AND2x4_ASAP7_75t_L g374 ( .A(n_352), .B(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g395 ( .A(n_352), .Y(n_395) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g380 ( .A(n_353), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g379 ( .A(n_355), .B(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g400 ( .A(n_355), .B(n_374), .Y(n_400) );
AND2x4_ASAP7_75t_L g454 ( .A(n_355), .B(n_380), .Y(n_454) );
AND2x2_ASAP7_75t_L g461 ( .A(n_355), .B(n_374), .Y(n_461) );
AND2x2_ASAP7_75t_L g540 ( .A(n_355), .B(n_374), .Y(n_540) );
AND2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_360), .Y(n_355) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_356), .Y(n_367) );
AND2x2_ASAP7_75t_L g373 ( .A(n_356), .B(n_361), .Y(n_373) );
INVx2_ASAP7_75t_L g391 ( .A(n_356), .Y(n_391) );
AND2x4_ASAP7_75t_L g406 ( .A(n_360), .B(n_391), .Y(n_406) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g390 ( .A(n_361), .B(n_391), .Y(n_390) );
BUFx2_ASAP7_75t_L g427 ( .A(n_361), .Y(n_427) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g615 ( .A(n_364), .Y(n_615) );
BUFx12f_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g477 ( .A(n_365), .Y(n_477) );
AND2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
AND2x4_ASAP7_75t_L g405 ( .A(n_366), .B(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g426 ( .A(n_366), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_SL g449 ( .A(n_366), .B(n_367), .Y(n_449) );
AND2x4_ASAP7_75t_L g458 ( .A(n_366), .B(n_406), .Y(n_458) );
AND2x4_ASAP7_75t_L g468 ( .A(n_366), .B(n_427), .Y(n_468) );
AND2x2_ASAP7_75t_SL g584 ( .A(n_366), .B(n_367), .Y(n_584) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx4_ASAP7_75t_SL g473 ( .A(n_371), .Y(n_473) );
INVx3_ASAP7_75t_L g559 ( .A(n_371), .Y(n_559) );
INVx3_ASAP7_75t_SL g611 ( .A(n_371), .Y(n_611) );
INVx3_ASAP7_75t_L g636 ( .A(n_371), .Y(n_636) );
INVx4_ASAP7_75t_SL g708 ( .A(n_371), .Y(n_708) );
INVx6_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
AND2x4_ASAP7_75t_L g383 ( .A(n_373), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g394 ( .A(n_373), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g446 ( .A(n_373), .B(n_374), .Y(n_446) );
AND2x2_ASAP7_75t_L g452 ( .A(n_373), .B(n_395), .Y(n_452) );
AND2x2_ASAP7_75t_L g455 ( .A(n_373), .B(n_384), .Y(n_455) );
AND2x2_ASAP7_75t_L g580 ( .A(n_373), .B(n_395), .Y(n_580) );
AND2x2_ASAP7_75t_L g582 ( .A(n_373), .B(n_384), .Y(n_582) );
AND2x2_ASAP7_75t_L g412 ( .A(n_374), .B(n_390), .Y(n_412) );
AND2x4_ASAP7_75t_L g433 ( .A(n_374), .B(n_406), .Y(n_433) );
AND2x2_ASAP7_75t_L g459 ( .A(n_374), .B(n_406), .Y(n_459) );
AND2x6_ASAP7_75t_L g464 ( .A(n_374), .B(n_390), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_386), .Y(n_376) );
BUFx6f_ASAP7_75t_SL g604 ( .A(n_378), .Y(n_604) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_379), .Y(n_482) );
INVx3_ASAP7_75t_L g566 ( .A(n_379), .Y(n_566) );
AND2x4_ASAP7_75t_L g415 ( .A(n_380), .B(n_406), .Y(n_415) );
AND2x2_ASAP7_75t_L g423 ( .A(n_380), .B(n_390), .Y(n_423) );
AND2x6_ASAP7_75t_L g465 ( .A(n_380), .B(n_406), .Y(n_465) );
AND2x2_ASAP7_75t_L g467 ( .A(n_380), .B(n_390), .Y(n_467) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_381), .Y(n_385) );
BUFx4f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g484 ( .A(n_383), .Y(n_484) );
INVx2_ASAP7_75t_L g607 ( .A(n_383), .Y(n_607) );
BUFx3_ASAP7_75t_L g630 ( .A(n_383), .Y(n_630) );
BUFx6f_ASAP7_75t_SL g710 ( .A(n_383), .Y(n_710) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx4f_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
BUFx2_ASAP7_75t_L g632 ( .A(n_388), .Y(n_632) );
BUFx2_ASAP7_75t_L g749 ( .A(n_388), .Y(n_749) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx2_ASAP7_75t_L g479 ( .A(n_389), .Y(n_479) );
BUFx2_ASAP7_75t_L g561 ( .A(n_389), .Y(n_561) );
BUFx3_ASAP7_75t_L g619 ( .A(n_389), .Y(n_619) );
INVx2_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g480 ( .A(n_393), .Y(n_480) );
INVx2_ASAP7_75t_L g620 ( .A(n_393), .Y(n_620) );
INVx2_ASAP7_75t_L g686 ( .A(n_393), .Y(n_686) );
INVx1_ASAP7_75t_L g706 ( .A(n_393), .Y(n_706) );
INVx2_ASAP7_75t_L g818 ( .A(n_393), .Y(n_818) );
INVx6_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_407), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_401), .B2(n_402), .Y(n_397) );
INVx3_ASAP7_75t_L g553 ( .A(n_399), .Y(n_553) );
INVx1_ASAP7_75t_SL g597 ( .A(n_399), .Y(n_597) );
INVx2_ASAP7_75t_L g689 ( .A(n_399), .Y(n_689) );
INVx2_ASAP7_75t_L g789 ( .A(n_399), .Y(n_789) );
INVx6_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g488 ( .A(n_400), .Y(n_488) );
BUFx3_ASAP7_75t_L g525 ( .A(n_400), .Y(n_525) );
INVxp67_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
BUFx3_ASAP7_75t_L g489 ( .A(n_405), .Y(n_489) );
BUFx2_ASAP7_75t_SL g647 ( .A(n_405), .Y(n_647) );
BUFx2_ASAP7_75t_SL g786 ( .A(n_405), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_413), .B2(n_414), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g492 ( .A(n_412), .Y(n_492) );
BUFx2_ASAP7_75t_L g642 ( .A(n_412), .Y(n_642) );
INVx2_ASAP7_75t_L g497 ( .A(n_414), .Y(n_497) );
INVx2_ASAP7_75t_L g551 ( .A(n_414), .Y(n_551) );
INVx2_ASAP7_75t_SL g595 ( .A(n_414), .Y(n_595) );
INVx2_ASAP7_75t_L g757 ( .A(n_414), .Y(n_757) );
INVx2_ASAP7_75t_L g781 ( .A(n_414), .Y(n_781) );
INVx8_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_428), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B1(n_424), .B2(n_425), .Y(n_417) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_421), .Y(n_783) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_421), .Y(n_852) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g645 ( .A(n_422), .Y(n_645) );
INVx1_ASAP7_75t_L g908 ( .A(n_422), .Y(n_908) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx3_ASAP7_75t_L g520 ( .A(n_423), .Y(n_520) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_423), .Y(n_555) );
INVx2_ASAP7_75t_L g600 ( .A(n_425), .Y(n_600) );
INVx3_ASAP7_75t_L g717 ( .A(n_425), .Y(n_717) );
INVx2_ASAP7_75t_L g909 ( .A(n_425), .Y(n_909) );
INVx5_ASAP7_75t_SL g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g556 ( .A(n_426), .Y(n_556) );
BUFx2_ASAP7_75t_L g798 ( .A(n_426), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_434), .B2(n_435), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
INVx3_ASAP7_75t_SL g522 ( .A(n_432), .Y(n_522) );
INVx2_ASAP7_75t_SL g548 ( .A(n_432), .Y(n_548) );
INVx4_ASAP7_75t_L g728 ( .A(n_432), .Y(n_728) );
INVx8_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g762 ( .A(n_435), .Y(n_762) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_436), .Y(n_788) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g494 ( .A(n_437), .Y(n_494) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_437), .Y(n_715) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_469), .B2(n_498), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_456), .Y(n_443) );
NAND4xp25_ASAP7_75t_SL g444 ( .A(n_445), .B(n_447), .C(n_450), .D(n_453), .Y(n_444) );
INVx2_ASAP7_75t_SL g510 ( .A(n_446), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g456 ( .A(n_457), .B(n_460), .C(n_463), .D(n_466), .Y(n_456) );
OR2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_485), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .C(n_478), .D(n_481), .Y(n_471) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_475), .Y(n_634) );
BUFx6f_ASAP7_75t_L g753 ( .A(n_476), .Y(n_753) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g681 ( .A(n_477), .Y(n_681) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .C(n_490), .D(n_495), .Y(n_485) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g713 ( .A(n_492), .Y(n_713) );
INVx2_ASAP7_75t_SL g780 ( .A(n_492), .Y(n_780) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g549 ( .A(n_494), .Y(n_549) );
INVx1_ASAP7_75t_L g649 ( .A(n_501), .Y(n_649) );
XNOR2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_570), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_528), .B1(n_568), .B2(n_569), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g568 ( .A(n_505), .Y(n_568) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
XOR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_527), .Y(n_506) );
NAND2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_513), .Y(n_508) );
OAI21xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_518), .B(n_523), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_521), .Y(n_518) );
BUFx2_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_526), .Y(n_523) );
INVx2_ASAP7_75t_L g569 ( .A(n_528), .Y(n_569) );
OA22x2_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_543), .B1(n_544), .B2(n_567), .Y(n_528) );
AO22x2_ASAP7_75t_L g573 ( .A1(n_529), .A2(n_530), .B1(n_574), .B2(n_590), .Y(n_573) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_530), .Y(n_567) );
OR2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .Y(n_531) );
NAND4xp25_ASAP7_75t_SL g532 ( .A(n_533), .B(n_534), .C(n_535), .D(n_536), .Y(n_532) );
NAND4xp25_ASAP7_75t_SL g537 ( .A(n_538), .B(n_539), .C(n_541), .D(n_542), .Y(n_537) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp67_ASAP7_75t_L g545 ( .A(n_546), .B(n_557), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .C(n_552), .D(n_554), .Y(n_546) );
NAND4xp25_ASAP7_75t_SL g557 ( .A(n_558), .B(n_560), .C(n_562), .D(n_564), .Y(n_557) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx4_ASAP7_75t_L g628 ( .A(n_566), .Y(n_628) );
INVx1_ASAP7_75t_L g678 ( .A(n_566), .Y(n_678) );
XOR2x1_ASAP7_75t_SL g570 ( .A(n_571), .B(n_623), .Y(n_570) );
AO22x2_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_573), .B1(n_591), .B2(n_622), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g590 ( .A(n_574), .Y(n_590) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_585), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .C(n_583), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_588), .D(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g622 ( .A(n_591), .Y(n_622) );
XOR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_621), .Y(n_591) );
NOR2x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_602), .Y(n_592) );
NAND4xp25_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .C(n_598), .D(n_601), .Y(n_593) );
NAND4xp25_ASAP7_75t_L g602 ( .A(n_603), .B(n_608), .C(n_612), .D(n_616), .Y(n_602) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g772 ( .A(n_607), .Y(n_772) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI21xp33_ASAP7_75t_SL g899 ( .A1(n_610), .A2(n_900), .B(n_901), .Y(n_899) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_611), .Y(n_777) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_637), .Y(n_625) );
NAND4xp25_ASAP7_75t_L g626 ( .A(n_627), .B(n_631), .C(n_633), .D(n_635), .Y(n_626) );
BUFx6f_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND4xp25_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .C(n_643), .D(n_646), .Y(n_637) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g872 ( .A(n_650), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_741), .B1(n_742), .B2(n_867), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_695), .B(n_737), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g867 ( .A1(n_653), .A2(n_868), .B(n_869), .Y(n_867) );
BUFx3_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g738 ( .A(n_654), .Y(n_738) );
OA21x2_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_672), .B(n_691), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_655), .B(n_692), .Y(n_691) );
OA22x2_ASAP7_75t_L g698 ( .A1(n_655), .A2(n_699), .B1(n_700), .B2(n_719), .Y(n_698) );
INVx3_ASAP7_75t_SL g719 ( .A(n_655), .Y(n_719) );
XOR2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_671), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_664), .Y(n_656) );
NOR2xp33_ASAP7_75t_L g657 ( .A(n_658), .B(n_661), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVxp67_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g694 ( .A(n_674), .Y(n_694) );
NAND4xp75_ASAP7_75t_L g674 ( .A(n_675), .B(n_682), .C(n_685), .D(n_687), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
BUFx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g868 ( .A(n_695), .Y(n_868) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OA22x2_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_698), .B1(n_720), .B2(n_736), .Y(n_696) );
OA22x2_ASAP7_75t_L g740 ( .A1(n_697), .A2(n_698), .B1(n_720), .B2(n_736), .Y(n_740) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
XNOR2x2_ASAP7_75t_SL g700 ( .A(n_701), .B(n_702), .Y(n_700) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_711), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .C(n_707), .D(n_709), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .C(n_716), .D(n_718), .Y(n_711) );
INVxp67_ASAP7_75t_L g736 ( .A(n_720), .Y(n_736) );
INVx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g735 ( .A(n_722), .Y(n_735) );
NOR2xp67_ASAP7_75t_L g722 ( .A(n_723), .B(n_729), .Y(n_722) );
NAND4xp25_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .C(n_726), .D(n_727), .Y(n_723) );
INVx2_ASAP7_75t_L g761 ( .A(n_728), .Y(n_761) );
BUFx6f_ASAP7_75t_L g785 ( .A(n_728), .Y(n_785) );
NAND4xp25_ASAP7_75t_SL g729 ( .A(n_730), .B(n_731), .C(n_732), .D(n_733), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g870 ( .A(n_738), .Y(n_870) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_740), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
XNOR2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_808), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_764), .B1(n_765), .B2(n_807), .Y(n_743) );
INVx1_ASAP7_75t_L g807 ( .A(n_744), .Y(n_807) );
NOR2x1_ASAP7_75t_L g745 ( .A(n_746), .B(n_755), .Y(n_745) );
NAND4xp25_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .C(n_750), .D(n_754), .Y(n_746) );
BUFx6f_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
NAND4xp25_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .C(n_759), .D(n_763), .Y(n_755) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
HB1xp67_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AO22x1_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_790), .B2(n_806), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NOR2xp67_ASAP7_75t_L g769 ( .A(n_770), .B(n_778), .Y(n_769) );
NAND4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .C(n_774), .D(n_776), .Y(n_770) );
NAND4xp25_ASAP7_75t_L g778 ( .A(n_779), .B(n_782), .C(n_784), .D(n_787), .Y(n_778) );
INVx1_ASAP7_75t_L g806 ( .A(n_790), .Y(n_806) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
NOR2xp67_ASAP7_75t_L g792 ( .A(n_793), .B(n_800), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_797), .C(n_799), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
NAND4xp25_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .C(n_803), .D(n_804), .Y(n_800) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
OA21x2_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_828), .B(n_865), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_812), .B(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g827 ( .A(n_814), .Y(n_827) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_815), .B(n_821), .Y(n_814) );
NAND4xp25_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .C(n_819), .D(n_820), .Y(n_815) );
NAND4xp25_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .C(n_824), .D(n_825), .Y(n_821) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g866 ( .A(n_829), .Y(n_866) );
XNOR2x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_843), .Y(n_829) );
NOR3xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_837), .C(n_840), .Y(n_831) );
NAND4xp25_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .C(n_835), .D(n_836), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_838), .B(n_839), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NAND4xp75_ASAP7_75t_L g843 ( .A(n_844), .B(n_861), .C(n_863), .D(n_864), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_853), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .C(n_851), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
NAND2xp5_ASAP7_75t_SL g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g862 ( .A(n_849), .Y(n_862) );
NOR2xp67_ASAP7_75t_L g853 ( .A(n_854), .B(n_858), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .C(n_857), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
INVx4_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_878), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_875), .B(n_879), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g875 ( .A(n_876), .B(n_877), .Y(n_875) );
INVx1_ASAP7_75t_L g924 ( .A(n_877), .Y(n_924) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
OAI21xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_891), .B(n_892), .Y(n_883) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_889), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NOR2xp33_ASAP7_75t_L g886 ( .A(n_887), .B(n_888), .Y(n_886) );
INVxp67_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
XNOR2x1_ASAP7_75t_L g896 ( .A(n_897), .B(n_914), .Y(n_896) );
HB1xp67_ASAP7_75t_L g920 ( .A(n_897), .Y(n_920) );
AND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_905), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_902), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_911), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_910), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_912), .B(n_913), .Y(n_911) );
CKINVDCx6p67_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
CKINVDCx20_ASAP7_75t_R g919 ( .A(n_920), .Y(n_919) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_923), .Y(n_922) );
endmodule