module fake_netlist_6_835_n_109 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_109);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_109;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_SL g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

INVxp33_ASAP7_75t_SL g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVxp67_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_2),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_23),
.B1(n_25),
.B2(n_29),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_40),
.B(n_41),
.C(n_38),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

O2A1O1Ixp5_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_46),
.B(n_39),
.C(n_49),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_45),
.B(n_29),
.Y(n_62)
);

CKINVDCx11_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_21),
.B1(n_56),
.B2(n_25),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_60),
.A2(n_23),
.B1(n_42),
.B2(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

O2A1O1Ixp5_ASAP7_75t_L g68 ( 
.A1(n_61),
.A2(n_57),
.B(n_55),
.C(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_42),
.B(n_30),
.C(n_33),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_43),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_73),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_74),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_82),
.B(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_74),
.B(n_75),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_63),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_77),
.B1(n_34),
.B2(n_35),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_31),
.B(n_33),
.Y(n_90)
);

AOI211xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_88),
.B(n_70),
.C(n_31),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_30),
.B(n_68),
.C(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_87),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_48),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_48),
.B1(n_39),
.B2(n_44),
.C(n_50),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_3),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_44),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_98),
.A2(n_52),
.B1(n_5),
.B2(n_6),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_57),
.C(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_4),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_16),
.Y(n_103)
);

AOI221xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_97),
.B1(n_9),
.B2(n_4),
.C(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_102),
.B1(n_99),
.B2(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_103),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_106),
.A2(n_54),
.B1(n_105),
.B2(n_91),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_54),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_54),
.B1(n_106),
.B2(n_107),
.Y(n_109)
);


endmodule