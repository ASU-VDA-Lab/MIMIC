module fake_jpeg_25618_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx8_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_6),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_34),
.B1(n_27),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_47),
.A2(n_50),
.B1(n_52),
.B2(n_30),
.Y(n_85)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_48),
.B(n_29),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_34),
.B1(n_27),
.B2(n_29),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_39),
.B1(n_38),
.B2(n_29),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_33),
.B1(n_26),
.B2(n_17),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_17),
.Y(n_74)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_64),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_31),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g66 ( 
.A(n_35),
.B(n_18),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_36),
.C(n_18),
.Y(n_77)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_74),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_78),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_28),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_49),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_28),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_33),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_23),
.C(n_32),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_63),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_58),
.B1(n_66),
.B2(n_59),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_116),
.B1(n_86),
.B2(n_81),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_66),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_99),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_73),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_66),
.B1(n_39),
.B2(n_51),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_64),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_107),
.Y(n_119)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_64),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g118 ( 
.A1(n_102),
.A2(n_111),
.B(n_96),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_23),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_110),
.Y(n_121)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_13),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_90),
.B1(n_84),
.B2(n_57),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_67),
.B1(n_56),
.B2(n_53),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_123),
.B1(n_65),
.B2(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_124),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_23),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_98),
.B(n_82),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_70),
.C(n_62),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_127),
.C(n_133),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_70),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_128),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_93),
.C(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_23),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_135),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_102),
.B1(n_94),
.B2(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_62),
.C(n_57),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_23),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_22),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_135),
.A2(n_107),
.B1(n_56),
.B2(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_164),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_136),
.A2(n_115),
.B1(n_111),
.B2(n_114),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_151),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_101),
.B1(n_108),
.B2(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_157),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_132),
.A2(n_101),
.B1(n_84),
.B2(n_61),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_122),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_61),
.B1(n_65),
.B2(n_22),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_30),
.B1(n_55),
.B2(n_21),
.Y(n_152)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_55),
.C(n_32),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_133),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_130),
.A2(n_0),
.B(n_1),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_160),
.B(n_119),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_55),
.B1(n_21),
.B2(n_20),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_137),
.A2(n_30),
.B(n_32),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_167),
.B(n_120),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_172),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_153),
.C(n_154),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_128),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_159),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_166),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_176),
.A2(n_180),
.B(n_187),
.Y(n_207)
);

HAxp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_119),
.CON(n_177),
.SN(n_177)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_142),
.C(n_160),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_162),
.B(n_117),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_184),
.B(n_188),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_0),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_123),
.B(n_138),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_18),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_189),
.A2(n_190),
.B1(n_176),
.B2(n_175),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_146),
.B(n_21),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_197),
.C(n_199),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_153),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_195),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_152),
.A3(n_150),
.B1(n_158),
.B2(n_157),
.C1(n_20),
.C2(n_13),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_32),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_186),
.C(n_183),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_20),
.C(n_16),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_181),
.A2(n_20),
.B1(n_16),
.B2(n_15),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_173),
.B1(n_174),
.B2(n_190),
.Y(n_223)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_168),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_181),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_208),
.C(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_210),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_218),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_223),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_178),
.B1(n_174),
.B2(n_190),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_216),
.A2(n_225),
.B1(n_196),
.B2(n_193),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_203),
.B(n_197),
.C(n_207),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_222),
.Y(n_238)
);

BUFx12_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_191),
.C(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_210),
.A2(n_187),
.B1(n_179),
.B2(n_15),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_14),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_208),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_216),
.C(n_220),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_213),
.C(n_224),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_234),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_232),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_12),
.C(n_4),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_12),
.C(n_4),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_6),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_1),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_225),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_240),
.B(n_246),
.Y(n_254)
);

NAND2xp33_ASAP7_75t_R g241 ( 
.A(n_231),
.B(n_217),
.Y(n_241)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_229),
.A2(n_211),
.B(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_233),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_220),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_235),
.A2(n_7),
.B(n_8),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_7),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_227),
.B1(n_233),
.B2(n_10),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_11),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_251),
.B(n_9),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_256),
.B(n_243),
.C(n_9),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_245),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_262),
.A3(n_11),
.B1(n_250),
.B2(n_251),
.C1(n_252),
.C2(n_259),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_260),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_253),
.B(n_239),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_9),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_11),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_265),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_268),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_266),
.Y(n_271)
);


endmodule