module fake_jpeg_31150_n_395 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_395);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_395;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_14),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_46),
.Y(n_90)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_14),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_51),
.Y(n_128)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_52),
.Y(n_100)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_53),
.B(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_13),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_61),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_13),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_77),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_67),
.Y(n_97)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g129 ( 
.A(n_66),
.B(n_68),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_19),
.B(n_13),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_70),
.Y(n_111)
);

CKINVDCx9p33_ASAP7_75t_R g70 ( 
.A(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_72),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_39),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_74),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_76),
.Y(n_117)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_79),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

CKINVDCx9p33_ASAP7_75t_R g84 ( 
.A(n_30),
.Y(n_84)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_24),
.B1(n_32),
.B2(n_2),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_42),
.B1(n_40),
.B2(n_28),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_86),
.A2(n_106),
.B1(n_125),
.B2(n_92),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_35),
.B1(n_40),
.B2(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_87),
.A2(n_116),
.B1(n_119),
.B2(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_60),
.B(n_21),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_93),
.B(n_94),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_21),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_20),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_20),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_22),
.B1(n_29),
.B2(n_16),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_102),
.A2(n_7),
.B1(n_8),
.B2(n_108),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_52),
.B(n_22),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_103),
.B(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_40),
.C(n_33),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_51),
.C(n_66),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_35),
.B1(n_16),
.B2(n_29),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_SL g160 ( 
.A(n_108),
.B(n_111),
.C(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_45),
.B(n_34),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_121),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_82),
.B(n_32),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_27),
.B1(n_25),
.B2(n_33),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_27),
.B1(n_31),
.B2(n_12),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_55),
.B(n_31),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_11),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_130),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_62),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_133),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_47),
.B(n_1),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_2),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_134),
.B(n_147),
.Y(n_214)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_98),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_135),
.Y(n_196)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_137),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_93),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_139),
.A2(n_101),
.B(n_115),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_140),
.B(n_120),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_97),
.A2(n_81),
.B1(n_65),
.B2(n_53),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_141),
.A2(n_143),
.B1(n_146),
.B2(n_169),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_108),
.A2(n_77),
.B1(n_4),
.B2(n_6),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_167),
.B1(n_178),
.B2(n_114),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_97),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_8),
.B1(n_111),
.B2(n_86),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_166),
.B1(n_117),
.B2(n_104),
.Y(n_184)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_123),
.Y(n_154)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_155),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_8),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_164),
.Y(n_193)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_160),
.B(n_88),
.Y(n_201)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_91),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_165),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_110),
.B1(n_91),
.B2(n_92),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_133),
.B1(n_131),
.B2(n_121),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_130),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_152),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

BUFx24_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_94),
.B(n_103),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_175),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g175 ( 
.A(n_107),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_105),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_177),
.Y(n_209)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_129),
.A2(n_85),
.B1(n_127),
.B2(n_88),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_150),
.Y(n_212)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_180),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_113),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_183),
.B(n_192),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_184),
.B(n_189),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_167),
.A2(n_117),
.B1(n_114),
.B2(n_120),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_152),
.B1(n_136),
.B2(n_149),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_174),
.B(n_132),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_200),
.B(n_181),
.Y(n_253)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_201),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_161),
.A2(n_85),
.B1(n_129),
.B2(n_107),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_135),
.B1(n_148),
.B2(n_159),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_180),
.A2(n_88),
.B1(n_127),
.B2(n_128),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_140),
.B(n_123),
.C(n_115),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_158),
.C(n_170),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_157),
.B(n_101),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_217),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_211),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_157),
.B(n_136),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_146),
.B(n_171),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_138),
.A2(n_168),
.B1(n_177),
.B2(n_163),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_221),
.Y(n_263)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_222),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_223),
.A2(n_224),
.B1(n_230),
.B2(n_243),
.Y(n_269)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_198),
.Y(n_225)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_185),
.Y(n_227)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_227),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_229),
.A2(n_231),
.B1(n_247),
.B2(n_196),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_234),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_172),
.B1(n_153),
.B2(n_154),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_237),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_155),
.B(n_137),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_196),
.B(n_187),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_253),
.C(n_205),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_200),
.B(n_176),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_244),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_175),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_214),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_246),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_216),
.A3(n_186),
.B1(n_201),
.B2(n_192),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_181),
.A2(n_216),
.B1(n_202),
.B2(n_208),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_252),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_197),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_191),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_183),
.B(n_175),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_193),
.B(n_199),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_182),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_194),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_255),
.B(n_228),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_215),
.B(n_188),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_256),
.B(n_270),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_257),
.A2(n_246),
.B1(n_222),
.B2(n_221),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_260),
.B(n_244),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_220),
.B(n_191),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_213),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_265),
.B(n_266),
.C(n_276),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_213),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_283),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_269),
.B(n_271),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_205),
.B(n_198),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_190),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_229),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_226),
.B(n_190),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_236),
.A2(n_182),
.B1(n_249),
.B2(n_235),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_238),
.B1(n_250),
.B2(n_240),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_182),
.C(n_242),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_280),
.B(n_251),
.C(n_237),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_282),
.B(n_227),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_226),
.B(n_182),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_252),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_245),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_268),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_292),
.Y(n_318)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_287),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_291),
.B(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_263),
.Y(n_290)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_290),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_282),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_223),
.Y(n_293)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_293),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_247),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_264),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_265),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_309),
.C(n_280),
.Y(n_312)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_304),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_233),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_273),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_307),
.B1(n_308),
.B2(n_279),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_255),
.B(n_254),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_312),
.B(n_316),
.C(n_320),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_284),
.C(n_278),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_324),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_276),
.C(n_266),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_298),
.B(n_251),
.C(n_269),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_298),
.B(n_251),
.C(n_279),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_323),
.B(n_327),
.C(n_328),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_262),
.B1(n_278),
.B2(n_257),
.Y(n_325)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_281),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_303),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_258),
.C(n_281),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_256),
.C(n_274),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_302),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_329),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_308),
.Y(n_332)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_332),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_293),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_333),
.B(n_335),
.C(n_341),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_267),
.B1(n_270),
.B2(n_288),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_334),
.A2(n_337),
.B(n_317),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_318),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_336),
.B(n_304),
.Y(n_360)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_297),
.B(n_292),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_297),
.B(n_274),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_259),
.B(n_260),
.C(n_317),
.Y(n_354)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_340),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_300),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_310),
.A2(n_294),
.B1(n_291),
.B2(n_289),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_342),
.A2(n_319),
.B1(n_321),
.B2(n_291),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_323),
.B(n_289),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_343),
.A2(n_315),
.B1(n_286),
.B2(n_290),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_307),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_314),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_305),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_347),
.B(n_326),
.C(n_328),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_349),
.B(n_355),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_351),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_352),
.A2(n_348),
.B1(n_343),
.B2(n_341),
.Y(n_368)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_320),
.C(n_311),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_358),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_261),
.C(n_301),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_361),
.Y(n_372)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_360),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_348),
.B(n_261),
.C(n_295),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_350),
.A2(n_344),
.B1(n_339),
.B2(n_338),
.Y(n_362)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_360),
.A2(n_346),
.B1(n_342),
.B2(n_296),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_370),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_272),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_353),
.A2(n_335),
.B1(n_333),
.B2(n_231),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_369),
.B(n_351),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_361),
.A2(n_275),
.B1(n_272),
.B2(n_232),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_377),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_357),
.B(n_354),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_SL g385 ( 
.A(n_375),
.B(n_369),
.C(n_371),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_345),
.Y(n_376)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_376),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_367),
.B(n_357),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_367),
.B(n_275),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_379),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_225),
.C(n_368),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_370),
.Y(n_384)
);

AOI21xp33_ASAP7_75t_L g383 ( 
.A1(n_374),
.A2(n_364),
.B(n_371),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_383),
.A2(n_373),
.B(n_381),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_385),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_380),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_388),
.B(n_390),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_379),
.Y(n_390)
);

AO21x2_ASAP7_75t_L g392 ( 
.A1(n_391),
.A2(n_384),
.B(n_372),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_392),
.A2(n_389),
.B(n_387),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_393),
.Y(n_395)
);


endmodule