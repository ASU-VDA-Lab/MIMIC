module fake_jpeg_29352_n_519 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_52),
.B(n_75),
.Y(n_148)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_62),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_64),
.Y(n_106)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_37),
.B(n_15),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_42),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_13),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_81),
.B(n_91),
.Y(n_151)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_84),
.Y(n_147)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_20),
.B(n_13),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_32),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_47),
.Y(n_135)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_96),
.Y(n_110)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

BUFx4f_ASAP7_75t_SL g98 ( 
.A(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_40),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_49),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_99),
.B(n_46),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_13),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_45),
.Y(n_137)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_31),
.B1(n_38),
.B2(n_47),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_102),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_68),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_111),
.B(n_117),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_74),
.B(n_36),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_68),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_143),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_125),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_53),
.B(n_36),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_129),
.B(n_137),
.Y(n_169)
);

BUFx12_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

BUFx4f_ASAP7_75t_SL g199 ( 
.A(n_132),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_135),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_55),
.Y(n_139)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_139),
.Y(n_189)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_57),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g194 ( 
.A(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_96),
.Y(n_143)
);

HAxp5_ASAP7_75t_SL g145 ( 
.A(n_88),
.B(n_22),
.CON(n_145),
.SN(n_145)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_26),
.B(n_18),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_58),
.B(n_28),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_155),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_28),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_54),
.B(n_46),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_159),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_92),
.A2(n_12),
.B(n_1),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_145),
.A2(n_61),
.B1(n_94),
.B2(n_69),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_163),
.A2(n_174),
.B1(n_195),
.B2(n_207),
.Y(n_237)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_164),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_168),
.B(n_203),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_153),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g258 ( 
.A(n_170),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_18),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_176),
.Y(n_235)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g229 ( 
.A(n_172),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_107),
.A2(n_73),
.B1(n_90),
.B2(n_89),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_137),
.B(n_45),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_183),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_44),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_213),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_122),
.A2(n_93),
.B1(n_51),
.B2(n_70),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_103),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_121),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_188),
.B(n_198),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_122),
.A2(n_51),
.B1(n_26),
.B2(n_43),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_130),
.A2(n_43),
.B1(n_44),
.B2(n_38),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_191),
.A2(n_214),
.B1(n_106),
.B2(n_140),
.Y(n_241)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_193),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_196),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_124),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_216),
.Y(n_228)
);

NOR2x1_ASAP7_75t_L g198 ( 
.A(n_135),
.B(n_29),
.Y(n_198)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_133),
.A2(n_97),
.B1(n_31),
.B2(n_40),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_206),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_134),
.A2(n_86),
.B1(n_79),
.B2(n_47),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_154),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_106),
.Y(n_244)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx8_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_113),
.B(n_41),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_210),
.B(n_211),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_113),
.B(n_41),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_41),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_130),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_103),
.Y(n_215)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_140),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_219),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_218),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_152),
.B(n_150),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_220),
.B(n_223),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_179),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_110),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_242),
.C(n_166),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_244),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_184),
.B(n_152),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_182),
.A2(n_134),
.B1(n_136),
.B2(n_161),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_245),
.A2(n_255),
.B1(n_209),
.B2(n_200),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_136),
.B1(n_160),
.B2(n_118),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_247),
.A2(n_254),
.B1(n_263),
.B2(n_218),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_169),
.B(n_132),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_193),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_161),
.B1(n_160),
.B2(n_127),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_L g255 ( 
.A1(n_187),
.A2(n_127),
.B1(n_138),
.B2(n_162),
.Y(n_255)
);

OAI21xp33_ASAP7_75t_L g257 ( 
.A1(n_175),
.A2(n_40),
.B(n_35),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_189),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_194),
.A2(n_138),
.B1(n_119),
.B2(n_123),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_198),
.Y(n_281)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_185),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_269),
.B(n_273),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_237),
.A2(n_194),
.B1(n_164),
.B2(n_181),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_270),
.A2(n_304),
.B1(n_308),
.B2(n_264),
.Y(n_313)
);

BUFx4f_ASAP7_75t_SL g271 ( 
.A(n_258),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_271),
.Y(n_345)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_231),
.A2(n_226),
.B1(n_250),
.B2(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_272),
.A2(n_115),
.B1(n_202),
.B2(n_189),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_262),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_213),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_292),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_276),
.B(n_286),
.Y(n_325)
);

INVx13_ASAP7_75t_L g277 ( 
.A(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_287),
.Y(n_317)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_279),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_203),
.B1(n_208),
.B2(n_192),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_280),
.B(n_301),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_281),
.B(n_282),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_228),
.B(n_259),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_283),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_242),
.B(n_166),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_284),
.B(n_289),
.C(n_226),
.Y(n_312)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_224),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_293),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_251),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_231),
.A2(n_215),
.B1(n_216),
.B2(n_173),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_290),
.A2(n_299),
.B(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_239),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_291),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_250),
.B(n_204),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_267),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_238),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_294),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_295),
.A2(n_261),
.B1(n_280),
.B2(n_308),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_235),
.B(n_170),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_296),
.B(n_297),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_243),
.B(n_170),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_224),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_298),
.Y(n_314)
);

AND2x6_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_199),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_302),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g301 ( 
.A1(n_245),
.A2(n_183),
.B1(n_172),
.B2(n_142),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_260),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_305),
.Y(n_326)
);

INVx13_ASAP7_75t_L g304 ( 
.A(n_258),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_257),
.B(n_199),
.CI(n_132),
.CON(n_305),
.SN(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_306),
.B(n_309),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_232),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_253),
.B(n_196),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_35),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_323),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_301),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_221),
.C(n_264),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_320),
.C(n_321),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_300),
.A2(n_261),
.B1(n_236),
.B2(n_123),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_319),
.A2(n_336),
.B1(n_342),
.B2(n_348),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_249),
.C(n_222),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_249),
.C(n_246),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_199),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_275),
.B(n_246),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_329),
.B(n_335),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_236),
.C(n_240),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_330),
.B(n_331),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_256),
.C(n_266),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g332 ( 
.A1(n_306),
.A2(n_266),
.B1(n_232),
.B2(n_119),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_332),
.A2(n_309),
.B1(n_293),
.B2(n_310),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_229),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_256),
.C(n_178),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_337),
.B(n_304),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_229),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_344),
.Y(n_362)
);

OA22x2_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_301),
.B1(n_280),
.B2(n_342),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_295),
.A2(n_115),
.B1(n_212),
.B2(n_35),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_299),
.A2(n_25),
.B1(n_12),
.B2(n_3),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_350),
.A2(n_357),
.B1(n_368),
.B2(n_372),
.Y(n_411)
);

BUFx12_ASAP7_75t_L g351 ( 
.A(n_345),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_356),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_353),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_5),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_305),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

INVx13_ASAP7_75t_L g356 ( 
.A(n_345),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_316),
.A2(n_330),
.B1(n_326),
.B2(n_331),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_271),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_363),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_305),
.Y(n_364)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_364),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_271),
.Y(n_365)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_365),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_314),
.B(n_302),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_366),
.B(n_375),
.Y(n_387)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_347),
.Y(n_367)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_326),
.A2(n_328),
.B1(n_312),
.B2(n_343),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_327),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_369),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_307),
.Y(n_370)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_370),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_328),
.A2(n_307),
.B1(n_280),
.B2(n_301),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_371),
.A2(n_311),
.B1(n_7),
.B2(n_8),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_343),
.A2(n_318),
.B1(n_341),
.B2(n_315),
.Y(n_372)
);

CKINVDCx10_ASAP7_75t_R g373 ( 
.A(n_317),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_373),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_318),
.A2(n_294),
.B1(n_279),
.B2(n_287),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_377),
.Y(n_392)
);

CKINVDCx12_ASAP7_75t_R g376 ( 
.A(n_322),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_376),
.B(n_381),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_334),
.A2(n_277),
.B1(n_1),
.B2(n_3),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_340),
.B(n_0),
.Y(n_378)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_378),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_0),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_380),
.Y(n_393)
);

INVx13_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_333),
.B(n_0),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_321),
.B(n_4),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_382),
.B(n_5),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_364),
.A2(n_334),
.B(n_335),
.C(n_348),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_383),
.A2(n_395),
.B(n_362),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_352),
.B(n_325),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_384),
.B(n_408),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_369),
.B(n_349),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_388),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_325),
.C(n_323),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_394),
.C(n_396),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_337),
.C(n_319),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_355),
.A2(n_339),
.B(n_324),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_346),
.C(n_311),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_397),
.B(n_11),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_401),
.A2(n_404),
.B1(n_350),
.B2(n_374),
.Y(n_426)
);

AO21x1_ASAP7_75t_L g427 ( 
.A1(n_403),
.A2(n_354),
.B(n_356),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_361),
.B(n_8),
.C(n_9),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_378),
.C(n_379),
.Y(n_436)
);

NOR4xp25_ASAP7_75t_L g407 ( 
.A(n_370),
.B(n_8),
.C(n_9),
.D(n_10),
.Y(n_407)
);

AOI21xp33_ASAP7_75t_L g420 ( 
.A1(n_407),
.A2(n_377),
.B(n_365),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_368),
.B(n_361),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_358),
.A2(n_9),
.B1(n_11),
.B2(n_376),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_410),
.A2(n_358),
.B1(n_373),
.B2(n_367),
.Y(n_417)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_414),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_415),
.Y(n_448)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_400),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_417),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_406),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_420),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_411),
.A2(n_355),
.B1(n_371),
.B2(n_362),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_437),
.B1(n_403),
.B2(n_401),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_403),
.C(n_385),
.Y(n_441)
);

INVx13_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_428),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_391),
.A2(n_388),
.B1(n_398),
.B2(n_386),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_425),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_426),
.A2(n_427),
.B1(n_392),
.B2(n_409),
.Y(n_442)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_351),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_430),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_386),
.A2(n_354),
.B1(n_360),
.B2(n_372),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_384),
.B(n_357),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_433),
.Y(n_443)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_432),
.A2(n_11),
.B(n_434),
.Y(n_457)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_434),
.A2(n_435),
.B(n_407),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_385),
.A2(n_354),
.B(n_351),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_396),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_411),
.A2(n_382),
.B1(n_351),
.B2(n_380),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_424),
.B(n_408),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_438),
.B(n_454),
.C(n_455),
.Y(n_460)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_441),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_442),
.A2(n_449),
.B1(n_435),
.B2(n_432),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_446),
.A2(n_450),
.B1(n_451),
.B2(n_426),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_428),
.A2(n_392),
.B1(n_409),
.B2(n_389),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_419),
.A2(n_389),
.B1(n_383),
.B2(n_412),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_437),
.A2(n_412),
.B1(n_387),
.B2(n_394),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_452),
.B(n_431),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_413),
.B(n_390),
.C(n_405),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_413),
.B(n_399),
.C(n_397),
.Y(n_455)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_456),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_457),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_422),
.Y(n_458)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_459),
.A2(n_468),
.B1(n_444),
.B2(n_453),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_445),
.B(n_415),
.Y(n_461)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_467),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_440),
.A2(n_415),
.B(n_427),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_443),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_448),
.Y(n_466)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_466),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_418),
.Y(n_467)
);

A2O1A1Ixp33_ASAP7_75t_SL g468 ( 
.A1(n_441),
.A2(n_427),
.B(n_421),
.C(n_423),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_424),
.C(n_436),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_471),
.C(n_443),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_414),
.C(n_416),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_446),
.A2(n_433),
.B1(n_450),
.B2(n_439),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_449),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_480),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_470),
.A2(n_451),
.B1(n_455),
.B2(n_442),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_479),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_481),
.B(n_483),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_464),
.A2(n_438),
.B1(n_459),
.B2(n_467),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_482),
.B(n_472),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_460),
.C(n_469),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_473),
.B(n_465),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_463),
.Y(n_492)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_466),
.Y(n_487)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_487),
.Y(n_493)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_489),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_461),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_491),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_494),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_460),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g495 ( 
.A(n_480),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_495),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_474),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_496),
.A2(n_497),
.B1(n_485),
.B2(n_478),
.Y(n_505)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_487),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_488),
.A2(n_485),
.B(n_476),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_505),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_481),
.C(n_484),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_503),
.B(n_490),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_509),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_490),
.C(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_508),
.B(n_499),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

AO21x1_ASAP7_75t_L g510 ( 
.A1(n_506),
.A2(n_504),
.B(n_458),
.Y(n_510)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_510),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_493),
.C(n_500),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_513),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_515),
.A2(n_511),
.B(n_514),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_502),
.C(n_486),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_517),
.B(n_468),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_468),
.B(n_512),
.Y(n_519)
);


endmodule