module fake_aes_11124_n_38 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_38);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_30;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_13), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_3), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_12), .B(n_8), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_3), .Y(n_20) );
BUFx6f_ASAP7_75t_L g21 ( .A(n_10), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_16), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_17), .B(n_1), .Y(n_23) );
OR2x6_ASAP7_75t_L g24 ( .A(n_20), .B(n_1), .Y(n_24) );
OAI21x1_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_19), .B(n_21), .Y(n_25) );
OAI21x1_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_19), .B(n_21), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_24), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_27), .B(n_24), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_24), .Y(n_29) );
OAI22xp33_ASAP7_75t_SL g30 ( .A1(n_28), .A2(n_18), .B1(n_15), .B2(n_27), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_25), .Y(n_31) );
INVxp33_ASAP7_75t_SL g32 ( .A(n_30), .Y(n_32) );
NOR2x1p5_ASAP7_75t_L g33 ( .A(n_32), .B(n_21), .Y(n_33) );
NAND2x1p5_ASAP7_75t_L g34 ( .A(n_31), .B(n_26), .Y(n_34) );
AOI21xp33_ASAP7_75t_SL g35 ( .A1(n_33), .A2(n_2), .B(n_4), .Y(n_35) );
OAI22xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_21), .B1(n_4), .B2(n_5), .Y(n_36) );
OAI22xp5_ASAP7_75t_SL g37 ( .A1(n_35), .A2(n_2), .B1(n_5), .B2(n_6), .Y(n_37) );
AOI322xp5_ASAP7_75t_L g38 ( .A1(n_37), .A2(n_36), .A3(n_7), .B1(n_6), .B2(n_11), .C1(n_14), .C2(n_9), .Y(n_38) );
endmodule