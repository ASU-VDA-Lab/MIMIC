module fake_netlist_6_3625_n_1704 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1704);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1704;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_50),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_80),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_28),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_37),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_26),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_148),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_136),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_44),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_19),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_39),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_104),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_90),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_71),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_132),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_20),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_53),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_54),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_147),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_55),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_96),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_6),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_114),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_87),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_156),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_24),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_3),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_56),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_119),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_146),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_57),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_64),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_43),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_125),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_133),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_45),
.Y(n_208)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_15),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_52),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_41),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_29),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_112),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_101),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_45),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_19),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_40),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_43),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_83),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_102),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_62),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_91),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_128),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_68),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_95),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_11),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_86),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_23),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_109),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_137),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_14),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_34),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_0),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_145),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_108),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_22),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_49),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_127),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_32),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_69),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_44),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_100),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_92),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_124),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_99),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_52),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_78),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_8),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_110),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_53),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_22),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_7),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_70),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_140),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_31),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_41),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_39),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_113),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_105),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_89),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_73),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_115),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_40),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_135),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_20),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_93),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_111),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_37),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_131),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_141),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_46),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_154),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_3),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_106),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_18),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_7),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_13),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_2),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_28),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_27),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_6),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_122),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_50),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_151),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_107),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_26),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_34),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_130),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_65),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g304 ( 
.A(n_84),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_67),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_9),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_116),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_35),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_63),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_38),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_117),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_207),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_251),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_255),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_209),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_209),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_191),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_209),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_253),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_209),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_209),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_254),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_209),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_209),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_209),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_181),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_181),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_181),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_181),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_181),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_239),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_289),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_198),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_218),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_218),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_218),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_241),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_289),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_241),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_218),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_162),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_187),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_164),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_188),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_162),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_190),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_192),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_300),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_234),
.Y(n_360)
);

BUFx5_ASAP7_75t_L g361 ( 
.A(n_158),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_170),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_241),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_235),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_205),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_270),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_164),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_235),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_182),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_252),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_195),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_215),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_208),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_259),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_270),
.Y(n_377)
);

INVxp33_ASAP7_75t_SL g378 ( 
.A(n_168),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_211),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_197),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_260),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_200),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_263),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g384 ( 
.A(n_215),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_274),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_281),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_284),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_286),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_212),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_324),
.A2(n_193),
.B1(n_310),
.B2(n_175),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_350),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_334),
.B(n_225),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_323),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_323),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_352),
.Y(n_395)
);

OAI21x1_ASAP7_75t_L g396 ( 
.A1(n_317),
.A2(n_219),
.B(n_179),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_318),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_374),
.B(n_173),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_265),
.C(n_161),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_334),
.B(n_225),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_173),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_314),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_325),
.Y(n_410)
);

INVx6_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_355),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_245),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_316),
.A2(n_168),
.B1(n_312),
.B2(n_175),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_354),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_325),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_341),
.B(n_233),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_351),
.B(n_245),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_316),
.A2(n_169),
.B1(n_312),
.B2(n_176),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_357),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_330),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_330),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_319),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_347),
.B(n_249),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_326),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_326),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_327),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_319),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_331),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_332),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_332),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_L g436 ( 
.A(n_336),
.B(n_169),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_335),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_315),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_373),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_337),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_337),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_369),
.B(n_163),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_176),
.B1(n_244),
.B2(n_294),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_338),
.Y(n_445)
);

OA21x2_ASAP7_75t_L g446 ( 
.A1(n_339),
.A2(n_219),
.B(n_179),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_341),
.B(n_233),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_321),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_384),
.B(n_163),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_346),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_368),
.A2(n_301),
.B1(n_297),
.B2(n_305),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_346),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_349),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_336),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_349),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_348),
.Y(n_457)
);

AND2x6_ASAP7_75t_L g458 ( 
.A(n_353),
.B(n_160),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_425),
.B(n_333),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_424),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_443),
.B(n_380),
.Y(n_461)
);

INVx5_ASAP7_75t_L g462 ( 
.A(n_458),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_390),
.B(n_382),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_416),
.A2(n_389),
.B1(n_379),
.B2(n_375),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_391),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_419),
.A2(n_354),
.B1(n_343),
.B2(n_293),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_358),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_359),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_304),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_433),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_392),
.B(n_264),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_399),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_392),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_399),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_411),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_450),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_392),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_455),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_393),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_356),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_394),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_403),
.B(n_377),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_405),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_444),
.A2(n_230),
.B1(n_213),
.B2(n_216),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_433),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_402),
.A2(n_364),
.B1(n_342),
.B2(n_372),
.Y(n_496)
);

INVxp67_ASAP7_75t_SL g497 ( 
.A(n_401),
.Y(n_497)
);

NAND3xp33_ASAP7_75t_L g498 ( 
.A(n_402),
.B(n_363),
.C(n_362),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_392),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_435),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_404),
.A2(n_295),
.B1(n_264),
.B2(n_361),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_401),
.B(n_361),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_455),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_435),
.Y(n_506)
);

AOI21x1_ASAP7_75t_L g507 ( 
.A1(n_446),
.A2(n_166),
.B(n_159),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_440),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_433),
.Y(n_510)
);

INVx8_ASAP7_75t_L g511 ( 
.A(n_458),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_401),
.B(n_361),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_431),
.B(n_356),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_444),
.A2(n_236),
.B1(n_308),
.B2(n_307),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_440),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_440),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g518 ( 
.A(n_406),
.B(n_381),
.C(n_376),
.Y(n_518)
);

CKINVDCx16_ASAP7_75t_R g519 ( 
.A(n_390),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_404),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_453),
.Y(n_521)
);

INVx8_ASAP7_75t_L g522 ( 
.A(n_458),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_404),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_401),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_434),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_404),
.A2(n_418),
.B1(n_447),
.B2(n_427),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_406),
.B(n_167),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_415),
.B(n_367),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_415),
.B(n_367),
.Y(n_530)
);

CKINVDCx6p67_ASAP7_75t_R g531 ( 
.A(n_407),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_405),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_409),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_418),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_410),
.B(n_361),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_418),
.B(n_360),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_420),
.B(n_375),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_409),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_420),
.B(n_379),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_R g541 ( 
.A(n_412),
.B(n_389),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_418),
.B(n_360),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_409),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_452),
.B(n_270),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_417),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_417),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_438),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_417),
.Y(n_549)
);

INVx4_ASAP7_75t_L g550 ( 
.A(n_411),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_L g552 ( 
.A1(n_413),
.A2(n_238),
.B1(n_217),
.B2(n_220),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_410),
.B(n_427),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_429),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_447),
.B(n_165),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_421),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_410),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_447),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_410),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_447),
.B(n_165),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_397),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_413),
.B(n_344),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_397),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_400),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_400),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_427),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_458),
.B(n_160),
.Y(n_572)
);

AOI21x1_ASAP7_75t_L g573 ( 
.A1(n_446),
.A2(n_194),
.B(n_189),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_434),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_408),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_427),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_428),
.B(n_361),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_428),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_428),
.B(n_361),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_408),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_449),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_434),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_414),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_428),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_414),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_430),
.B(n_361),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_430),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_430),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_430),
.B(n_422),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_422),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_446),
.A2(n_388),
.B1(n_383),
.B2(n_385),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_457),
.B(n_171),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_434),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_423),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_423),
.B(n_201),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_426),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_426),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_457),
.B(n_345),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_432),
.B(n_171),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_437),
.B(n_172),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_437),
.B(n_386),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_441),
.B(n_172),
.Y(n_605)
);

OAI21xp33_ASAP7_75t_SL g606 ( 
.A1(n_441),
.A2(n_371),
.B(n_370),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_442),
.B(n_202),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_R g608 ( 
.A(n_442),
.B(n_204),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_482),
.B(n_445),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_482),
.A2(n_446),
.B1(n_160),
.B2(n_183),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_461),
.B(n_177),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_537),
.A2(n_183),
.B1(n_160),
.B2(n_313),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_459),
.B(n_177),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_540),
.B(n_467),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_585),
.B(n_445),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_481),
.A2(n_456),
.B(n_448),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_530),
.A2(n_301),
.B1(n_297),
.B2(n_305),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_473),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_585),
.B(n_448),
.Y(n_621)
);

BUFx8_ASAP7_75t_L g622 ( 
.A(n_516),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

NOR3xp33_ASAP7_75t_L g624 ( 
.A(n_466),
.B(n_371),
.C(n_242),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_542),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_469),
.B(n_456),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_451),
.Y(n_627)
);

BUFx5_ASAP7_75t_L g628 ( 
.A(n_561),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_479),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_478),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_481),
.B(n_160),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_485),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_485),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_481),
.B(n_183),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_499),
.B(n_451),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_499),
.B(n_451),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_478),
.B(n_386),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_483),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_487),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_481),
.B(n_183),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_487),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_474),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_387),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_520),
.B(n_451),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_486),
.B(n_178),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_520),
.A2(n_226),
.B1(n_206),
.B2(n_210),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_463),
.A2(n_183),
.B1(n_313),
.B2(n_227),
.Y(n_647)
);

NOR2xp67_ASAP7_75t_L g648 ( 
.A(n_513),
.B(n_223),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_491),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_463),
.A2(n_313),
.B1(n_268),
.B2(n_196),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_523),
.A2(n_534),
.B1(n_562),
.B2(n_471),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_550),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_463),
.A2(n_477),
.B1(n_471),
.B2(n_528),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_491),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_523),
.B(n_451),
.Y(n_655)
);

BUFx5_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_527),
.A2(n_229),
.B1(n_203),
.B2(n_214),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_484),
.B(n_387),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_566),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_582),
.B(n_221),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_550),
.B(n_463),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_550),
.B(n_313),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_529),
.B(n_530),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_483),
.B(n_365),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_550),
.B(n_313),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_534),
.B(n_451),
.Y(n_666)
);

NAND2x1p5_ASAP7_75t_L g667 ( 
.A(n_562),
.B(n_222),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_497),
.B(n_454),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_484),
.B(n_365),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_524),
.B(n_567),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_463),
.B(n_224),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_492),
.Y(n_672)
);

AO22x2_ASAP7_75t_L g673 ( 
.A1(n_544),
.A2(n_476),
.B1(n_488),
.B2(n_474),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

NOR2xp67_ASAP7_75t_L g675 ( 
.A(n_498),
.B(n_231),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_536),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_492),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_477),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_591),
.B(n_595),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_546),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_591),
.B(n_454),
.Y(n_681)
);

CKINVDCx14_ASAP7_75t_R g682 ( 
.A(n_531),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_471),
.A2(n_273),
.B1(n_232),
.B2(n_240),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_471),
.A2(n_276),
.B1(n_247),
.B2(n_248),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_474),
.Y(n_685)
);

NOR3xp33_ASAP7_75t_L g686 ( 
.A(n_496),
.B(n_228),
.C(n_290),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_536),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_477),
.B(n_237),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_595),
.B(n_454),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_471),
.B(n_494),
.Y(n_690)
);

INVxp33_ASAP7_75t_L g691 ( 
.A(n_505),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_546),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_505),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_599),
.B(n_454),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_600),
.Y(n_695)
);

BUFx5_ASAP7_75t_L g696 ( 
.A(n_563),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_599),
.B(n_454),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_600),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_528),
.A2(n_279),
.B1(n_296),
.B2(n_258),
.Y(n_699)
);

INVx5_ASAP7_75t_L g700 ( 
.A(n_597),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_496),
.B(n_178),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_563),
.B(n_454),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_571),
.B(n_411),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_571),
.B(n_411),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_576),
.B(n_578),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_477),
.B(n_243),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_460),
.B(n_366),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_596),
.B(n_180),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_576),
.B(n_411),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_604),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_607),
.B(n_180),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_578),
.B(n_588),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_588),
.B(n_250),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_R g714 ( 
.A(n_541),
.B(n_184),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_477),
.A2(n_528),
.B1(n_592),
.B2(n_575),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_516),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_589),
.B(n_256),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_555),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_589),
.B(n_303),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_554),
.B(n_311),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_590),
.B(n_261),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_566),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_601),
.B(n_269),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_559),
.Y(n_724)
);

INVx2_ASAP7_75t_SL g725 ( 
.A(n_460),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_568),
.B(n_271),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_568),
.B(n_272),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_557),
.B(n_184),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_559),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_569),
.B(n_278),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_460),
.Y(n_731)
);

NAND3xp33_ASAP7_75t_L g732 ( 
.A(n_468),
.B(n_292),
.C(n_277),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_528),
.A2(n_287),
.B1(n_282),
.B2(n_283),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_597),
.B(n_285),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_597),
.B(n_185),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_L g736 ( 
.A(n_501),
.B(n_185),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_604),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_528),
.A2(n_294),
.B1(n_244),
.B2(n_307),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_569),
.B(n_186),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_570),
.B(n_186),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_597),
.B(n_298),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_564),
.B(n_309),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_460),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_570),
.B(n_298),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_575),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_581),
.B(n_584),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_548),
.A2(n_366),
.B1(n_370),
.B2(n_8),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_584),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_560),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_603),
.B(n_288),
.C(n_246),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_531),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_586),
.B(n_309),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_560),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_586),
.B(n_299),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_598),
.B(n_299),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_552),
.B(n_302),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_598),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_605),
.B(n_593),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_462),
.B(n_602),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_602),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_519),
.B(n_267),
.C(n_257),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_608),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_462),
.B(n_302),
.Y(n_764)
);

BUFx3_ASAP7_75t_L g765 ( 
.A(n_467),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_565),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_465),
.B(n_306),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_465),
.B(n_306),
.Y(n_768)
);

NAND2x1p5_ASAP7_75t_L g769 ( 
.A(n_462),
.B(n_98),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_565),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_579),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_SL g772 ( 
.A(n_558),
.B(n_308),
.Y(n_772)
);

NAND3xp33_ASAP7_75t_L g773 ( 
.A(n_514),
.B(n_291),
.C(n_275),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_475),
.B(n_458),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_514),
.B(n_266),
.Y(n_775)
);

AOI22xp5_ASAP7_75t_L g776 ( 
.A1(n_498),
.A2(n_458),
.B1(n_262),
.B2(n_236),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_500),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_678),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_716),
.B(n_511),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_670),
.B(n_475),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_678),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_690),
.A2(n_757),
.B1(n_663),
.B2(n_611),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_658),
.B(n_558),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_678),
.B(n_480),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_669),
.B(n_707),
.Y(n_785)
);

OR2x2_ASAP7_75t_SL g786 ( 
.A(n_773),
.B(n_519),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_611),
.A2(n_606),
.B1(n_533),
.B2(n_532),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_693),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_710),
.B(n_518),
.Y(n_789)
);

AO22x1_ASAP7_75t_L g790 ( 
.A1(n_690),
.A2(n_464),
.B1(n_606),
.B2(n_458),
.Y(n_790)
);

AO22x1_ASAP7_75t_L g791 ( 
.A1(n_663),
.A2(n_775),
.B1(n_757),
.B2(n_645),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_678),
.B(n_480),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_676),
.Y(n_793)
);

CKINVDCx16_ASAP7_75t_R g794 ( 
.A(n_682),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_645),
.A2(n_543),
.B1(n_532),
.B2(n_533),
.Y(n_795)
);

A2O1A1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_613),
.A2(n_518),
.B(n_587),
.C(n_512),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_612),
.A2(n_553),
.B1(n_539),
.B2(n_543),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_679),
.B(n_489),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_759),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_659),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_659),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_715),
.B(n_489),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_745),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_745),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_SL g805 ( 
.A(n_613),
.B(n_580),
.C(n_503),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_643),
.Y(n_806)
);

OR2x6_ASAP7_75t_L g807 ( 
.A(n_716),
.B(n_511),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_765),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_715),
.B(n_490),
.Y(n_809)
);

HB1xp67_ASAP7_75t_L g810 ( 
.A(n_643),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_687),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_691),
.B(n_464),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_691),
.B(n_490),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_664),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_674),
.Y(n_815)
);

NOR3xp33_ASAP7_75t_SL g816 ( 
.A(n_617),
.B(n_535),
.C(n_577),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_626),
.B(n_610),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_682),
.Y(n_818)
);

CKINVDCx11_ASAP7_75t_R g819 ( 
.A(n_752),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_763),
.B(n_462),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_661),
.A2(n_522),
.B(n_511),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_737),
.B(n_472),
.Y(n_822)
);

CKINVDCx14_ASAP7_75t_R g823 ( 
.A(n_714),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_708),
.B(n_462),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_610),
.B(n_695),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_661),
.A2(n_522),
.B(n_511),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_643),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_759),
.A2(n_549),
.B1(n_539),
.B2(n_547),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_664),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_637),
.Y(n_830)
);

NOR2x1_ASAP7_75t_L g831 ( 
.A(n_765),
.B(n_472),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_612),
.A2(n_556),
.B1(n_509),
.B2(n_502),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_674),
.B(n_698),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_708),
.B(n_462),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_L g835 ( 
.A(n_700),
.B(n_511),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_622),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_653),
.A2(n_507),
.B1(n_573),
.B2(n_556),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_614),
.B(n_502),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_623),
.B(n_506),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_SL g840 ( 
.A1(n_738),
.A2(n_2),
.B1(n_5),
.B2(n_10),
.Y(n_840)
);

NAND2x1p5_ASAP7_75t_L g841 ( 
.A(n_700),
.B(n_652),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_738),
.B(n_772),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_625),
.B(n_506),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_637),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_722),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_722),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_609),
.B(n_521),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_622),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_657),
.A2(n_521),
.B1(n_509),
.B2(n_515),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_615),
.B(n_538),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_515),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_621),
.B(n_628),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_642),
.A2(n_472),
.B1(n_493),
.B2(n_574),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_748),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_660),
.Y(n_855)
);

OR2x6_ASAP7_75t_L g856 ( 
.A(n_752),
.B(n_522),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_628),
.B(n_525),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_777),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_660),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_660),
.Y(n_860)
);

AND2x6_ASAP7_75t_SL g861 ( 
.A(n_701),
.B(n_12),
.Y(n_861)
);

AO22x1_ASAP7_75t_L g862 ( 
.A1(n_762),
.A2(n_493),
.B1(n_495),
.B2(n_504),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_711),
.B(n_594),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_749),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_628),
.B(n_525),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_685),
.B(n_493),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_628),
.B(n_517),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_777),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_628),
.B(n_517),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_628),
.B(n_656),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_656),
.B(n_538),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_761),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_746),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_711),
.A2(n_495),
.B1(n_504),
.B2(n_574),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_630),
.B(n_495),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_705),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_712),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_656),
.B(n_504),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_755),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_771),
.B(n_12),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_656),
.B(n_545),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_651),
.A2(n_545),
.B1(n_508),
.B2(n_574),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_725),
.Y(n_884)
);

INVxp33_ASAP7_75t_SL g885 ( 
.A(n_683),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_638),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_618),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_769),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_724),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_656),
.B(n_508),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_731),
.B(n_743),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_751),
.B(n_545),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_671),
.A2(n_572),
.B(n_508),
.C(n_510),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_648),
.B(n_594),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_619),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_747),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_624),
.B(n_510),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_700),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_620),
.Y(n_899)
);

AND2x6_ASAP7_75t_L g900 ( 
.A(n_774),
.B(n_594),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_656),
.B(n_510),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_755),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_747),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_696),
.B(n_594),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_769),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_667),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_700),
.B(n_594),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_728),
.B(n_583),
.Y(n_908)
);

INVx1_ASAP7_75t_SL g909 ( 
.A(n_756),
.Y(n_909)
);

AND2x2_ASAP7_75t_SL g910 ( 
.A(n_653),
.B(n_583),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_723),
.B(n_583),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_729),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_629),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_686),
.A2(n_522),
.B1(n_551),
.B2(n_526),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_673),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_736),
.A2(n_701),
.B1(n_742),
.B2(n_728),
.Y(n_916)
);

AND2x2_ASAP7_75t_SL g917 ( 
.A(n_742),
.B(n_583),
.Y(n_917)
);

BUFx8_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_652),
.B(n_583),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_673),
.B(n_573),
.Y(n_920)
);

AO21x1_ASAP7_75t_L g921 ( 
.A1(n_671),
.A2(n_507),
.B(n_14),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_756),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_667),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_750),
.Y(n_924)
);

INVxp33_ASAP7_75t_L g925 ( 
.A(n_732),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_675),
.B(n_551),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_684),
.B(n_733),
.Y(n_927)
);

CKINVDCx20_ASAP7_75t_R g928 ( 
.A(n_721),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_696),
.B(n_551),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_760),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_754),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_696),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_699),
.A2(n_522),
.B1(n_551),
.B2(n_526),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_SL g934 ( 
.A1(n_673),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_739),
.B(n_16),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_740),
.B(n_744),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_688),
.A2(n_551),
.B1(n_526),
.B2(n_157),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_696),
.B(n_526),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_688),
.A2(n_526),
.B1(n_21),
.B2(n_23),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_753),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_696),
.B(n_155),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_696),
.B(n_85),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_767),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_776),
.B(n_17),
.Y(n_944)
);

NOR3xp33_ASAP7_75t_SL g945 ( 
.A(n_721),
.B(n_768),
.C(n_720),
.Y(n_945)
);

OR2x6_ASAP7_75t_L g946 ( 
.A(n_760),
.B(n_17),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_632),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_627),
.B(n_77),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_650),
.B(n_153),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_766),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_650),
.B(n_76),
.Y(n_951)
);

INVx4_ASAP7_75t_L g952 ( 
.A(n_680),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_668),
.B(n_152),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_647),
.B(n_72),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_726),
.B(n_21),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_727),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_770),
.Y(n_957)
);

AOI22xp5_ASAP7_75t_L g958 ( 
.A1(n_734),
.A2(n_149),
.B1(n_142),
.B2(n_120),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_706),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_734),
.A2(n_88),
.B1(n_61),
.B2(n_59),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_633),
.Y(n_961)
);

NAND2x1p5_ASAP7_75t_L g962 ( 
.A(n_706),
.B(n_58),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_692),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_730),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_785),
.B(n_647),
.Y(n_965)
);

NAND2x1p5_ASAP7_75t_L g966 ( 
.A(n_778),
.B(n_718),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_932),
.A2(n_644),
.B(n_655),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_932),
.A2(n_636),
.B(n_635),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_793),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_835),
.A2(n_666),
.B(n_703),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_782),
.A2(n_741),
.B1(n_735),
.B2(n_713),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_871),
.A2(n_704),
.B(n_709),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_877),
.B(n_735),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_918),
.A2(n_719),
.B1(n_717),
.B2(n_689),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_871),
.A2(n_741),
.B(n_665),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_799),
.B(n_646),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_811),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_878),
.B(n_677),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_842),
.B(n_694),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_839),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_839),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_799),
.B(n_764),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_788),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_791),
.B(n_672),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_L g985 ( 
.A(n_783),
.B(n_764),
.C(n_681),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_940),
.B(n_641),
.Y(n_986)
);

OAI22x1_ASAP7_75t_L g987 ( 
.A1(n_927),
.A2(n_631),
.B1(n_665),
.B2(n_662),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_930),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_L g989 ( 
.A(n_812),
.B(n_697),
.C(n_640),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_818),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_940),
.B(n_639),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_943),
.B(n_649),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_964),
.B(n_654),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_R g994 ( 
.A(n_823),
.B(n_702),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_885),
.B(n_662),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_916),
.B(n_640),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_810),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_843),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_863),
.A2(n_634),
.B(n_631),
.C(n_616),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_915),
.A2(n_634),
.B(n_30),
.C(n_31),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_843),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_800),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_904),
.A2(n_29),
.B(n_30),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_817),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_874),
.B(n_33),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_801),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_803),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_789),
.B(n_36),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_880),
.A2(n_38),
.B(n_42),
.C(n_46),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_904),
.A2(n_51),
.B(n_47),
.Y(n_1010)
);

AOI221xp5_ASAP7_75t_L g1011 ( 
.A1(n_840),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.C(n_49),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_804),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_789),
.B(n_817),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_858),
.Y(n_1014)
);

OR2x6_ASAP7_75t_SL g1015 ( 
.A(n_881),
.B(n_813),
.Y(n_1015)
);

BUFx2_ASAP7_75t_L g1016 ( 
.A(n_808),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_910),
.B(n_917),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_815),
.B(n_833),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_909),
.B(n_880),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_778),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_859),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_854),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_864),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_833),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_929),
.A2(n_938),
.B(n_852),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_928),
.A2(n_956),
.B1(n_922),
.B2(n_902),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_778),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_852),
.B(n_908),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_819),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_814),
.B(n_829),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_830),
.B(n_844),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_955),
.A2(n_816),
.B(n_945),
.C(n_935),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_873),
.Y(n_1033)
);

INVx2_ASAP7_75t_SL g1034 ( 
.A(n_806),
.Y(n_1034)
);

AO32x1_ASAP7_75t_L g1035 ( 
.A1(n_837),
.A2(n_920),
.A3(n_937),
.B1(n_944),
.B2(n_897),
.Y(n_1035)
);

BUFx10_ASAP7_75t_L g1036 ( 
.A(n_827),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_851),
.B(n_891),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_887),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_929),
.A2(n_938),
.B(n_821),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_781),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_866),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_815),
.B(n_906),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_918),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_925),
.B(n_896),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_816),
.A2(n_936),
.B(n_796),
.C(n_825),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_838),
.Y(n_1046)
);

AOI33xp33_ASAP7_75t_L g1047 ( 
.A1(n_934),
.A2(n_959),
.A3(n_939),
.B1(n_855),
.B2(n_886),
.B3(n_914),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_780),
.B(n_850),
.Y(n_1048)
);

A2O1A1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_825),
.A2(n_953),
.B(n_949),
.C(n_951),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_802),
.A2(n_809),
.B1(n_934),
.B2(n_903),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_815),
.B(n_906),
.Y(n_1051)
);

INVxp67_ASAP7_75t_L g1052 ( 
.A(n_860),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_802),
.A2(n_809),
.B1(n_780),
.B2(n_949),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_821),
.A2(n_826),
.B(n_870),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_906),
.B(n_923),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_850),
.B(n_847),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_794),
.Y(n_1057)
);

BUFx8_ASAP7_75t_L g1058 ( 
.A(n_836),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_895),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_786),
.B(n_790),
.Y(n_1060)
);

OAI21x1_ASAP7_75t_L g1061 ( 
.A1(n_879),
.A2(n_882),
.B(n_890),
.Y(n_1061)
);

OA22x2_ASAP7_75t_L g1062 ( 
.A1(n_946),
.A2(n_861),
.B1(n_787),
.B2(n_958),
.Y(n_1062)
);

BUFx6f_ASAP7_75t_L g1063 ( 
.A(n_781),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_884),
.B(n_923),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_889),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_954),
.A2(n_798),
.B1(n_797),
.B2(n_869),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_SL g1067 ( 
.A(n_926),
.B(n_805),
.C(n_931),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_869),
.B(n_822),
.Y(n_1068)
);

OA22x2_ASAP7_75t_L g1069 ( 
.A1(n_946),
.A2(n_960),
.B1(n_822),
.B2(n_883),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_846),
.B(n_953),
.Y(n_1070)
);

BUFx8_ASAP7_75t_L g1071 ( 
.A(n_848),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_846),
.B(n_845),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_826),
.A2(n_868),
.B(n_872),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_857),
.A2(n_868),
.B(n_872),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_856),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_892),
.A2(n_876),
.B1(n_805),
.B2(n_961),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_898),
.B(n_779),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_779),
.A2(n_807),
.B1(n_784),
.B2(n_792),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_912),
.B(n_963),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_857),
.A2(n_865),
.B(n_870),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_924),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_950),
.B(n_957),
.Y(n_1082)
);

NAND2x1p5_ASAP7_75t_L g1083 ( 
.A(n_930),
.B(n_888),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_831),
.B(n_952),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_952),
.B(n_865),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_898),
.A2(n_841),
.B(n_942),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_892),
.A2(n_876),
.B1(n_947),
.B2(n_913),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_879),
.A2(n_890),
.B(n_882),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_779),
.A2(n_807),
.B1(n_792),
.B2(n_784),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_899),
.Y(n_1090)
);

NOR2x1_ASAP7_75t_L g1091 ( 
.A(n_856),
.B(n_807),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_828),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_867),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_SL g1094 ( 
.A1(n_911),
.A2(n_894),
.B(n_824),
.C(n_834),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_948),
.A2(n_946),
.B(n_921),
.C(n_942),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_901),
.A2(n_948),
.B(n_941),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_856),
.Y(n_1097)
);

OR2x6_ASAP7_75t_L g1098 ( 
.A(n_888),
.B(n_905),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_867),
.A2(n_905),
.B1(n_888),
.B2(n_941),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_795),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_905),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_901),
.B(n_862),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_832),
.A2(n_893),
.B(n_849),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_841),
.A2(n_907),
.B(n_919),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_907),
.A2(n_933),
.B(n_893),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_962),
.A2(n_853),
.B1(n_875),
.B2(n_820),
.Y(n_1106)
);

NAND3xp33_ASAP7_75t_SL g1107 ( 
.A(n_962),
.B(n_782),
.C(n_614),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_900),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_900),
.A2(n_782),
.B(n_611),
.C(n_799),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_900),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1096),
.A2(n_900),
.B(n_1028),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1045),
.A2(n_900),
.B(n_1049),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1039),
.A2(n_1054),
.B(n_1061),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1048),
.A2(n_1073),
.B(n_1056),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1020),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1088),
.A2(n_970),
.B(n_972),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_1105),
.A2(n_1025),
.B(n_1102),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1037),
.B(n_1046),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_980),
.B(n_981),
.Y(n_1119)
);

O2A1O1Ixp5_ASAP7_75t_L g1120 ( 
.A1(n_1032),
.A2(n_996),
.B(n_971),
.C(n_974),
.Y(n_1120)
);

O2A1O1Ixp5_ASAP7_75t_L g1121 ( 
.A1(n_971),
.A2(n_1106),
.B(n_1103),
.C(n_1060),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_998),
.B(n_1001),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_967),
.A2(n_968),
.B(n_1080),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1013),
.B(n_1053),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1095),
.A2(n_1074),
.B(n_975),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1104),
.A2(n_1091),
.B(n_999),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1094),
.A2(n_1078),
.B(n_1089),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1053),
.B(n_1050),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_1020),
.Y(n_1129)
);

NAND3xp33_ASAP7_75t_L g1130 ( 
.A(n_1011),
.B(n_1109),
.C(n_995),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1044),
.B(n_1024),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1018),
.B(n_1064),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_987),
.A2(n_1106),
.A3(n_1066),
.B(n_1050),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1022),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_976),
.B(n_982),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1066),
.A2(n_984),
.A3(n_1004),
.B(n_1108),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1019),
.B(n_1015),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_993),
.B(n_986),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_1057),
.B(n_990),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1103),
.A2(n_1076),
.B(n_1086),
.Y(n_1140)
);

OAI22x1_ASAP7_75t_L g1141 ( 
.A1(n_1026),
.A2(n_1043),
.B1(n_1099),
.B2(n_1062),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1107),
.A2(n_1047),
.B(n_989),
.C(n_1067),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1085),
.A2(n_1070),
.B(n_966),
.Y(n_1143)
);

AO32x2_ASAP7_75t_L g1144 ( 
.A1(n_1004),
.A2(n_1035),
.A3(n_1097),
.B1(n_1069),
.B2(n_1062),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_991),
.B(n_992),
.Y(n_1145)
);

INVxp67_ASAP7_75t_L g1146 ( 
.A(n_1021),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_983),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1069),
.A2(n_965),
.B(n_1077),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1092),
.A2(n_1100),
.B(n_1084),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1008),
.A2(n_977),
.B1(n_1023),
.B2(n_1041),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1030),
.B(n_1031),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_978),
.B(n_1005),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1097),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_966),
.A2(n_1072),
.B(n_1079),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_979),
.A2(n_985),
.B(n_1110),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1082),
.A2(n_1083),
.B(n_1087),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1017),
.A2(n_1068),
.B(n_979),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1033),
.B(n_1065),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_997),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1081),
.A2(n_1090),
.B1(n_1059),
.B2(n_1038),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1002),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1093),
.B(n_1014),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1035),
.A2(n_1010),
.A3(n_1003),
.B(n_1007),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_983),
.Y(n_1164)
);

NOR4xp25_ASAP7_75t_L g1165 ( 
.A(n_1009),
.B(n_1000),
.C(n_1012),
.D(n_1006),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1055),
.B(n_988),
.Y(n_1166)
);

BUFx2_ASAP7_75t_SL g1167 ( 
.A(n_1016),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1098),
.A2(n_1051),
.B(n_1042),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1098),
.A2(n_1083),
.B(n_1101),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1034),
.B(n_1101),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1098),
.A2(n_1101),
.B(n_1075),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1020),
.A2(n_1040),
.B(n_1027),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1052),
.B(n_1040),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1027),
.B(n_1040),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_994),
.B(n_1027),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1063),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1063),
.A2(n_1036),
.B(n_1029),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1063),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1036),
.B(n_1058),
.Y(n_1179)
);

OAI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1058),
.A2(n_782),
.B1(n_612),
.B2(n_916),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1071),
.A2(n_1039),
.B(n_1054),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_1071),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_R g1183 ( 
.A(n_994),
.B(n_467),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_SL g1184 ( 
.A(n_1017),
.B(n_842),
.Y(n_1184)
);

O2A1O1Ixp5_ASAP7_75t_L g1185 ( 
.A1(n_1032),
.A2(n_791),
.B(n_645),
.C(n_611),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1024),
.B(n_1046),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_980),
.B(n_981),
.Y(n_1187)
);

AOI221x1_ASAP7_75t_L g1188 ( 
.A1(n_1032),
.A2(n_1107),
.B1(n_1004),
.B2(n_971),
.C(n_1045),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_1058),
.Y(n_1189)
);

NAND2x1_ASAP7_75t_L g1190 ( 
.A(n_1098),
.B(n_678),
.Y(n_1190)
);

NAND2x1p5_ASAP7_75t_L g1191 ( 
.A(n_1091),
.B(n_1097),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_976),
.B(n_314),
.Y(n_1192)
);

INVxp67_ASAP7_75t_SL g1193 ( 
.A(n_1068),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1096),
.A2(n_932),
.B(n_652),
.Y(n_1194)
);

O2A1O1Ixp5_ASAP7_75t_SL g1195 ( 
.A1(n_1004),
.A2(n_915),
.B(n_996),
.C(n_863),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_995),
.B(n_783),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1096),
.A2(n_932),
.B(n_652),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1050),
.A2(n_782),
.B1(n_612),
.B2(n_916),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1024),
.B(n_1046),
.Y(n_1199)
);

OAI22x1_ASAP7_75t_L g1200 ( 
.A1(n_1044),
.A2(n_464),
.B1(n_663),
.B2(n_1060),
.Y(n_1200)
);

OAI22xp5_ASAP7_75t_L g1201 ( 
.A1(n_1050),
.A2(n_782),
.B1(n_612),
.B2(n_916),
.Y(n_1201)
);

O2A1O1Ixp5_ASAP7_75t_L g1202 ( 
.A1(n_1032),
.A2(n_791),
.B(n_645),
.C(n_611),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1020),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_980),
.B(n_981),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_976),
.B(n_314),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_987),
.A2(n_1045),
.A3(n_1054),
.B(n_1096),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_969),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1049),
.A2(n_932),
.B(n_1053),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_983),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1096),
.A2(n_1073),
.B(n_1039),
.Y(n_1210)
);

NOR2x1_ASAP7_75t_SL g1211 ( 
.A(n_1098),
.B(n_779),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1058),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1097),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1109),
.A2(n_782),
.B(n_916),
.C(n_611),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1045),
.A2(n_1049),
.B(n_782),
.Y(n_1215)
);

NAND2xp33_ASAP7_75t_L g1216 ( 
.A(n_973),
.B(n_782),
.Y(n_1216)
);

AOI221xp5_ASAP7_75t_L g1217 ( 
.A1(n_1011),
.A2(n_540),
.B1(n_537),
.B2(n_663),
.C(n_782),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1045),
.A2(n_1049),
.B(n_782),
.Y(n_1218)
);

AOI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1105),
.A2(n_975),
.B(n_1039),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1096),
.A2(n_932),
.B(n_652),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_969),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1020),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_976),
.B(n_314),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1096),
.A2(n_932),
.B(n_652),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_969),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_990),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_SL g1227 ( 
.A(n_1011),
.B(n_782),
.C(n_614),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_995),
.B(n_783),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_976),
.B(n_314),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1096),
.A2(n_932),
.B(n_652),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_SL g1231 ( 
.A(n_1029),
.B(n_765),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1032),
.A2(n_927),
.B(n_1049),
.C(n_1045),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_969),
.Y(n_1233)
);

INVx2_ASAP7_75t_SL g1234 ( 
.A(n_983),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1037),
.B(n_785),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1037),
.B(n_785),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1037),
.B(n_785),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1020),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_987),
.A2(n_1045),
.A3(n_1054),
.B(n_1096),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_969),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1045),
.A2(n_1049),
.B(n_782),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1037),
.B(n_785),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1037),
.B(n_785),
.Y(n_1243)
);

OAI21xp33_ASAP7_75t_L g1244 ( 
.A1(n_995),
.A2(n_782),
.B(n_614),
.Y(n_1244)
);

BUFx8_ASAP7_75t_L g1245 ( 
.A(n_1189),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_1159),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1211),
.B(n_1132),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1139),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1135),
.B(n_1242),
.Y(n_1249)
);

OR2x6_ASAP7_75t_L g1250 ( 
.A(n_1208),
.B(n_1112),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1151),
.Y(n_1251)
);

INVx3_ASAP7_75t_SL g1252 ( 
.A(n_1226),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1217),
.A2(n_1227),
.B1(n_1244),
.B2(n_1130),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1129),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1181),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1114),
.A2(n_1197),
.B(n_1194),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1123),
.A2(n_1126),
.B(n_1113),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1130),
.A2(n_1244),
.B1(n_1228),
.B2(n_1196),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1125),
.A2(n_1188),
.B(n_1121),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1185),
.A2(n_1202),
.B(n_1214),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1119),
.B(n_1122),
.Y(n_1261)
);

A2O1A1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1215),
.A2(n_1218),
.B(n_1241),
.C(n_1201),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1116),
.A2(n_1219),
.B(n_1230),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_1112),
.B(n_1215),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1153),
.B(n_1213),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1198),
.A2(n_1201),
.B(n_1241),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1132),
.B(n_1153),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1198),
.A2(n_1180),
.B1(n_1232),
.B2(n_1200),
.C(n_1216),
.Y(n_1268)
);

OA21x2_ASAP7_75t_L g1269 ( 
.A1(n_1127),
.A2(n_1140),
.B(n_1128),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1220),
.A2(n_1224),
.B(n_1111),
.Y(n_1270)
);

CKINVDCx20_ASAP7_75t_R g1271 ( 
.A(n_1212),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1128),
.B(n_1124),
.Y(n_1272)
);

AND2x6_ASAP7_75t_SL g1273 ( 
.A(n_1179),
.B(n_1192),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1138),
.B(n_1145),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1142),
.A2(n_1180),
.B(n_1152),
.C(n_1124),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1184),
.B(n_1148),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1120),
.A2(n_1149),
.B(n_1155),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1207),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1143),
.A2(n_1154),
.B(n_1210),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1210),
.A2(n_1156),
.B(n_1117),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1118),
.B(n_1235),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1117),
.A2(n_1195),
.B(n_1155),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1221),
.Y(n_1283)
);

OA21x2_ASAP7_75t_L g1284 ( 
.A1(n_1157),
.A2(n_1187),
.B(n_1119),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1184),
.A2(n_1229),
.B1(n_1223),
.B2(n_1205),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1137),
.A2(n_1141),
.B1(n_1199),
.B2(n_1186),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1186),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1122),
.B(n_1187),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1204),
.A2(n_1150),
.B(n_1160),
.Y(n_1289)
);

AOI222xp33_ASAP7_75t_L g1290 ( 
.A1(n_1236),
.A2(n_1243),
.B1(n_1237),
.B2(n_1131),
.C1(n_1150),
.C2(n_1199),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1168),
.A2(n_1191),
.B(n_1169),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1182),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1193),
.A2(n_1190),
.B(n_1165),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1146),
.A2(n_1231),
.B1(n_1167),
.B2(n_1161),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1165),
.A2(n_1206),
.B(n_1239),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1225),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1173),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1129),
.Y(n_1298)
);

AOI221xp5_ASAP7_75t_L g1299 ( 
.A1(n_1233),
.A2(n_1240),
.B1(n_1158),
.B2(n_1177),
.C(n_1162),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1166),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1176),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1147),
.A2(n_1234),
.B1(n_1209),
.B2(n_1164),
.Y(n_1302)
);

XNOR2xp5_ASAP7_75t_L g1303 ( 
.A(n_1175),
.B(n_1171),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1191),
.A2(n_1172),
.B(n_1178),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1206),
.A2(n_1239),
.B(n_1133),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1170),
.A2(n_1174),
.B1(n_1183),
.B2(n_1115),
.Y(n_1307)
);

AO21x2_ASAP7_75t_L g1308 ( 
.A1(n_1206),
.A2(n_1239),
.B(n_1133),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1133),
.A2(n_1163),
.B(n_1136),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1163),
.A2(n_1136),
.B(n_1144),
.Y(n_1310)
);

AOI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1174),
.A2(n_1115),
.B1(n_1203),
.B2(n_1222),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1115),
.B(n_1203),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_R g1313 ( 
.A(n_1203),
.B(n_1222),
.Y(n_1313)
);

AOI21xp33_ASAP7_75t_L g1314 ( 
.A1(n_1238),
.A2(n_1144),
.B(n_1163),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1238),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1316)
);

BUFx2_ASAP7_75t_R g1317 ( 
.A(n_1147),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1211),
.B(n_1097),
.Y(n_1318)
);

INVx4_ASAP7_75t_SL g1319 ( 
.A(n_1136),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1139),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1135),
.B(n_915),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1135),
.B(n_915),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1137),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1324)
);

NAND2x1p5_ASAP7_75t_L g1325 ( 
.A(n_1153),
.B(n_1091),
.Y(n_1325)
);

AND2x4_ASAP7_75t_L g1326 ( 
.A(n_1211),
.B(n_1097),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1149),
.A2(n_1111),
.B(n_987),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1134),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1211),
.B(n_1097),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1134),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1129),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1134),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1226),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1125),
.A2(n_1188),
.B(n_1121),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1135),
.B(n_915),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1134),
.Y(n_1339)
);

AO21x2_ASAP7_75t_L g1340 ( 
.A1(n_1125),
.A2(n_1218),
.B(n_1215),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1135),
.B(n_915),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1217),
.A2(n_1227),
.B1(n_1244),
.B2(n_842),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1159),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1125),
.A2(n_1188),
.B(n_1121),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1129),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1125),
.A2(n_1188),
.B(n_1121),
.Y(n_1348)
);

NOR3xp33_ASAP7_75t_L g1349 ( 
.A(n_1217),
.B(n_791),
.C(n_459),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1193),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1217),
.A2(n_1227),
.B1(n_1244),
.B2(n_842),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1129),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_SL g1353 ( 
.A1(n_1214),
.A2(n_1201),
.B(n_1198),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1126),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1134),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1125),
.A2(n_1218),
.B(n_1215),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1318),
.A2(n_1331),
.B(n_1326),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1253),
.A2(n_1351),
.B1(n_1343),
.B2(n_1285),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1336),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1256),
.A2(n_1250),
.B(n_1262),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1350),
.A2(n_1262),
.B(n_1250),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1251),
.B(n_1281),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1287),
.Y(n_1363)
);

O2A1O1Ixp33_ASAP7_75t_L g1364 ( 
.A1(n_1349),
.A2(n_1275),
.B(n_1266),
.C(n_1258),
.Y(n_1364)
);

A2O1A1Ixp33_ASAP7_75t_L g1365 ( 
.A1(n_1268),
.A2(n_1260),
.B(n_1276),
.C(n_1293),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1294),
.A2(n_1286),
.B1(n_1250),
.B2(n_1323),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1250),
.A2(n_1264),
.B(n_1356),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1280),
.A2(n_1282),
.B(n_1279),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1274),
.B(n_1261),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1261),
.B(n_1288),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1247),
.B(n_1267),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1288),
.B(n_1249),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1321),
.B(n_1322),
.Y(n_1374)
);

AND2x2_ASAP7_75t_SL g1375 ( 
.A(n_1259),
.B(n_1337),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1248),
.B(n_1320),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1338),
.B(n_1341),
.Y(n_1377)
);

INVx1_ASAP7_75t_SL g1378 ( 
.A(n_1297),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_SL g1379 ( 
.A1(n_1247),
.A2(n_1338),
.B(n_1341),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1264),
.A2(n_1303),
.B1(n_1272),
.B2(n_1302),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1290),
.B(n_1267),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1336),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1267),
.B(n_1300),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1264),
.A2(n_1272),
.B1(n_1353),
.B2(n_1276),
.Y(n_1384)
);

NOR2xp67_ASAP7_75t_L g1385 ( 
.A(n_1248),
.B(n_1320),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1246),
.B(n_1345),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1299),
.A2(n_1305),
.B(n_1291),
.C(n_1275),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1291),
.A2(n_1278),
.B(n_1283),
.C(n_1296),
.Y(n_1388)
);

OR2x6_ASAP7_75t_L g1389 ( 
.A(n_1255),
.B(n_1289),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1315),
.B(n_1301),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1307),
.A2(n_1317),
.B1(n_1311),
.B2(n_1252),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1252),
.A2(n_1325),
.B1(n_1355),
.B2(n_1330),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1315),
.B(n_1332),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1335),
.B(n_1339),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1340),
.A2(n_1337),
.B(n_1346),
.C(n_1259),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1265),
.A2(n_1289),
.B1(n_1254),
.B2(n_1347),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1284),
.B(n_1273),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1284),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1295),
.B(n_1308),
.Y(n_1399)
);

O2A1O1Ixp5_ASAP7_75t_L g1400 ( 
.A1(n_1328),
.A2(n_1314),
.B(n_1255),
.C(n_1298),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1277),
.B(n_1348),
.Y(n_1401)
);

OA21x2_ASAP7_75t_L g1402 ( 
.A1(n_1263),
.A2(n_1354),
.B(n_1334),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1292),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1312),
.B(n_1295),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1333),
.B(n_1352),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1308),
.B(n_1313),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1309),
.A2(n_1310),
.B(n_1270),
.C(n_1304),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1292),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1308),
.B(n_1269),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1306),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_SL g1411 ( 
.A1(n_1319),
.A2(n_1309),
.B(n_1310),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1304),
.B(n_1319),
.Y(n_1412)
);

INVx1_ASAP7_75t_SL g1413 ( 
.A(n_1271),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1245),
.Y(n_1414)
);

AND2x6_ASAP7_75t_L g1415 ( 
.A(n_1245),
.B(n_1257),
.Y(n_1415)
);

O2A1O1Ixp5_ASAP7_75t_L g1416 ( 
.A1(n_1316),
.A2(n_1327),
.B(n_1344),
.C(n_1342),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1245),
.A2(n_1329),
.B(n_1344),
.C(n_1342),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1257),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1324),
.B(n_1329),
.Y(n_1419)
);

NOR2xp67_ASAP7_75t_L g1420 ( 
.A(n_1248),
.B(n_1320),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1274),
.B(n_1135),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1349),
.A2(n_1217),
.B(n_1227),
.C(n_1244),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1253),
.A2(n_1217),
.B1(n_782),
.B2(n_842),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1398),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1365),
.B(n_1375),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1423),
.B(n_1358),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1389),
.B(n_1418),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1388),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1389),
.B(n_1412),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1375),
.B(n_1409),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1368),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1401),
.B(n_1367),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1401),
.B(n_1404),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1388),
.Y(n_1434)
);

BUFx2_ASAP7_75t_L g1435 ( 
.A(n_1389),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1399),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1365),
.B(n_1360),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1384),
.B(n_1370),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1413),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1396),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1395),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1397),
.B(n_1407),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1406),
.B(n_1419),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1416),
.A2(n_1387),
.B(n_1400),
.Y(n_1444)
);

OAI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1364),
.A2(n_1422),
.B(n_1387),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1374),
.B(n_1377),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_1380),
.B(n_1392),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1415),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1371),
.B(n_1415),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1417),
.A2(n_1361),
.B(n_1411),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1402),
.B(n_1373),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1381),
.B(n_1366),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1369),
.B(n_1421),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1426),
.A2(n_1362),
.B1(n_1378),
.B2(n_1391),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1433),
.B(n_1383),
.Y(n_1455)
);

AOI33xp33_ASAP7_75t_L g1456 ( 
.A1(n_1441),
.A2(n_1394),
.A3(n_1393),
.B1(n_1390),
.B2(n_1371),
.B3(n_1405),
.Y(n_1456)
);

NAND2xp5_ASAP7_75t_L g1457 ( 
.A(n_1451),
.B(n_1372),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1433),
.B(n_1390),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1442),
.B(n_1386),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1431),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1426),
.A2(n_1363),
.B1(n_1394),
.B2(n_1414),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1442),
.B(n_1393),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1424),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1424),
.Y(n_1464)
);

INVx3_ASAP7_75t_L g1465 ( 
.A(n_1427),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1451),
.B(n_1415),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1451),
.B(n_1415),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1443),
.B(n_1414),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1442),
.B(n_1408),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1431),
.Y(n_1470)
);

BUFx6f_ASAP7_75t_SL g1471 ( 
.A(n_1448),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1430),
.B(n_1379),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1442),
.B(n_1382),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1427),
.Y(n_1474)
);

INVx5_ASAP7_75t_SL g1475 ( 
.A(n_1450),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1451),
.B(n_1359),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1430),
.B(n_1379),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1427),
.B(n_1357),
.Y(n_1478)
);

INVx1_ASAP7_75t_SL g1479 ( 
.A(n_1432),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1430),
.B(n_1357),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1469),
.Y(n_1481)
);

AOI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1469),
.A2(n_1437),
.B(n_1445),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1463),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1480),
.B(n_1430),
.Y(n_1484)
);

BUFx2_ASAP7_75t_SL g1485 ( 
.A(n_1471),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1459),
.B(n_1438),
.Y(n_1486)
);

NOR2x1_ASAP7_75t_L g1487 ( 
.A(n_1469),
.B(n_1437),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1463),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1463),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1454),
.A2(n_1437),
.B(n_1445),
.Y(n_1490)
);

NAND3xp33_ASAP7_75t_L g1491 ( 
.A(n_1454),
.B(n_1445),
.C(n_1440),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1461),
.A2(n_1447),
.B1(n_1425),
.B2(n_1452),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1478),
.B(n_1474),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1479),
.B(n_1441),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1464),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1473),
.A2(n_1447),
.B1(n_1452),
.B2(n_1438),
.Y(n_1496)
);

NAND3xp33_ASAP7_75t_L g1497 ( 
.A(n_1473),
.B(n_1440),
.C(n_1438),
.Y(n_1497)
);

AOI211xp5_ASAP7_75t_L g1498 ( 
.A1(n_1473),
.A2(n_1425),
.B(n_1441),
.C(n_1432),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1480),
.B(n_1432),
.Y(n_1499)
);

BUFx6f_ASAP7_75t_L g1500 ( 
.A(n_1478),
.Y(n_1500)
);

AND4x1_ASAP7_75t_L g1501 ( 
.A(n_1456),
.B(n_1425),
.C(n_1428),
.D(n_1434),
.Y(n_1501)
);

AOI221xp5_ASAP7_75t_L g1502 ( 
.A1(n_1476),
.A2(n_1453),
.B1(n_1434),
.B2(n_1428),
.C(n_1446),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1479),
.B(n_1436),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1476),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1472),
.B(n_1429),
.Y(n_1505)
);

OAI31xp33_ASAP7_75t_L g1506 ( 
.A1(n_1472),
.A2(n_1434),
.A3(n_1428),
.B(n_1435),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1461),
.A2(n_1453),
.B1(n_1448),
.B2(n_1449),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1474),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_L g1509 ( 
.A(n_1459),
.B(n_1439),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1472),
.A2(n_1429),
.B1(n_1439),
.B2(n_1450),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1483),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1490),
.A2(n_1450),
.B(n_1444),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1483),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1488),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1499),
.B(n_1465),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1494),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1488),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1465),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1489),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1489),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1495),
.Y(n_1522)
);

INVx8_ASAP7_75t_L g1523 ( 
.A(n_1500),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1500),
.Y(n_1524)
);

AOI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1487),
.A2(n_1470),
.B(n_1460),
.Y(n_1525)
);

NOR3xp33_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1456),
.C(n_1376),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1500),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1498),
.B(n_1478),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1494),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1484),
.B(n_1465),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1487),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1511),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1511),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1513),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1513),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1524),
.B(n_1493),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1516),
.B(n_1459),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1516),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1526),
.B(n_1482),
.Y(n_1541)
);

NOR3xp33_ASAP7_75t_L g1542 ( 
.A(n_1526),
.B(n_1492),
.C(n_1497),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1529),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1525),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1518),
.B(n_1509),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1518),
.B(n_1403),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1514),
.Y(n_1547)
);

AOI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1512),
.A2(n_1496),
.B1(n_1498),
.B2(n_1502),
.C(n_1504),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1531),
.B(n_1481),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1531),
.B(n_1481),
.Y(n_1550)
);

NOR2x1_ASAP7_75t_L g1551 ( 
.A(n_1528),
.B(n_1485),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1527),
.B(n_1505),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1527),
.B(n_1505),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1514),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1528),
.B(n_1484),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1517),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1517),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1520),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1512),
.B(n_1455),
.Y(n_1560)
);

AND3x2_ASAP7_75t_L g1561 ( 
.A(n_1530),
.B(n_1506),
.C(n_1508),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1530),
.B(n_1500),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1520),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1530),
.B(n_1500),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1523),
.B(n_1410),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1525),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1521),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

NAND4xp25_ASAP7_75t_SL g1570 ( 
.A(n_1515),
.B(n_1510),
.C(n_1477),
.D(n_1467),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1523),
.B(n_1468),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1515),
.B(n_1508),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.B(n_1462),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1543),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1542),
.A2(n_1548),
.B1(n_1570),
.B2(n_1551),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1551),
.B(n_1515),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1533),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1533),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1534),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1545),
.B(n_1468),
.Y(n_1581)
);

INVxp33_ASAP7_75t_L g1582 ( 
.A(n_1565),
.Y(n_1582)
);

OAI32xp33_ASAP7_75t_L g1583 ( 
.A1(n_1549),
.A2(n_1466),
.A3(n_1467),
.B1(n_1503),
.B2(n_1462),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1550),
.B(n_1560),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1544),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1546),
.B(n_1468),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1556),
.B(n_1519),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1540),
.B(n_1457),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1539),
.B(n_1455),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1556),
.B(n_1519),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1535),
.Y(n_1591)
);

INVxp67_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1539),
.B(n_1503),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1544),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1536),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1536),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1553),
.B(n_1446),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1547),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1553),
.B(n_1554),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1571),
.B(n_1507),
.C(n_1477),
.D(n_1385),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1547),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1532),
.B(n_1537),
.Y(n_1602)
);

NOR2x1_ASAP7_75t_L g1603 ( 
.A(n_1544),
.B(n_1566),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1532),
.B(n_1519),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1554),
.B(n_1458),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1561),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1602),
.B(n_1537),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1591),
.Y(n_1608)
);

INVx2_ASAP7_75t_SL g1609 ( 
.A(n_1602),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1606),
.B(n_1538),
.Y(n_1610)
);

NAND3xp33_ASAP7_75t_L g1611 ( 
.A(n_1575),
.B(n_1501),
.C(n_1566),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1606),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1582),
.Y(n_1613)
);

NAND2x1p5_ASAP7_75t_L g1614 ( 
.A(n_1606),
.B(n_1501),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1590),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1591),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_L g1617 ( 
.A1(n_1600),
.A2(n_1582),
.B1(n_1573),
.B2(n_1584),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1574),
.A2(n_1475),
.B1(n_1538),
.B2(n_1552),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1576),
.B(n_1552),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1577),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1578),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1562),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1599),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1579),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1562),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1592),
.A2(n_1475),
.B1(n_1450),
.B2(n_1477),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1588),
.B(n_1555),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_R g1630 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1592),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1611),
.A2(n_1581),
.B1(n_1604),
.B2(n_1598),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1623),
.B(n_1604),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1613),
.B(n_1597),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1631),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1631),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1612),
.Y(n_1637)
);

INVxp67_ASAP7_75t_SL g1638 ( 
.A(n_1612),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1608),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1608),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1616),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1610),
.B(n_1572),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1616),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1572),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1624),
.B(n_1580),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1609),
.B(n_1595),
.Y(n_1646)
);

NAND2x1_ASAP7_75t_L g1647 ( 
.A(n_1610),
.B(n_1603),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1614),
.A2(n_1586),
.B1(n_1605),
.B2(n_1589),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1621),
.Y(n_1649)
);

NAND4xp25_ASAP7_75t_SL g1650 ( 
.A(n_1611),
.B(n_1593),
.C(n_1596),
.D(n_1601),
.Y(n_1650)
);

AOI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1614),
.B1(n_1609),
.B2(n_1632),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1634),
.B(n_1615),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1642),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1633),
.A2(n_1614),
.B1(n_1610),
.B2(n_1626),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1645),
.B(n_1615),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1638),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1642),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1644),
.B(n_1623),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1644),
.B(n_1619),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1636),
.B(n_1619),
.Y(n_1661)
);

NOR3xp33_ASAP7_75t_L g1662 ( 
.A(n_1659),
.B(n_1637),
.C(n_1638),
.Y(n_1662)
);

OAI31xp33_ASAP7_75t_L g1663 ( 
.A1(n_1656),
.A2(n_1648),
.A3(n_1637),
.B(n_1640),
.Y(n_1663)
);

AOI321xp33_ASAP7_75t_L g1664 ( 
.A1(n_1651),
.A2(n_1643),
.A3(n_1641),
.B1(n_1639),
.B2(n_1646),
.C(n_1649),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1656),
.Y(n_1665)
);

OAI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1654),
.A2(n_1647),
.B(n_1628),
.Y(n_1666)
);

AOI222xp33_ASAP7_75t_L g1667 ( 
.A1(n_1661),
.A2(n_1625),
.B1(n_1621),
.B2(n_1622),
.C1(n_1630),
.C2(n_1626),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1627),
.Y(n_1668)
);

OAI31xp33_ASAP7_75t_L g1669 ( 
.A1(n_1657),
.A2(n_1626),
.A3(n_1630),
.B(n_1620),
.Y(n_1669)
);

OAI32xp33_ASAP7_75t_L g1670 ( 
.A1(n_1655),
.A2(n_1653),
.A3(n_1652),
.B1(n_1660),
.B2(n_1622),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1659),
.A2(n_1626),
.B1(n_1620),
.B2(n_1607),
.Y(n_1671)
);

AOI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1665),
.A2(n_1625),
.B(n_1594),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1668),
.Y(n_1673)
);

A2O1A1Ixp33_ASAP7_75t_SL g1674 ( 
.A1(n_1662),
.A2(n_1585),
.B(n_1594),
.C(n_1618),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1671),
.B(n_1607),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_SL g1676 ( 
.A1(n_1666),
.A2(n_1627),
.B1(n_1583),
.B2(n_1523),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_SL g1677 ( 
.A(n_1676),
.B(n_1663),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1672),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1675),
.A2(n_1667),
.B(n_1669),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1673),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1674),
.B(n_1670),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1629),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1678),
.B(n_1585),
.Y(n_1683)
);

INVxp67_ASAP7_75t_SL g1684 ( 
.A(n_1682),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1680),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1679),
.B(n_1629),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1681),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1685),
.B(n_1677),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1686),
.B(n_1687),
.Y(n_1689)
);

NAND3xp33_ASAP7_75t_L g1690 ( 
.A(n_1686),
.B(n_1664),
.C(n_1628),
.Y(n_1690)
);

NOR3x2_ASAP7_75t_L g1691 ( 
.A(n_1689),
.B(n_1684),
.C(n_1683),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1691),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1692),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1692),
.Y(n_1694)
);

INVxp67_ASAP7_75t_SL g1695 ( 
.A(n_1693),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1694),
.B(n_1688),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1696),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1695),
.A2(n_1690),
.B1(n_1566),
.B2(n_1569),
.Y(n_1698)
);

OAI22xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1697),
.A2(n_1420),
.B1(n_1569),
.B2(n_1568),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1698),
.B(n_1563),
.Y(n_1700)
);

NAND2x1p5_ASAP7_75t_L g1701 ( 
.A(n_1700),
.B(n_1555),
.Y(n_1701)
);

AO21x2_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1557),
.B(n_1568),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1558),
.B1(n_1567),
.B2(n_1563),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1567),
.B(n_1559),
.C(n_1558),
.Y(n_1704)
);


endmodule