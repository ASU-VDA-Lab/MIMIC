module fake_aes_9216_n_716 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_716);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_235;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_75), .Y(n_80) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_60), .Y(n_81) );
INVxp33_ASAP7_75t_SL g82 ( .A(n_55), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_52), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_54), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_4), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_14), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_1), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_7), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_19), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_13), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_6), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_24), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_7), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_18), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_27), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_5), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_37), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_6), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_3), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_2), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_48), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_26), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_15), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_39), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_61), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_18), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_64), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVxp67_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_19), .Y(n_111) );
BUFx3_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_35), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_22), .Y(n_114) );
BUFx3_ASAP7_75t_L g115 ( .A(n_65), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_56), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_34), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_70), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_11), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_67), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_78), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_30), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_23), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_32), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_45), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_62), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_44), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_122), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_116), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_121), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g132 ( .A(n_113), .B(n_0), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_100), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_80), .B(n_0), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_95), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_90), .B(n_1), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_123), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_95), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_84), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_106), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_107), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_113), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_110), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_85), .B(n_2), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_106), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_114), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_119), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_114), .Y(n_157) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_92), .A2(n_38), .B(n_77), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_86), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_126), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_86), .B(n_87), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_89), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_113), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_126), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_89), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_91), .B(n_4), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_81), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_91), .Y(n_170) );
INVxp67_ASAP7_75t_L g171 ( .A(n_101), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_93), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_135), .B(n_93), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_151), .B(n_99), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_151), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_138), .B(n_109), .Y(n_178) );
OR2x2_ASAP7_75t_L g179 ( .A(n_150), .B(n_94), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_161), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_171), .B(n_94), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_161), .B(n_144), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_133), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_161), .B(n_96), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_156), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_138), .B(n_102), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_133), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_167), .A2(n_104), .B1(n_96), .B2(n_99), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_133), .Y(n_191) );
NAND3xp33_ASAP7_75t_L g192 ( .A(n_139), .B(n_98), .C(n_127), .Y(n_192) );
INVx5_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_162), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_167), .A2(n_129), .B1(n_152), .B2(n_165), .Y(n_195) );
INVx8_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_144), .B(n_98), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_149), .B(n_120), .Y(n_199) );
NAND3xp33_ASAP7_75t_L g200 ( .A(n_160), .B(n_127), .C(n_97), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_169), .B(n_82), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_163), .B(n_111), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_165), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_147), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_172), .Y(n_210) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_129), .Y(n_213) );
AND2x6_ASAP7_75t_L g214 ( .A(n_149), .B(n_97), .Y(n_214) );
INVx5_ASAP7_75t_L g215 ( .A(n_147), .Y(n_215) );
INVx5_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_154), .B(n_103), .Y(n_218) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_136), .B(n_117), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_153), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_140), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_143), .Y(n_223) );
AND2x4_ASAP7_75t_L g224 ( .A(n_134), .B(n_117), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_143), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_137), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_148), .B(n_120), .Y(n_227) );
NAND2x1p5_ASAP7_75t_L g228 ( .A(n_132), .B(n_105), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_164), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_155), .A2(n_124), .B1(n_115), .B2(n_112), .Y(n_230) );
AND2x4_ASAP7_75t_L g231 ( .A(n_158), .B(n_115), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_158), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_157), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_164), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_164), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_169), .A2(n_128), .B1(n_125), .B2(n_118), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_166), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_180), .Y(n_238) );
INVx4_ASAP7_75t_L g239 ( .A(n_196), .Y(n_239) );
BUFx8_ASAP7_75t_L g240 ( .A(n_233), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_180), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_231), .B(n_112), .Y(n_242) );
OR2x4_ASAP7_75t_L g243 ( .A(n_202), .B(n_146), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_231), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
NOR3xp33_ASAP7_75t_SL g246 ( .A(n_195), .B(n_130), .C(n_131), .Y(n_246) );
BUFx4f_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
INVx3_ASAP7_75t_SL g248 ( .A(n_196), .Y(n_248) );
INVx5_ASAP7_75t_L g249 ( .A(n_214), .Y(n_249) );
INVx1_ASAP7_75t_SL g250 ( .A(n_196), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_222), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_231), .B(n_108), .Y(n_252) );
INVx2_ASAP7_75t_SL g253 ( .A(n_175), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_175), .Y(n_254) );
NOR2xp33_ASAP7_75t_R g255 ( .A(n_213), .B(n_141), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_187), .B(n_166), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_179), .B(n_146), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_232), .A2(n_166), .B(n_40), .Y(n_258) );
AOI21x1_ASAP7_75t_L g259 ( .A1(n_198), .A2(n_166), .B(n_41), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_205), .Y(n_261) );
INVx4_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_184), .Y(n_263) );
OAI22xp5_ASAP7_75t_SL g264 ( .A1(n_213), .A2(n_5), .B1(n_8), .B2(n_9), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_187), .Y(n_266) );
XOR2xp5_ASAP7_75t_L g267 ( .A(n_205), .B(n_8), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_178), .B(n_166), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_185), .B(n_42), .Y(n_270) );
BUFx8_ASAP7_75t_L g271 ( .A(n_173), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_190), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_182), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_232), .B(n_43), .Y(n_276) );
INVx6_ASAP7_75t_L g277 ( .A(n_224), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_226), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_186), .B(n_47), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_214), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_173), .B(n_10), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_211), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_179), .B(n_12), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_194), .B(n_49), .Y(n_285) );
INVx5_ASAP7_75t_L g286 ( .A(n_214), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_209), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_219), .A2(n_12), .B1(n_13), .B2(n_14), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_181), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_220), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_176), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
AND2x4_ASAP7_75t_L g293 ( .A(n_181), .B(n_16), .Y(n_293) );
INVx6_ASAP7_75t_L g294 ( .A(n_224), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_177), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_207), .B(n_53), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_224), .Y(n_297) );
INVx4_ASAP7_75t_L g298 ( .A(n_214), .Y(n_298) );
BUFx3_ASAP7_75t_L g299 ( .A(n_204), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_204), .B(n_17), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_210), .Y(n_301) );
INVx4_ASAP7_75t_L g302 ( .A(n_214), .Y(n_302) );
AND2x4_ASAP7_75t_L g303 ( .A(n_197), .B(n_20), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_228), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_228), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_188), .B(n_21), .Y(n_306) );
BUFx6f_ASAP7_75t_L g307 ( .A(n_214), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_239), .B(n_212), .Y(n_310) );
AOI21x1_ASAP7_75t_L g311 ( .A1(n_242), .A2(n_198), .B(n_199), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_266), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_260), .Y(n_313) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_239), .B(n_227), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_242), .A2(n_218), .B(n_199), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_260), .Y(n_317) );
BUFx6f_ASAP7_75t_L g318 ( .A(n_244), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_244), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_271), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_244), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_277), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_253), .B(n_200), .Y(n_323) );
OAI21x1_ASAP7_75t_L g324 ( .A1(n_258), .A2(n_227), .B(n_230), .Y(n_324) );
INVx6_ASAP7_75t_L g325 ( .A(n_262), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_245), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_298), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_298), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_301), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_254), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_252), .A2(n_192), .B(n_219), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_307), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_297), .B(n_236), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
CKINVDCx8_ASAP7_75t_R g336 ( .A(n_283), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_265), .Y(n_338) );
NOR2x1_ASAP7_75t_L g339 ( .A(n_284), .B(n_234), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_307), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_247), .B(n_216), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
NAND2x1p5_ASAP7_75t_L g343 ( .A(n_247), .B(n_216), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_248), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_262), .B(n_25), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_289), .A2(n_237), .B(n_189), .Y(n_346) );
INVx4_ASAP7_75t_L g347 ( .A(n_248), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_277), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_277), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_294), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_249), .Y(n_351) );
INVx5_ASAP7_75t_L g352 ( .A(n_249), .Y(n_352) );
AOI222xp33_ASAP7_75t_L g353 ( .A1(n_299), .A2(n_193), .B1(n_215), .B2(n_216), .C1(n_217), .C2(n_201), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_281), .B(n_28), .Y(n_354) );
CKINVDCx11_ASAP7_75t_R g355 ( .A(n_261), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_294), .A2(n_206), .B1(n_189), .B2(n_201), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_294), .Y(n_357) );
BUFx4f_ASAP7_75t_L g358 ( .A(n_293), .Y(n_358) );
AND2x4_ASAP7_75t_L g359 ( .A(n_293), .B(n_29), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_306), .B(n_216), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_278), .Y(n_361) );
OR2x6_ASAP7_75t_L g362 ( .A(n_347), .B(n_303), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_358), .B(n_300), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_344), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_359), .A2(n_288), .B1(n_291), .B2(n_306), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_344), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_358), .B(n_250), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_358), .B(n_250), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_330), .B(n_295), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_361), .Y(n_370) );
CKINVDCx11_ASAP7_75t_R g371 ( .A(n_336), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_326), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_326), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_359), .A2(n_257), .B1(n_261), .B2(n_240), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_347), .B(n_305), .Y(n_375) );
CKINVDCx6p67_ASAP7_75t_R g376 ( .A(n_347), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_310), .B(n_304), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g379 ( .A(n_339), .B(n_291), .C(n_258), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_312), .Y(n_381) );
INVx2_ASAP7_75t_SL g382 ( .A(n_325), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_318), .Y(n_383) );
NOR2xp33_ASAP7_75t_R g384 ( .A(n_355), .B(n_240), .Y(n_384) );
NOR2xp33_ASAP7_75t_R g385 ( .A(n_355), .B(n_249), .Y(n_385) );
OR2x6_ASAP7_75t_L g386 ( .A(n_359), .B(n_303), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_329), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_323), .A2(n_252), .B1(n_255), .B2(n_251), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_334), .A2(n_273), .B1(n_264), .B2(n_246), .C(n_267), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_310), .B(n_282), .Y(n_390) );
AOI21x1_ASAP7_75t_L g391 ( .A1(n_360), .A2(n_259), .B(n_276), .Y(n_391) );
INVx3_ASAP7_75t_L g392 ( .A(n_342), .Y(n_392) );
INVx2_ASAP7_75t_SL g393 ( .A(n_325), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_310), .B(n_272), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_315), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_386), .B(n_309), .Y(n_396) );
OAI22xp5_ASAP7_75t_SL g397 ( .A1(n_374), .A2(n_243), .B1(n_336), .B2(n_273), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_372), .Y(n_398) );
BUFx12f_ASAP7_75t_L g399 ( .A(n_371), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_389), .A2(n_323), .B1(n_255), .B2(n_320), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_386), .B(n_290), .Y(n_401) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_386), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_389), .A2(n_323), .B1(n_332), .B2(n_349), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_370), .B(n_316), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_386), .B(n_292), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_372), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_373), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_365), .A2(n_349), .B1(n_360), .B2(n_348), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_365), .A2(n_357), .B1(n_350), .B2(n_322), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_379), .A2(n_276), .B(n_324), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_386), .A2(n_350), .B1(n_322), .B2(n_325), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_362), .A2(n_345), .B1(n_354), .B2(n_243), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_SL g415 ( .A1(n_392), .A2(n_345), .B(n_268), .C(n_351), .Y(n_415) );
AO31x2_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_268), .A3(n_285), .B(n_270), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_369), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_390), .B(n_269), .Y(n_419) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_362), .A2(n_246), .B1(n_238), .B2(n_256), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
OAI21x1_ASAP7_75t_L g422 ( .A1(n_391), .A2(n_324), .B(n_313), .Y(n_422) );
INVx4_ASAP7_75t_L g423 ( .A(n_376), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_424), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_397), .A2(n_388), .B1(n_363), .B2(n_362), .C(n_377), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_409), .A2(n_362), .B1(n_408), .B2(n_418), .Y(n_427) );
OA21x2_ASAP7_75t_L g428 ( .A1(n_422), .A2(n_404), .B(n_379), .Y(n_428) );
OAI33xp33_ASAP7_75t_L g429 ( .A1(n_397), .A2(n_377), .A3(n_380), .B1(n_256), .B2(n_395), .B3(n_381), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_414), .A2(n_400), .B1(n_403), .B2(n_418), .C(n_417), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_417), .B(n_380), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_423), .B(n_383), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_406), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_390), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_415), .A2(n_362), .B(n_387), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_407), .B(n_381), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_407), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_414), .A2(n_395), .B1(n_363), .B2(n_384), .C(n_394), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_410), .B(n_366), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_402), .Y(n_442) );
NAND3xp33_ASAP7_75t_SL g443 ( .A(n_420), .B(n_385), .C(n_366), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_423), .B(n_387), .Y(n_446) );
NOR4xp25_ASAP7_75t_SL g447 ( .A(n_423), .B(n_376), .C(n_346), .D(n_364), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_423), .A2(n_394), .B1(n_378), .B2(n_364), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_424), .Y(n_449) );
NOR2xp33_ASAP7_75t_R g450 ( .A(n_399), .B(n_364), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
OAI332xp33_ASAP7_75t_L g452 ( .A1(n_396), .A2(n_275), .A3(n_393), .B1(n_382), .B2(n_287), .B3(n_274), .C1(n_285), .C2(n_296), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
NAND3xp33_ASAP7_75t_L g454 ( .A(n_420), .B(n_353), .C(n_270), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_419), .B(n_378), .Y(n_455) );
OR2x2_ASAP7_75t_L g456 ( .A(n_402), .B(n_378), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_396), .B(n_378), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_411), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_401), .A2(n_367), .B1(n_368), .B2(n_375), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_401), .A2(n_367), .B1(n_368), .B2(n_375), .Y(n_460) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_440), .B(n_413), .C(n_401), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_434), .B(n_411), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_451), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_441), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_429), .A2(n_419), .B1(n_405), .B2(n_331), .C(n_382), .Y(n_465) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_437), .A2(n_412), .B(n_422), .Y(n_466) );
OAI33xp33_ASAP7_75t_L g467 ( .A1(n_433), .A2(n_296), .A3(n_279), .B1(n_421), .B2(n_206), .B3(n_174), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_426), .A2(n_405), .B1(n_375), .B2(n_419), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_431), .B(n_405), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_431), .B(n_421), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_451), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_433), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_436), .B(n_421), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_436), .B(n_375), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_430), .A2(n_393), .B1(n_399), .B2(n_392), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_434), .B(n_412), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_439), .B(n_412), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_441), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_452), .B(n_399), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_445), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_425), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_439), .B(n_412), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_444), .B(n_416), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_458), .B(n_422), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_446), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_444), .B(n_416), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_438), .B(n_416), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_445), .Y(n_490) );
AOI22xp5_ASAP7_75t_L g491 ( .A1(n_427), .A2(n_279), .B1(n_392), .B2(n_241), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g492 ( .A(n_454), .B(n_392), .C(n_183), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_SL g493 ( .A1(n_453), .A2(n_351), .B(n_416), .C(n_391), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
NOR2x1p5_ASAP7_75t_L g495 ( .A(n_443), .B(n_387), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_455), .A2(n_321), .B1(n_318), .B2(n_319), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_438), .Y(n_497) );
AOI33xp33_ASAP7_75t_L g498 ( .A1(n_459), .A2(n_174), .A3(n_237), .B1(n_208), .B2(n_217), .B3(n_319), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_455), .B(n_416), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g500 ( .A(n_448), .B(n_235), .C(n_183), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_428), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_442), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_442), .Y(n_503) );
INVx3_ASAP7_75t_L g504 ( .A(n_432), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_449), .B(n_416), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_428), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_456), .B(n_416), .Y(n_507) );
INVxp67_ASAP7_75t_L g508 ( .A(n_457), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_460), .B(n_356), .C(n_208), .D(n_351), .Y(n_509) );
OAI321xp33_ASAP7_75t_L g510 ( .A1(n_456), .A2(n_457), .A3(n_311), .B1(n_314), .B2(n_341), .C(n_343), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_428), .B(n_31), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_472), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_472), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_481), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_487), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_497), .B(n_464), .Y(n_516) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_505), .B(n_449), .Y(n_517) );
NOR3xp33_ASAP7_75t_L g518 ( .A(n_479), .B(n_449), .C(n_432), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_481), .Y(n_519) );
BUFx2_ASAP7_75t_L g520 ( .A(n_487), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_483), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_483), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_494), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_508), .B(n_432), .Y(n_524) );
NAND3xp33_ASAP7_75t_L g525 ( .A(n_482), .B(n_428), .C(n_447), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_497), .B(n_478), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_463), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_469), .B(n_446), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_470), .B(n_446), .Y(n_529) );
INVxp67_ASAP7_75t_L g530 ( .A(n_503), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_473), .B(n_450), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_463), .Y(n_532) );
INVxp67_ASAP7_75t_L g533 ( .A(n_503), .Y(n_533) );
INVxp67_ASAP7_75t_L g534 ( .A(n_502), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_461), .B(n_33), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_480), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_461), .B(n_36), .Y(n_537) );
NOR2xp67_ASAP7_75t_SL g538 ( .A(n_510), .B(n_352), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_499), .B(n_314), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_499), .B(n_50), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g541 ( .A(n_475), .B(n_327), .C(n_328), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_471), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_471), .B(n_318), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_507), .B(n_51), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_504), .B(n_57), .Y(n_545) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_480), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_462), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_507), .B(n_321), .Y(n_548) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_491), .A2(n_229), .B(n_191), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g550 ( .A1(n_492), .A2(n_341), .B(n_343), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_462), .Y(n_551) );
OAI31xp33_ASAP7_75t_L g552 ( .A1(n_468), .A2(n_337), .A3(n_327), .B(n_328), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_474), .B(n_58), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_490), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_490), .Y(n_555) );
INVx1_ASAP7_75t_SL g556 ( .A(n_504), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_486), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_486), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_489), .B(n_59), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_485), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_488), .B(n_321), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_476), .Y(n_562) );
NOR2x1_ASAP7_75t_L g563 ( .A(n_500), .B(n_337), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_509), .B(n_63), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_492), .A2(n_280), .B(n_286), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_476), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_477), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_504), .B(n_66), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_477), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_465), .B(n_69), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_516), .B(n_505), .Y(n_571) );
INVxp67_ASAP7_75t_SL g572 ( .A(n_523), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_560), .B(n_484), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_526), .B(n_505), .Y(n_574) );
AO22x1_ASAP7_75t_L g575 ( .A1(n_515), .A2(n_505), .B1(n_511), .B2(n_484), .Y(n_575) );
AOI32xp33_ASAP7_75t_L g576 ( .A1(n_535), .A2(n_511), .A3(n_506), .B1(n_496), .B2(n_501), .Y(n_576) );
OAI221xp5_ASAP7_75t_L g577 ( .A1(n_535), .A2(n_491), .B1(n_500), .B2(n_506), .C(n_501), .Y(n_577) );
OAI211xp5_ASAP7_75t_L g578 ( .A1(n_520), .A2(n_495), .B(n_352), .C(n_498), .Y(n_578) );
OAI21xp33_ASAP7_75t_L g579 ( .A1(n_537), .A2(n_493), .B(n_235), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_528), .B(n_466), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_512), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_518), .A2(n_495), .B1(n_467), .B2(n_466), .Y(n_582) );
OAI22xp33_ASAP7_75t_L g583 ( .A1(n_544), .A2(n_493), .B1(n_318), .B2(n_321), .Y(n_583) );
OAI211xp5_ASAP7_75t_SL g584 ( .A1(n_531), .A2(n_337), .B(n_328), .C(n_327), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_534), .A2(n_466), .B1(n_235), .B2(n_229), .C(n_183), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g586 ( .A1(n_515), .A2(n_352), .B1(n_317), .B2(n_313), .C1(n_308), .C2(n_286), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_558), .B(n_71), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_524), .B(n_547), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_540), .A2(n_342), .B1(n_352), .B2(n_340), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_L g590 ( .A1(n_537), .A2(n_308), .B(n_317), .C(n_79), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_551), .B(n_73), .Y(n_591) );
OAI322xp33_ASAP7_75t_L g592 ( .A1(n_534), .A2(n_203), .A3(n_235), .B1(n_183), .B2(n_191), .C1(n_229), .C2(n_74), .Y(n_592) );
AOI31xp33_ASAP7_75t_SL g593 ( .A1(n_518), .A2(n_193), .A3(n_215), .B(n_216), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_562), .B(n_191), .Y(n_594) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_517), .B(n_342), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_513), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_523), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_514), .Y(n_598) );
AOI221x1_ASAP7_75t_L g599 ( .A1(n_525), .A2(n_191), .B1(n_229), .B2(n_203), .C(n_340), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_517), .B(n_193), .Y(n_600) );
OAI21xp5_ASAP7_75t_SL g601 ( .A1(n_552), .A2(n_342), .B(n_340), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_519), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_521), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_566), .B(n_203), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_567), .B(n_203), .Y(n_605) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_564), .A2(n_352), .B(n_286), .C(n_249), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_557), .B(n_203), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_546), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_529), .B(n_329), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_570), .A2(n_329), .B1(n_333), .B2(n_340), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_556), .Y(n_611) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_545), .B(n_329), .Y(n_612) );
AOI21xp33_ASAP7_75t_SL g613 ( .A1(n_564), .A2(n_280), .B(n_286), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_522), .Y(n_614) );
OAI21xp33_ASAP7_75t_SL g615 ( .A1(n_563), .A2(n_333), .B(n_280), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g616 ( .A1(n_570), .A2(n_280), .B1(n_333), .B2(n_193), .C(n_215), .Y(n_616) );
OAI221xp5_ASAP7_75t_SL g617 ( .A1(n_539), .A2(n_193), .B1(n_215), .B2(n_333), .C(n_533), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g618 ( .A1(n_550), .A2(n_215), .B(n_549), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g619 ( .A1(n_541), .A2(n_538), .B(n_533), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_527), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_532), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_542), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_541), .A2(n_530), .B(n_545), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g624 ( .A(n_530), .B(n_568), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_580), .B(n_569), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_594), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_581), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_588), .B(n_546), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_571), .B(n_536), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_596), .Y(n_630) );
NOR3xp33_ASAP7_75t_SL g631 ( .A(n_619), .B(n_548), .C(n_561), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_574), .B(n_536), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_598), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_573), .B(n_602), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_608), .B(n_554), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_597), .B(n_555), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_603), .B(n_559), .Y(n_637) );
NOR4xp25_ASAP7_75t_SL g638 ( .A(n_601), .B(n_565), .C(n_543), .D(n_553), .Y(n_638) );
AOI21xp5_ASAP7_75t_SL g639 ( .A1(n_623), .A2(n_618), .B(n_578), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_614), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_611), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_620), .B(n_622), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g643 ( .A(n_595), .B(n_612), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_621), .B(n_572), .Y(n_644) );
OAI222xp33_ASAP7_75t_L g645 ( .A1(n_576), .A2(n_624), .B1(n_577), .B2(n_582), .C1(n_617), .C2(n_616), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_594), .Y(n_646) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_600), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_604), .Y(n_648) );
INVx2_ASAP7_75t_SL g649 ( .A(n_575), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_604), .B(n_605), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_605), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_585), .B(n_607), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_587), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_587), .B(n_591), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_577), .B(n_609), .Y(n_655) );
XNOR2xp5_ASAP7_75t_L g656 ( .A(n_616), .B(n_610), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_615), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_579), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_585), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_593), .Y(n_660) );
NOR2xp33_ASAP7_75t_R g661 ( .A(n_584), .B(n_589), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_628), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_644), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_627), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_641), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_655), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_650), .B(n_583), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_645), .A2(n_590), .B(n_613), .C(n_592), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g669 ( .A1(n_649), .A2(n_606), .B(n_599), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_659), .A2(n_586), .B1(n_656), .B2(n_652), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_642), .B(n_634), .Y(n_672) );
AOI211xp5_ASAP7_75t_L g673 ( .A1(n_639), .A2(n_649), .B(n_643), .C(n_660), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_630), .Y(n_674) );
XOR2x2_ASAP7_75t_L g675 ( .A(n_656), .B(n_654), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_630), .B(n_640), .Y(n_676) );
AOI32xp33_ASAP7_75t_L g677 ( .A1(n_657), .A2(n_659), .A3(n_652), .B1(n_625), .B2(n_629), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_633), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_633), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_647), .Y(n_680) );
INVx1_ASAP7_75t_SL g681 ( .A(n_629), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_640), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_666), .B(n_650), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g684 ( .A1(n_670), .A2(n_631), .B1(n_657), .B2(n_653), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_676), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_673), .A2(n_639), .B(n_638), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_665), .B(n_646), .Y(n_687) );
AO22x1_ASAP7_75t_L g688 ( .A1(n_672), .A2(n_658), .B1(n_637), .B2(n_653), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_668), .A2(n_638), .B(n_658), .Y(n_689) );
NOR3xp33_ASAP7_75t_L g690 ( .A(n_669), .B(n_646), .C(n_651), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_676), .Y(n_691) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_670), .B(n_637), .Y(n_692) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_677), .B(n_661), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_666), .B(n_625), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_664), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_681), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g697 ( .A1(n_672), .A2(n_632), .B1(n_651), .B2(n_626), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g698 ( .A1(n_663), .A2(n_635), .B1(n_636), .B2(n_626), .C(n_648), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_667), .A2(n_626), .B(n_648), .C(n_636), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_671), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_674), .A2(n_679), .B1(n_682), .B2(n_678), .C(n_662), .Y(n_701) );
NAND4xp75_ASAP7_75t_L g702 ( .A(n_675), .B(n_649), .C(n_631), .D(n_643), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_692), .B(n_684), .Y(n_703) );
CKINVDCx12_ASAP7_75t_R g704 ( .A(n_680), .Y(n_704) );
AOI22xp33_ASAP7_75t_R g705 ( .A1(n_702), .A2(n_689), .B1(n_684), .B2(n_693), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_686), .A2(n_690), .B1(n_688), .B2(n_687), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_687), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_707), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_703), .B(n_699), .C(n_697), .D(n_694), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_706), .A2(n_685), .B1(n_691), .B2(n_683), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_708), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_710), .Y(n_712) );
INVxp33_ASAP7_75t_SL g713 ( .A(n_711), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_711), .Y(n_714) );
AOI322xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_712), .A3(n_705), .B1(n_696), .B2(n_709), .C1(n_704), .C2(n_698), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_713), .B1(n_701), .B2(n_700), .C(n_695), .Y(n_716) );
endmodule