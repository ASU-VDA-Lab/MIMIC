module fake_jpeg_19721_n_344 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_344);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_344;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx24_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_39),
.Y(n_65)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_29),
.B1(n_34),
.B2(n_21),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_29),
.B1(n_34),
.B2(n_21),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_52),
.B1(n_66),
.B2(n_36),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_17),
.B1(n_33),
.B2(n_23),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_41),
.B(n_22),
.Y(n_63)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_63),
.B(n_42),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_68),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_72),
.Y(n_101)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_73),
.B(n_88),
.Y(n_122)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_61),
.A2(n_48),
.B1(n_47),
.B2(n_41),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_96),
.B1(n_48),
.B2(n_44),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_82),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_85),
.B(n_86),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_90),
.B1(n_92),
.B2(n_37),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

CKINVDCx6p67_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_42),
.Y(n_94)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_97),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_98),
.B(n_25),
.Y(n_131)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_104),
.A2(n_120),
.B1(n_124),
.B2(n_128),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_113),
.B1(n_68),
.B2(n_90),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_114),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_43),
.B1(n_44),
.B2(n_37),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_45),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_23),
.B1(n_20),
.B2(n_17),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_45),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_38),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_44),
.B1(n_45),
.B2(n_43),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_94),
.A2(n_45),
.B(n_38),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_28),
.B1(n_20),
.B2(n_32),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_131),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_93),
.C(n_89),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_142),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_121),
.B(n_116),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_138),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_35),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_120),
.B1(n_127),
.B2(n_102),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_76),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_122),
.B(n_101),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_35),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_38),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_75),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_40),
.Y(n_191)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_152),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_100),
.B1(n_97),
.B2(n_71),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_154),
.A2(n_42),
.B1(n_40),
.B2(n_95),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_25),
.B1(n_27),
.B2(n_26),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_27),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_35),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_158),
.A2(n_38),
.B(n_42),
.Y(n_182)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_159),
.A2(n_123),
.B1(n_109),
.B2(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_35),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_170),
.B1(n_175),
.B2(n_177),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_114),
.B1(n_118),
.B2(n_102),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_169),
.B1(n_174),
.B2(n_181),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_153),
.A2(n_105),
.B1(n_131),
.B2(n_115),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_125),
.B1(n_130),
.B2(n_109),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_146),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_171),
.B(n_24),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_185),
.B(n_191),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_157),
.A2(n_105),
.B1(n_126),
.B2(n_101),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_126),
.B1(n_124),
.B2(n_129),
.Y(n_175)
);

AO22x2_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_129),
.B1(n_69),
.B2(n_111),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_183),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_134),
.A2(n_111),
.B1(n_116),
.B2(n_132),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_142),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_132),
.B1(n_12),
.B2(n_2),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_151),
.B(n_148),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_140),
.A2(n_40),
.B(n_95),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_176),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_189),
.B(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_195),
.B(n_202),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_196),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_166),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_140),
.B1(n_144),
.B2(n_158),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_200),
.A2(n_216),
.B1(n_183),
.B2(n_176),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_163),
.B(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_203),
.B(n_206),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_209),
.B(n_213),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_189),
.B(n_136),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_207),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_210),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_185),
.B(n_174),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_150),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_212),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_173),
.A2(n_152),
.B(n_147),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_173),
.A2(n_159),
.B(n_19),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_217),
.B(n_221),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_222),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_190),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_9),
.B(n_13),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_219),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_31),
.C(n_30),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_181),
.C(n_168),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_167),
.A2(n_0),
.B(n_1),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_4),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_228),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_178),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_237),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_246),
.C(n_214),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_176),
.B1(n_169),
.B2(n_162),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_227),
.A2(n_242),
.B1(n_201),
.B2(n_221),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_176),
.C(n_31),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_233),
.Y(n_264)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_198),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_24),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_0),
.B1(n_1),
.B2(n_12),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_199),
.B1(n_204),
.B2(n_216),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_204),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_222),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_220),
.B(n_4),
.C(n_6),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_205),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_247),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_257),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_262),
.C(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_200),
.Y(n_259)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_260),
.A2(n_267),
.B1(n_224),
.B2(n_227),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_231),
.B1(n_248),
.B2(n_211),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_192),
.C(n_209),
.Y(n_262)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

INVx11_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_266),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_226),
.B(n_198),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_234),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_212),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_270),
.B(n_225),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_271),
.A2(n_252),
.B1(n_263),
.B2(n_254),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_274),
.B1(n_285),
.B2(n_261),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_229),
.B(n_230),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_242),
.B1(n_201),
.B2(n_202),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_276),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_229),
.B(n_230),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_12),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_260),
.A2(n_194),
.B1(n_207),
.B2(n_232),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_275),
.Y(n_294)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_262),
.C(n_258),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_292),
.C(n_295),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_270),
.C(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_294),
.B(n_297),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_264),
.C(n_194),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_298),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_246),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_218),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_252),
.B(n_219),
.Y(n_299)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_236),
.C(n_217),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_295),
.C(n_293),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_280),
.Y(n_306)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_289),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_306),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_284),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_309),
.B(n_310),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_279),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_292),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_289),
.C(n_284),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_288),
.C(n_8),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_305),
.A2(n_287),
.B(n_281),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_316),
.A2(n_302),
.B1(n_300),
.B2(n_282),
.Y(n_318)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_301),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_319),
.B(n_10),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_325),
.C(n_311),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_315),
.B(n_288),
.Y(n_321)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_321),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_308),
.A2(n_313),
.B1(n_307),
.B2(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_324),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_317),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_312),
.B(n_311),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_328),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_333),
.Y(n_335)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_325),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_331),
.Y(n_336)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_334),
.C(n_320),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_330),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_330),
.B(n_335),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_324),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_329),
.B(n_323),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_10),
.Y(n_344)
);


endmodule