module fake_jpeg_4654_n_16 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_16);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_16;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_7;

CKINVDCx5p33_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_0),
.Y(n_9)
);

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_8),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_10)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_10),
.A2(n_11),
.B1(n_8),
.B2(n_7),
.Y(n_13)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_9),
.B(n_7),
.Y(n_11)
);

CKINVDCx16_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

AO221x1_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_13),
.B1(n_0),
.B2(n_1),
.C(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_14),
.B(n_13),
.Y(n_15)
);

O2A1O1Ixp33_ASAP7_75t_SL g16 ( 
.A1(n_15),
.A2(n_4),
.B(n_5),
.C(n_14),
.Y(n_16)
);


endmodule