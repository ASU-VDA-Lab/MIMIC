module fake_netlist_6_3228_n_1405 (n_52, n_1, n_91, n_326, n_256, n_209, n_63, n_223, n_278, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_125, n_168, n_297, n_77, n_106, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_78, n_84, n_142, n_143, n_180, n_62, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_280, n_287, n_65, n_230, n_141, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_111, n_314, n_35, n_183, n_79, n_338, n_56, n_119, n_235, n_147, n_191, n_39, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_189, n_213, n_294, n_302, n_129, n_197, n_11, n_137, n_17, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_9, n_107, n_6, n_14, n_89, n_103, n_272, n_185, n_69, n_293, n_31, n_334, n_53, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_166, n_184, n_216, n_83, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_231, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_317, n_149, n_90, n_24, n_54, n_328, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_315, n_64, n_288, n_135, n_165, n_259, n_177, n_295, n_190, n_262, n_187, n_60, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1405);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_63;
input n_223;
input n_278;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_125;
input n_168;
input n_297;
input n_77;
input n_106;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_78;
input n_84;
input n_142;
input n_143;
input n_180;
input n_62;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_280;
input n_287;
input n_65;
input n_230;
input n_141;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_111;
input n_314;
input n_35;
input n_183;
input n_79;
input n_338;
input n_56;
input n_119;
input n_235;
input n_147;
input n_191;
input n_39;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_189;
input n_213;
input n_294;
input n_302;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_103;
input n_272;
input n_185;
input n_69;
input n_293;
input n_31;
input n_334;
input n_53;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_166;
input n_184;
input n_216;
input n_83;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_231;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_317;
input n_149;
input n_90;
input n_24;
input n_54;
input n_328;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_259;
input n_177;
input n_295;
input n_190;
input n_262;
input n_187;
input n_60;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1405;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1370;
wire n_369;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_1393;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_606;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_1052;
wire n_462;
wire n_1033;
wire n_1296;
wire n_694;
wire n_1294;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1384;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_1368;
wire n_958;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_1382;
wire n_1372;
wire n_505;
wire n_1339;
wire n_537;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_463;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1316;
wire n_1287;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1272;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_482;
wire n_934;
wire n_420;
wire n_1341;
wire n_394;
wire n_942;
wire n_543;
wire n_1271;
wire n_1355;
wire n_1225;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_1343;
wire n_548;
wire n_833;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_1248;
wire n_902;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_591;
wire n_1377;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1324;
wire n_1399;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_1028;
wire n_576;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_1311;
wire n_670;
wire n_1089;
wire n_1365;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_160),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_45),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_78),
.Y(n_342)
);

BUFx2_ASAP7_75t_L g343 ( 
.A(n_313),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_194),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_34),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_252),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_235),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_190),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_305),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_32),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_291),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_212),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_175),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_155),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_258),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_185),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_323),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_329),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_213),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_146),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_196),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_82),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_36),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_95),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_328),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_333),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_263),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_86),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_214),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_128),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_24),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_136),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_79),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_246),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_327),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_278),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_96),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_173),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_22),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_311),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_295),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_195),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_88),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_73),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_147),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_26),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_158),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_44),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_25),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_253),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_145),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_234),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_331),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_207),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_132),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_285),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_317),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_138),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_276),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_123),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_334),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_116),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_264),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_218),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_238),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_26),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_236),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_71),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_1),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_23),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_74),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_319),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_49),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_188),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_259),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_270),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_204),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_191),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_100),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_172),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_23),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_245),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_104),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_83),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_247),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_15),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_22),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_34),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_85),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_60),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_7),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_162),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_14),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_168),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_27),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_66),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_169),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_325),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_42),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_76),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_144),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_299),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_261),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_151),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_55),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_121),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_89),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_61),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_54),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_198),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_93),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_208),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_108),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_81),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_220),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_332),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_240),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_326),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_64),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_99),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_20),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_135),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_154),
.Y(n_468)
);

BUFx10_ASAP7_75t_L g469 ( 
.A(n_255),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_337),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_39),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_3),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_307),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_260),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_117),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_293),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_227),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_164),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_233),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_48),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_183),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_51),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_321),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_186),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_280),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_256),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_103),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_25),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_231),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_14),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_152),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_38),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_68),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_254),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_39),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_17),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_3),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_308),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_48),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_57),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_141),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_49),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_304),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_273),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_189),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_244),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_90),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_10),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_300),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_69),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_306),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_314),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g513 ( 
.A(n_274),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_271),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_113),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_125),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_139),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_118),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_106),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_322),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_102),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_222),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_267),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_210),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_10),
.Y(n_525)
);

INVx4_ASAP7_75t_R g526 ( 
.A(n_266),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_114),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_463),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_350),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_350),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_463),
.B(n_0),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_350),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_350),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_374),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_358),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_466),
.B(n_0),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_374),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_374),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_358),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_343),
.B(n_1),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_476),
.B(n_2),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_374),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_508),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_358),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_466),
.B(n_2),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_358),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_398),
.Y(n_547)
);

INVx5_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

BUFx8_ASAP7_75t_SL g549 ( 
.A(n_382),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_429),
.B(n_4),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_398),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_373),
.B(n_4),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_508),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_476),
.B(n_5),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_508),
.Y(n_556)
);

AND2x6_ASAP7_75t_L g557 ( 
.A(n_416),
.B(n_65),
.Y(n_557)
);

INVx5_ASAP7_75t_L g558 ( 
.A(n_398),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_416),
.B(n_5),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_371),
.B(n_6),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_357),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_487),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_341),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_433),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_391),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_513),
.B(n_6),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_433),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_487),
.B(n_7),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_377),
.B(n_8),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_400),
.B(n_8),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_357),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_527),
.B(n_9),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_340),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_415),
.Y(n_575)
);

BUFx8_ASAP7_75t_L g576 ( 
.A(n_471),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_377),
.B(n_9),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_430),
.B(n_11),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_430),
.B(n_67),
.Y(n_579)
);

XNOR2x2_ASAP7_75t_L g580 ( 
.A(n_418),
.B(n_11),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_342),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_357),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_403),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_394),
.B(n_12),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_514),
.B(n_12),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_494),
.B(n_403),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_514),
.B(n_70),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_403),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_461),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_347),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_426),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_339),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_431),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_376),
.B(n_13),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_432),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_461),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_346),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_461),
.Y(n_598)
);

INVx2_ASAP7_75t_SL g599 ( 
.A(n_469),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_469),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_469),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_512),
.B(n_13),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_450),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_397),
.B(n_15),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_454),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_414),
.B(n_378),
.Y(n_606)
);

BUFx12f_ASAP7_75t_L g607 ( 
.A(n_512),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_512),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_344),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_345),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_R g611 ( 
.A(n_402),
.B(n_445),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_526),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_423),
.B(n_16),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_472),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_349),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_352),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_366),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_389),
.Y(n_619)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_500),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_392),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_348),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_353),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_351),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_410),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_525),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_356),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_442),
.B(n_16),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_574),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_606),
.A2(n_451),
.B1(n_473),
.B2(n_470),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_534),
.Y(n_631)
);

AND2x2_ASAP7_75t_SL g632 ( 
.A(n_552),
.B(n_367),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_538),
.Y(n_633)
);

OA22x2_ASAP7_75t_L g634 ( 
.A1(n_586),
.A2(n_435),
.B1(n_436),
.B2(n_413),
.Y(n_634)
);

OA22x2_ASAP7_75t_L g635 ( 
.A1(n_599),
.A2(n_440),
.B1(n_444),
.B2(n_438),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_561),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_596),
.B(n_478),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_581),
.B(n_369),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_561),
.Y(n_639)
);

OAI22xp33_ASAP7_75t_L g640 ( 
.A1(n_552),
.A2(n_453),
.B1(n_490),
.B2(n_488),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_530),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_543),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_540),
.A2(n_451),
.B1(n_489),
.B2(n_483),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_600),
.B(n_608),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_566),
.A2(n_511),
.B1(n_520),
.B2(n_504),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_L g646 ( 
.A1(n_536),
.A2(n_596),
.B1(n_589),
.B2(n_559),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_537),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_536),
.A2(n_492),
.B1(n_497),
.B2(n_496),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_612),
.B(n_523),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_612),
.B(n_589),
.Y(n_650)
);

NAND3x1_ASAP7_75t_L g651 ( 
.A(n_602),
.B(n_387),
.C(n_386),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_530),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_545),
.A2(n_502),
.B1(n_499),
.B2(n_495),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_612),
.B(n_563),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_354),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_559),
.A2(n_482),
.B1(n_407),
.B2(n_409),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_550),
.A2(n_359),
.B1(n_360),
.B2(n_355),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_530),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_604),
.A2(n_421),
.B1(n_434),
.B2(n_388),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_537),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

AO22x2_ASAP7_75t_L g662 ( 
.A1(n_531),
.A2(n_447),
.B1(n_458),
.B2(n_441),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_533),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_590),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_L g665 ( 
.A1(n_604),
.A2(n_462),
.B1(n_464),
.B2(n_460),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_533),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_560),
.A2(n_362),
.B1(n_363),
.B2(n_361),
.Y(n_667)
);

OAI22xp33_ASAP7_75t_L g668 ( 
.A1(n_569),
.A2(n_477),
.B1(n_479),
.B2(n_467),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_570),
.A2(n_365),
.B1(n_368),
.B2(n_364),
.Y(n_669)
);

AO22x2_ASAP7_75t_L g670 ( 
.A1(n_531),
.A2(n_486),
.B1(n_493),
.B2(n_484),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_542),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_611),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_583),
.B(n_509),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_613),
.A2(n_372),
.B1(n_375),
.B2(n_370),
.Y(n_674)
);

OA22x2_ASAP7_75t_L g675 ( 
.A1(n_620),
.A2(n_519),
.B1(n_517),
.B2(n_380),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_553),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_379),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_569),
.A2(n_383),
.B1(n_384),
.B2(n_381),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_561),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_616),
.B(n_385),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_625),
.A2(n_393),
.B1(n_395),
.B2(n_390),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_553),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_584),
.A2(n_399),
.B1(n_401),
.B2(n_396),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_555),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_572),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_628),
.A2(n_405),
.B1(n_406),
.B2(n_404),
.Y(n_686)
);

AO22x2_ASAP7_75t_L g687 ( 
.A1(n_541),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_621),
.A2(n_411),
.B1(n_412),
.B2(n_408),
.Y(n_688)
);

OAI22xp33_ASAP7_75t_L g689 ( 
.A1(n_572),
.A2(n_419),
.B1(n_420),
.B2(n_417),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_607),
.B(n_18),
.Y(n_690)
);

AND2x2_ASAP7_75t_SL g691 ( 
.A(n_573),
.B(n_19),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_SL g692 ( 
.A1(n_594),
.A2(n_424),
.B1(n_425),
.B2(n_422),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_541),
.A2(n_428),
.B1(n_437),
.B2(n_427),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_555),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_622),
.B(n_524),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_528),
.B(n_439),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_533),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_572),
.B(n_443),
.Y(n_698)
);

OA22x2_ASAP7_75t_L g699 ( 
.A1(n_565),
.A2(n_448),
.B1(n_449),
.B2(n_446),
.Y(n_699)
);

OAI22xp33_ASAP7_75t_L g700 ( 
.A1(n_582),
.A2(n_455),
.B1(n_456),
.B2(n_452),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_582),
.B(n_457),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_535),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_554),
.A2(n_568),
.B1(n_578),
.B2(n_577),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_SL g704 ( 
.A1(n_554),
.A2(n_522),
.B1(n_521),
.B2(n_518),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_598),
.A2(n_516),
.B1(n_515),
.B2(n_510),
.Y(n_705)
);

OR2x6_ASAP7_75t_L g706 ( 
.A(n_601),
.B(n_20),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_556),
.Y(n_707)
);

AO22x2_ASAP7_75t_L g708 ( 
.A1(n_568),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_577),
.A2(n_507),
.B1(n_506),
.B2(n_505),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_562),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_575),
.B(n_21),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_582),
.B(n_459),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_694),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_694),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_641),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_641),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_653),
.B(n_624),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_654),
.B(n_588),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_633),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_702),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_703),
.B(n_627),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_702),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_650),
.B(n_529),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_638),
.B(n_588),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_652),
.Y(n_725)
);

INVxp33_ASAP7_75t_L g726 ( 
.A(n_630),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_658),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_663),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_666),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_697),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_647),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_672),
.Y(n_732)
);

XOR2xp5_ASAP7_75t_L g733 ( 
.A(n_645),
.B(n_643),
.Y(n_733)
);

CKINVDCx20_ASAP7_75t_R g734 ( 
.A(n_629),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_660),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_661),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_671),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_676),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_682),
.Y(n_739)
);

CKINVDCx16_ASAP7_75t_R g740 ( 
.A(n_644),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_684),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_703),
.B(n_627),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_707),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_631),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_649),
.B(n_696),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_637),
.B(n_529),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_642),
.Y(n_747)
);

XOR2xp5_ASAP7_75t_L g748 ( 
.A(n_664),
.B(n_465),
.Y(n_748)
);

INVx2_ASAP7_75t_SL g749 ( 
.A(n_632),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_710),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_710),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_699),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_655),
.Y(n_753)
);

INVxp33_ASAP7_75t_L g754 ( 
.A(n_680),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_675),
.B(n_588),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_662),
.Y(n_756)
);

XOR2xp5_ASAP7_75t_L g757 ( 
.A(n_634),
.B(n_468),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_662),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_670),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_670),
.Y(n_760)
);

AND2x2_ASAP7_75t_SL g761 ( 
.A(n_691),
.B(n_578),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_698),
.B(n_529),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_711),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_R g764 ( 
.A(n_644),
.B(n_585),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_711),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_695),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_701),
.Y(n_767)
);

XNOR2xp5_ASAP7_75t_L g768 ( 
.A(n_656),
.B(n_580),
.Y(n_768)
);

XOR2x2_ASAP7_75t_L g769 ( 
.A(n_635),
.B(n_549),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_712),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_659),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_648),
.B(n_562),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_646),
.B(n_640),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_693),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_687),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_636),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_687),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_708),
.B(n_585),
.Y(n_778)
);

XOR2xp5_ASAP7_75t_L g779 ( 
.A(n_705),
.B(n_474),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_708),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_681),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_639),
.B(n_564),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_706),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_678),
.B(n_562),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_679),
.B(n_564),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_709),
.A2(n_557),
.B(n_579),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_685),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_685),
.B(n_618),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_651),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_706),
.Y(n_790)
);

CKINVDCx16_ASAP7_75t_R g791 ( 
.A(n_673),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_692),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_688),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_674),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_686),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_677),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_667),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_669),
.B(n_657),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_673),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_668),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_690),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_767),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_721),
.B(n_593),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_721),
.B(n_603),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_744),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_713),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_767),
.B(n_557),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_742),
.B(n_614),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_713),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_742),
.B(n_617),
.Y(n_810)
);

AND2x2_ASAP7_75t_SL g811 ( 
.A(n_761),
.B(n_557),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_764),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_714),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_745),
.B(n_591),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_764),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_714),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_719),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_734),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_736),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_782),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_796),
.B(n_591),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_744),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_719),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_766),
.B(n_557),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_796),
.B(n_595),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_771),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_704),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_736),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_741),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_741),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_752),
.B(n_595),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_731),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_778),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_749),
.B(n_605),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_749),
.B(n_605),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_724),
.B(n_770),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_784),
.B(n_665),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_735),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_734),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_747),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_737),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_738),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_761),
.B(n_626),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_739),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_754),
.B(n_689),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_756),
.B(n_626),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_743),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_725),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_727),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_728),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_729),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_730),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_715),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_784),
.B(n_683),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_758),
.B(n_571),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_716),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_772),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_786),
.A2(n_700),
.B(n_587),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_753),
.B(n_571),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_773),
.B(n_571),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_720),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_793),
.B(n_579),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_773),
.B(n_567),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_722),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_782),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_785),
.Y(n_866)
);

HB1xp67_ASAP7_75t_L g867 ( 
.A(n_789),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_785),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_797),
.B(n_579),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_754),
.B(n_567),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_794),
.B(n_579),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_795),
.B(n_587),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_763),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_750),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_781),
.B(n_717),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_798),
.A2(n_587),
.B(n_556),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_787),
.Y(n_877)
);

AND2x2_ASAP7_75t_SL g878 ( 
.A(n_798),
.B(n_587),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_787),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_800),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_789),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_778),
.B(n_618),
.Y(n_882)
);

AND2x2_ASAP7_75t_SL g883 ( 
.A(n_774),
.B(n_592),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_759),
.B(n_690),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_778),
.B(n_618),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_760),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_755),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_746),
.B(n_619),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_755),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_792),
.B(n_718),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_763),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_778),
.B(n_775),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_777),
.B(n_619),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_762),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_723),
.A2(n_481),
.B(n_475),
.Y(n_895)
);

AND2x2_ASAP7_75t_SL g896 ( 
.A(n_780),
.B(n_592),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_776),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_860),
.B(n_768),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_802),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_875),
.B(n_726),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_884),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_834),
.B(n_726),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_887),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_833),
.B(n_790),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_809),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_809),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_834),
.B(n_733),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_860),
.B(n_765),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_833),
.B(n_790),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_806),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_806),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_816),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_SL g913 ( 
.A(n_811),
.B(n_732),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_SL g914 ( 
.A(n_811),
.B(n_878),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_833),
.B(n_783),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_843),
.B(n_748),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_889),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_812),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_897),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_818),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_802),
.Y(n_921)
);

OR2x2_ASAP7_75t_L g922 ( 
.A(n_843),
.B(n_740),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_892),
.B(n_801),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_835),
.B(n_776),
.Y(n_924)
);

OR2x2_ASAP7_75t_L g925 ( 
.A(n_857),
.B(n_801),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_879),
.Y(n_926)
);

BUFx3_ASAP7_75t_L g927 ( 
.A(n_889),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_863),
.B(n_757),
.Y(n_928)
);

NAND2x1p5_ASAP7_75t_L g929 ( 
.A(n_897),
.B(n_751),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_879),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_867),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_863),
.B(n_779),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_816),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_878),
.Y(n_934)
);

BUFx5_ASAP7_75t_L g935 ( 
.A(n_877),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_813),
.Y(n_936)
);

OR2x6_ASAP7_75t_L g937 ( 
.A(n_892),
.B(n_732),
.Y(n_937)
);

INVx4_ASAP7_75t_L g938 ( 
.A(n_897),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_897),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_880),
.B(n_592),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_873),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_897),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_815),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_837),
.B(n_609),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_881),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_866),
.B(n_485),
.Y(n_946)
);

BUFx2_ASAP7_75t_L g947 ( 
.A(n_884),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_877),
.Y(n_948)
);

NAND2x1_ASAP7_75t_SL g949 ( 
.A(n_882),
.B(n_769),
.Y(n_949)
);

BUFx8_ASAP7_75t_SL g950 ( 
.A(n_884),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_802),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_802),
.Y(n_952)
);

HB1xp67_ASAP7_75t_L g953 ( 
.A(n_826),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_883),
.B(n_802),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_835),
.B(n_791),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_813),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_883),
.B(n_821),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_891),
.B(n_799),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_846),
.B(n_799),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_886),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_854),
.B(n_619),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_828),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_821),
.B(n_609),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_825),
.B(n_609),
.Y(n_964)
);

OR2x2_ASAP7_75t_L g965 ( 
.A(n_839),
.B(n_769),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_870),
.B(n_610),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_813),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_870),
.B(n_610),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_846),
.B(n_788),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_944),
.B(n_825),
.Y(n_970)
);

CKINVDCx8_ASAP7_75t_R g971 ( 
.A(n_947),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_944),
.B(n_814),
.Y(n_972)
);

CKINVDCx14_ASAP7_75t_R g973 ( 
.A(n_920),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_951),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_901),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_948),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_905),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_951),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_919),
.Y(n_979)
);

CKINVDCx16_ASAP7_75t_R g980 ( 
.A(n_937),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_918),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_934),
.B(n_814),
.Y(n_982)
);

INVx6_ASAP7_75t_L g983 ( 
.A(n_958),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_925),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_919),
.Y(n_985)
);

INVx2_ASAP7_75t_SL g986 ( 
.A(n_903),
.Y(n_986)
);

INVx8_ASAP7_75t_L g987 ( 
.A(n_923),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_919),
.Y(n_988)
);

BUFx2_ASAP7_75t_SL g989 ( 
.A(n_958),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_951),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_939),
.Y(n_991)
);

INVx6_ASAP7_75t_SL g992 ( 
.A(n_937),
.Y(n_992)
);

OR2x6_ASAP7_75t_L g993 ( 
.A(n_937),
.B(n_820),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_950),
.Y(n_994)
);

INVx6_ASAP7_75t_L g995 ( 
.A(n_959),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_906),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_959),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_953),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_962),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_934),
.B(n_866),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_910),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_902),
.B(n_868),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_915),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_939),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_952),
.Y(n_1005)
);

INVx1_ASAP7_75t_SL g1006 ( 
.A(n_943),
.Y(n_1006)
);

BUFx2_ASAP7_75t_R g1007 ( 
.A(n_898),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_922),
.Y(n_1008)
);

BUFx2_ASAP7_75t_R g1009 ( 
.A(n_898),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_915),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_955),
.Y(n_1011)
);

BUFx12f_ASAP7_75t_L g1012 ( 
.A(n_923),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_924),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_923),
.B(n_846),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_952),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_907),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_939),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_904),
.B(n_803),
.Y(n_1018)
);

INVx1_ASAP7_75t_SL g1019 ( 
.A(n_908),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_917),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_926),
.Y(n_1021)
);

BUFx2_ASAP7_75t_SL g1022 ( 
.A(n_927),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_914),
.B(n_841),
.Y(n_1023)
);

BUFx2_ASAP7_75t_SL g1024 ( 
.A(n_942),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_952),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_SL g1026 ( 
.A(n_904),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_909),
.B(n_803),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_911),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_976),
.Y(n_1029)
);

AOI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_1016),
.A2(n_900),
.B1(n_932),
.B2(n_913),
.Y(n_1030)
);

CKINVDCx11_ASAP7_75t_R g1031 ( 
.A(n_971),
.Y(n_1031)
);

INVx6_ASAP7_75t_L g1032 ( 
.A(n_995),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_981),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1018),
.A2(n_932),
.B1(n_928),
.B2(n_845),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_979),
.Y(n_1035)
);

INVx6_ASAP7_75t_L g1036 ( 
.A(n_995),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_977),
.Y(n_1037)
);

OAI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_1016),
.A2(n_913),
.B1(n_914),
.B2(n_916),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_996),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_999),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_SL g1041 ( 
.A(n_992),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_980),
.A2(n_928),
.B1(n_1011),
.B2(n_973),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_1019),
.A2(n_957),
.B1(n_954),
.B2(n_908),
.Y(n_1043)
);

CKINVDCx20_ASAP7_75t_R g1044 ( 
.A(n_994),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_979),
.Y(n_1045)
);

INVx1_ASAP7_75t_SL g1046 ( 
.A(n_981),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1001),
.Y(n_1047)
);

CKINVDCx12_ASAP7_75t_R g1048 ( 
.A(n_993),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1028),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1021),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_1015),
.B(n_938),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1002),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1018),
.A2(n_890),
.B1(n_957),
.B2(n_858),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_997),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1013),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1013),
.B(n_1019),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_SL g1057 ( 
.A(n_992),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1027),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_982),
.B(n_966),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_1027),
.A2(n_909),
.B1(n_961),
.B2(n_941),
.Y(n_1060)
);

BUFx12f_ASAP7_75t_L g1061 ( 
.A(n_1012),
.Y(n_1061)
);

BUFx12f_ASAP7_75t_L g1062 ( 
.A(n_998),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1008),
.A2(n_827),
.B1(n_894),
.B2(n_804),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_982),
.B(n_968),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_979),
.Y(n_1065)
);

CKINVDCx11_ASAP7_75t_R g1066 ( 
.A(n_975),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_1000),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_SL g1068 ( 
.A1(n_1006),
.A2(n_965),
.B1(n_896),
.B2(n_945),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_972),
.B(n_868),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1000),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_1015),
.Y(n_1071)
);

INVx6_ASAP7_75t_L g1072 ( 
.A(n_983),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1006),
.B(n_804),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_1014),
.A2(n_894),
.B1(n_810),
.B2(n_808),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_974),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1014),
.A2(n_810),
.B1(n_808),
.B2(n_882),
.Y(n_1076)
);

OAI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_1023),
.A2(n_836),
.B1(n_931),
.B2(n_820),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_974),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_972),
.A2(n_859),
.B1(n_896),
.B2(n_865),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_993),
.A2(n_885),
.B1(n_893),
.B2(n_831),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_SL g1081 ( 
.A1(n_1022),
.A2(n_874),
.B1(n_859),
.B2(n_876),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_970),
.A2(n_824),
.B(n_807),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_970),
.B(n_963),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1050),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1030),
.A2(n_1007),
.B1(n_1009),
.B2(n_993),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_1071),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1030),
.A2(n_1009),
.B1(n_1007),
.B2(n_984),
.Y(n_1087)
);

OAI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_1063),
.A2(n_946),
.B(n_949),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1068),
.A2(n_838),
.B1(n_832),
.B2(n_963),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_1073),
.B(n_893),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_1055),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1068),
.A2(n_838),
.B1(n_832),
.B2(n_964),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1029),
.Y(n_1093)
);

BUFx2_ASAP7_75t_SL g1094 ( 
.A(n_1054),
.Y(n_1094)
);

OAI222xp33_ASAP7_75t_L g1095 ( 
.A1(n_1079),
.A2(n_1023),
.B1(n_964),
.B2(n_929),
.C1(n_986),
.C2(n_940),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1038),
.A2(n_842),
.B1(n_940),
.B2(n_987),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1034),
.A2(n_842),
.B1(n_987),
.B2(n_847),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1060),
.A2(n_874),
.B1(n_1026),
.B2(n_989),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1037),
.Y(n_1099)
);

NOR2x1_ASAP7_75t_R g1100 ( 
.A(n_1031),
.B(n_983),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1052),
.B(n_1020),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1059),
.A2(n_987),
.B1(n_844),
.B2(n_829),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_1041),
.A2(n_1026),
.B1(n_1003),
.B2(n_1010),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1039),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1064),
.A2(n_829),
.B1(n_830),
.B2(n_828),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1042),
.A2(n_960),
.B1(n_855),
.B2(n_938),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1053),
.A2(n_830),
.B1(n_852),
.B2(n_848),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1040),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1043),
.A2(n_1056),
.B1(n_1069),
.B2(n_1077),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1083),
.A2(n_848),
.B1(n_852),
.B2(n_840),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1058),
.B(n_885),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_1046),
.B(n_978),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_1046),
.B(n_831),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1067),
.A2(n_851),
.B1(n_850),
.B2(n_822),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1047),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1070),
.A2(n_850),
.B1(n_851),
.B2(n_805),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1049),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1048),
.A2(n_969),
.B1(n_831),
.B2(n_841),
.Y(n_1118)
);

OAI21xp5_ASAP7_75t_SL g1119 ( 
.A1(n_1081),
.A2(n_895),
.B(n_969),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_1066),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_1033),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1078),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1075),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1035),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_SL g1125 ( 
.A1(n_1057),
.A2(n_576),
.B1(n_960),
.B2(n_807),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1079),
.A2(n_960),
.B1(n_819),
.B2(n_849),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1071),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1035),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_1035),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_1045),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1076),
.B(n_855),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1045),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1074),
.A2(n_855),
.B1(n_871),
.B2(n_869),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1080),
.B(n_886),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_1032),
.B(n_856),
.Y(n_1135)
);

AOI222xp33_ASAP7_75t_L g1136 ( 
.A1(n_1061),
.A2(n_576),
.B1(n_864),
.B2(n_856),
.C1(n_872),
.C2(n_862),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1062),
.B(n_841),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_1072),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1045),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1065),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1072),
.A2(n_807),
.B1(n_1024),
.B2(n_935),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_SL g1142 ( 
.A1(n_1032),
.A2(n_935),
.B1(n_942),
.B2(n_841),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1036),
.B(n_841),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_1036),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1065),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1082),
.A2(n_819),
.B1(n_933),
.B2(n_912),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1093),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1088),
.A2(n_861),
.B1(n_864),
.B2(n_853),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1136),
.A2(n_861),
.B1(n_853),
.B2(n_823),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1087),
.A2(n_853),
.B1(n_823),
.B2(n_817),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1121),
.B(n_1065),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_SL g1152 ( 
.A1(n_1085),
.A2(n_1044),
.B1(n_1051),
.B2(n_942),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1089),
.A2(n_1092),
.B1(n_1097),
.B2(n_1131),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1089),
.A2(n_853),
.B1(n_817),
.B2(n_888),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1092),
.A2(n_853),
.B1(n_921),
.B2(n_899),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1097),
.A2(n_921),
.B1(n_899),
.B2(n_935),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1108),
.B(n_978),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1090),
.A2(n_935),
.B1(n_956),
.B2(n_936),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1096),
.A2(n_935),
.B1(n_967),
.B2(n_930),
.Y(n_1159)
);

OAI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1102),
.A2(n_1051),
.B1(n_1025),
.B2(n_1015),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1118),
.A2(n_1025),
.B1(n_1015),
.B2(n_990),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1096),
.A2(n_491),
.B1(n_501),
.B2(n_498),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1115),
.B(n_990),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1102),
.A2(n_503),
.B1(n_610),
.B2(n_615),
.Y(n_1164)
);

NAND3xp33_ASAP7_75t_L g1165 ( 
.A(n_1119),
.B(n_1125),
.C(n_1109),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1134),
.A2(n_623),
.B1(n_615),
.B2(n_1005),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1111),
.A2(n_1098),
.B1(n_1109),
.B2(n_1094),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1113),
.A2(n_623),
.B1(n_615),
.B2(n_1005),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1135),
.A2(n_623),
.B1(n_1017),
.B2(n_1004),
.Y(n_1169)
);

OAI211xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1101),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1103),
.A2(n_1025),
.B1(n_1017),
.B2(n_1004),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1099),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1106),
.A2(n_1137),
.B1(n_1138),
.B2(n_1143),
.Y(n_1173)
);

OAI222xp33_ASAP7_75t_L g1174 ( 
.A1(n_1110),
.A2(n_1126),
.B1(n_1107),
.B2(n_1114),
.C1(n_1116),
.C2(n_1141),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1133),
.A2(n_1017),
.B1(n_1004),
.B2(n_991),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1110),
.A2(n_1025),
.B1(n_991),
.B2(n_988),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1120),
.A2(n_991),
.B1(n_988),
.B2(n_985),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1107),
.A2(n_988),
.B1(n_985),
.B2(n_535),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1112),
.A2(n_985),
.B1(n_546),
.B2(n_551),
.Y(n_1179)
);

AOI222xp33_ASAP7_75t_L g1180 ( 
.A1(n_1100),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C1(n_31),
.C2(n_32),
.Y(n_1180)
);

AOI22xp33_ASAP7_75t_L g1181 ( 
.A1(n_1112),
.A2(n_546),
.B1(n_551),
.B2(n_535),
.Y(n_1181)
);

OAI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1091),
.A2(n_546),
.B1(n_551),
.B2(n_548),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1084),
.B(n_31),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1091),
.B(n_33),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_SL g1185 ( 
.A(n_1126),
.B(n_1104),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_SL g1186 ( 
.A1(n_1117),
.A2(n_558),
.B1(n_548),
.B2(n_547),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1105),
.A2(n_558),
.B1(n_548),
.B2(n_547),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1122),
.B(n_1123),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1105),
.A2(n_547),
.B1(n_544),
.B2(n_539),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1128),
.B(n_33),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1144),
.A2(n_558),
.B1(n_544),
.B2(n_539),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1143),
.A2(n_75),
.B(n_72),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1116),
.A2(n_544),
.B1(n_539),
.B2(n_532),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1095),
.A2(n_35),
.B(n_36),
.Y(n_1194)
);

OAI222xp33_ASAP7_75t_L g1195 ( 
.A1(n_1114),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C1(n_40),
.C2(n_41),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1146),
.Y(n_1196)
);

NAND3xp33_ASAP7_75t_L g1197 ( 
.A(n_1146),
.B(n_532),
.C(n_37),
.Y(n_1197)
);

AOI222xp33_ASAP7_75t_L g1198 ( 
.A1(n_1132),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.C1(n_43),
.C2(n_44),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1145),
.A2(n_532),
.B1(n_45),
.B2(n_46),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1140),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1124),
.B(n_47),
.Y(n_1201)
);

OAI221xp5_ASAP7_75t_SL g1202 ( 
.A1(n_1139),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.C(n_53),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_L g1203 ( 
.A(n_1142),
.B(n_1130),
.C(n_1129),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1086),
.A2(n_1127),
.B1(n_1130),
.B2(n_1129),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1086),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1165),
.B(n_1180),
.C(n_1198),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1194),
.A2(n_1127),
.B(n_1129),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1188),
.B(n_1129),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1188),
.B(n_1130),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_L g1210 ( 
.A(n_1202),
.B(n_1130),
.C(n_54),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1170),
.B(n_55),
.C(n_56),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_L g1212 ( 
.A(n_1205),
.B(n_56),
.C(n_57),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1153),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1147),
.B(n_1172),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1147),
.B(n_58),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1172),
.B(n_59),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1173),
.B(n_61),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_SL g1218 ( 
.A(n_1185),
.B(n_77),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_SL g1219 ( 
.A1(n_1149),
.A2(n_62),
.B(n_63),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1157),
.B(n_62),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1157),
.B(n_63),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1151),
.B(n_1167),
.Y(n_1222)
);

NAND3xp33_ASAP7_75t_L g1223 ( 
.A(n_1200),
.B(n_80),
.C(n_84),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1163),
.B(n_1184),
.Y(n_1224)
);

OAI221xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1199),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.C(n_94),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1195),
.B(n_97),
.C(n_98),
.Y(n_1226)
);

NAND3xp33_ASAP7_75t_L g1227 ( 
.A(n_1162),
.B(n_101),
.C(n_105),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1185),
.B(n_107),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1197),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.C(n_112),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1163),
.B(n_336),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1152),
.B(n_115),
.C(n_119),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1160),
.A2(n_120),
.B1(n_122),
.B2(n_124),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1196),
.B(n_126),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1196),
.B(n_127),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1161),
.B(n_1148),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1204),
.B(n_335),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1150),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1154),
.A2(n_133),
.B1(n_134),
.B2(n_137),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_1174),
.B(n_140),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1192),
.A2(n_142),
.B(n_143),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1183),
.B(n_148),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1190),
.B(n_149),
.Y(n_1242)
);

NAND4xp25_ASAP7_75t_L g1243 ( 
.A(n_1201),
.B(n_150),
.C(n_153),
.D(n_156),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1155),
.B(n_157),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1164),
.A2(n_159),
.B(n_161),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1175),
.B(n_163),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1203),
.B(n_1166),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1177),
.A2(n_165),
.B(n_166),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1169),
.B(n_167),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1159),
.B(n_1158),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1156),
.B(n_1171),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1176),
.B(n_170),
.Y(n_1252)
);

OR2x2_ASAP7_75t_L g1253 ( 
.A(n_1214),
.B(n_1168),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1208),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1224),
.B(n_1192),
.Y(n_1255)
);

NAND4xp75_ASAP7_75t_L g1256 ( 
.A(n_1218),
.B(n_1186),
.C(n_1182),
.D(n_1191),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1209),
.B(n_1179),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1206),
.A2(n_1178),
.B1(n_1189),
.B2(n_1187),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1216),
.Y(n_1259)
);

NOR3xp33_ASAP7_75t_L g1260 ( 
.A(n_1218),
.B(n_1181),
.C(n_1193),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1215),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1222),
.B(n_171),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1220),
.Y(n_1263)
);

OA211x2_ASAP7_75t_L g1264 ( 
.A1(n_1228),
.A2(n_1239),
.B(n_1217),
.C(n_1235),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1217),
.B(n_174),
.Y(n_1265)
);

NAND4xp75_ASAP7_75t_L g1266 ( 
.A(n_1228),
.B(n_176),
.C(n_177),
.D(n_178),
.Y(n_1266)
);

NAND3xp33_ASAP7_75t_SL g1267 ( 
.A(n_1210),
.B(n_179),
.C(n_180),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_1239),
.B(n_181),
.C(n_182),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1226),
.A2(n_184),
.B1(n_187),
.B2(n_192),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1207),
.B(n_193),
.Y(n_1270)
);

NAND3xp33_ASAP7_75t_L g1271 ( 
.A(n_1211),
.B(n_197),
.C(n_199),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1221),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1233),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1229),
.B(n_200),
.C(n_202),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1230),
.B(n_203),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1234),
.B(n_205),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1251),
.B(n_206),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1247),
.B(n_209),
.Y(n_1278)
);

XNOR2xp5_ASAP7_75t_L g1279 ( 
.A(n_1242),
.B(n_211),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1254),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1264),
.A2(n_1235),
.B1(n_1219),
.B2(n_1213),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1254),
.B(n_1236),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1267),
.A2(n_1245),
.B1(n_1248),
.B2(n_1231),
.Y(n_1283)
);

XNOR2xp5_ASAP7_75t_L g1284 ( 
.A(n_1279),
.B(n_1243),
.Y(n_1284)
);

NOR4xp25_ASAP7_75t_L g1285 ( 
.A(n_1265),
.B(n_1212),
.C(n_1225),
.D(n_1223),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1272),
.B(n_1250),
.Y(n_1286)
);

INVx4_ASAP7_75t_L g1287 ( 
.A(n_1275),
.Y(n_1287)
);

AND2x2_ASAP7_75t_SL g1288 ( 
.A(n_1255),
.B(n_1238),
.Y(n_1288)
);

NAND4xp75_ASAP7_75t_L g1289 ( 
.A(n_1270),
.B(n_1240),
.C(n_1252),
.D(n_1249),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1272),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1259),
.Y(n_1291)
);

NAND4xp75_ASAP7_75t_L g1292 ( 
.A(n_1270),
.B(n_1241),
.C(n_1246),
.D(n_1244),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1273),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1261),
.Y(n_1294)
);

NAND4xp75_ASAP7_75t_L g1295 ( 
.A(n_1255),
.B(n_1278),
.C(n_1262),
.D(n_1263),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_L g1296 ( 
.A(n_1277),
.B(n_1227),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1253),
.Y(n_1297)
);

INVxp67_ASAP7_75t_L g1298 ( 
.A(n_1257),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1271),
.Y(n_1299)
);

BUFx3_ASAP7_75t_L g1300 ( 
.A(n_1290),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1293),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1286),
.Y(n_1302)
);

INVxp67_ASAP7_75t_L g1303 ( 
.A(n_1297),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_R g1304 ( 
.A(n_1299),
.B(n_1275),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1282),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1287),
.Y(n_1306)
);

XOR2x2_ASAP7_75t_L g1307 ( 
.A(n_1284),
.B(n_1256),
.Y(n_1307)
);

XOR2x2_ASAP7_75t_L g1308 ( 
.A(n_1295),
.B(n_1266),
.Y(n_1308)
);

XNOR2x1_ASAP7_75t_L g1309 ( 
.A(n_1289),
.B(n_1268),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1293),
.Y(n_1310)
);

XNOR2x1_ASAP7_75t_L g1311 ( 
.A(n_1307),
.B(n_1292),
.Y(n_1311)
);

AOI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1309),
.A2(n_1281),
.B1(n_1296),
.B2(n_1288),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1300),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1303),
.Y(n_1314)
);

XOR2x2_ASAP7_75t_L g1315 ( 
.A(n_1308),
.B(n_1288),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1303),
.Y(n_1316)
);

AO22x2_ASAP7_75t_SL g1317 ( 
.A1(n_1304),
.A2(n_1298),
.B1(n_1291),
.B2(n_1306),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1304),
.A2(n_1296),
.B1(n_1283),
.B2(n_1298),
.Y(n_1318)
);

AO22x2_ASAP7_75t_L g1319 ( 
.A1(n_1300),
.A2(n_1294),
.B1(n_1287),
.B2(n_1280),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1302),
.Y(n_1320)
);

INVxp33_ASAP7_75t_SL g1321 ( 
.A(n_1305),
.Y(n_1321)
);

OA22x2_ASAP7_75t_L g1322 ( 
.A1(n_1310),
.A2(n_1287),
.B1(n_1280),
.B2(n_1276),
.Y(n_1322)
);

AOI22x1_ASAP7_75t_L g1323 ( 
.A1(n_1301),
.A2(n_1285),
.B1(n_1269),
.B2(n_1274),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1319),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1314),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1319),
.Y(n_1326)
);

AOI322xp5_ASAP7_75t_L g1327 ( 
.A1(n_1312),
.A2(n_1269),
.A3(n_1258),
.B1(n_1260),
.B2(n_1301),
.C1(n_1238),
.C2(n_1237),
.Y(n_1327)
);

INVx2_ASAP7_75t_SL g1328 ( 
.A(n_1313),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1316),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1320),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1322),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1330),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1325),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1328),
.A2(n_1315),
.B1(n_1311),
.B2(n_1318),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1329),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1331),
.A2(n_1321),
.B1(n_1317),
.B2(n_1258),
.Y(n_1336)
);

NAND4xp25_ASAP7_75t_L g1337 ( 
.A(n_1327),
.B(n_1331),
.C(n_1324),
.D(n_1323),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1334),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1332),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1337),
.A2(n_1326),
.B1(n_1324),
.B2(n_1232),
.Y(n_1340)
);

AOI31xp33_ASAP7_75t_L g1341 ( 
.A1(n_1336),
.A2(n_1335),
.A3(n_1333),
.B(n_1326),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1332),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1332),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1338),
.B(n_215),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1340),
.A2(n_1237),
.B1(n_217),
.B2(n_219),
.Y(n_1345)
);

NOR2x1_ASAP7_75t_L g1346 ( 
.A(n_1341),
.B(n_216),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1342),
.Y(n_1347)
);

NOR3xp33_ASAP7_75t_L g1348 ( 
.A(n_1343),
.B(n_221),
.C(n_223),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1339),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1342),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1342),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1347),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1350),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_1346),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1345),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1351),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1344),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1349),
.Y(n_1358)
);

OAI211xp5_ASAP7_75t_L g1359 ( 
.A1(n_1354),
.A2(n_1348),
.B(n_237),
.C(n_239),
.Y(n_1359)
);

AOI22xp5_ASAP7_75t_L g1360 ( 
.A1(n_1354),
.A2(n_232),
.B1(n_241),
.B2(n_242),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1352),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1357),
.B(n_243),
.Y(n_1362)
);

OR3x2_ASAP7_75t_L g1363 ( 
.A(n_1358),
.B(n_248),
.C(n_249),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1353),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1356),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1362),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1364),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1365),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1363),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1361),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1360),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1359),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1364),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1364),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1364),
.Y(n_1375)
);

AOI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1372),
.A2(n_1355),
.B1(n_251),
.B2(n_257),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1369),
.A2(n_250),
.B1(n_262),
.B2(n_265),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1366),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1370),
.A2(n_268),
.B1(n_269),
.B2(n_272),
.Y(n_1379)
);

OAI22x1_ASAP7_75t_L g1380 ( 
.A1(n_1367),
.A2(n_275),
.B1(n_277),
.B2(n_279),
.Y(n_1380)
);

OAI22x1_ASAP7_75t_L g1381 ( 
.A1(n_1368),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1370),
.Y(n_1382)
);

HB1xp67_ASAP7_75t_L g1383 ( 
.A(n_1373),
.Y(n_1383)
);

OAI22x1_ASAP7_75t_L g1384 ( 
.A1(n_1374),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_1384)
);

AO22x2_ASAP7_75t_L g1385 ( 
.A1(n_1375),
.A2(n_289),
.B1(n_290),
.B2(n_292),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1371),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1382),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1383),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1378),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1385),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1386),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1385),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1377),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1388),
.A2(n_1376),
.B1(n_1381),
.B2(n_1380),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1389),
.A2(n_1379),
.B1(n_1384),
.B2(n_297),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1390),
.A2(n_294),
.B1(n_296),
.B2(n_298),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1396),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1394),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1398),
.A2(n_1393),
.B1(n_1391),
.B2(n_1392),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1397),
.A2(n_1395),
.B1(n_1387),
.B2(n_303),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1398),
.A2(n_301),
.B1(n_302),
.B2(n_309),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1399),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1400),
.Y(n_1403)
);

AOI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1402),
.A2(n_1401),
.B1(n_310),
.B2(n_312),
.C(n_315),
.Y(n_1404)
);

AOI211xp5_ASAP7_75t_L g1405 ( 
.A1(n_1404),
.A2(n_1403),
.B(n_318),
.C(n_320),
.Y(n_1405)
);


endmodule