module fake_netlist_6_4394_n_1714 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1714);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1714;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_44),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_36),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_57),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_18),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_35),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_23),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_98),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_76),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_27),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_32),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_100),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_12),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_47),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_43),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_12),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_109),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_93),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_22),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_133),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_73),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_49),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_77),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_34),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_1),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_54),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_38),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_58),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_68),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_143),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_151),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_36),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_7),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_14),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_55),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_43),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_137),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_92),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_28),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_146),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_95),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_67),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_128),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_41),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_56),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_114),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_69),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_33),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_70),
.Y(n_233)
);

INVx5_ASAP7_75t_SL g234 ( 
.A(n_18),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_86),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_55),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_121),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_103),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_125),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_50),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_30),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_89),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_118),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_80),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_64),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_78),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_2),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_96),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_15),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_135),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_16),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_0),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_15),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_123),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_31),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_11),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_99),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_50),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_152),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_58),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_14),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_38),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_163),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_162),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_91),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_134),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_66),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_40),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_1),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_65),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_57),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_124),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_7),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_37),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_31),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_44),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_37),
.Y(n_280)
);

BUFx2_ASAP7_75t_SL g281 ( 
.A(n_85),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_9),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_52),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_149),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_108),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_136),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_25),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_147),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_122),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_75),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_19),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_60),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_156),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_111),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_117),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_141),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_25),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_13),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_54),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_46),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_48),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_48),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_160),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_61),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_27),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_34),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_17),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_84),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_105),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_11),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_154),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_106),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_97),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_127),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_10),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_120),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_81),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_8),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_9),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_10),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_79),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_23),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_307),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_204),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_170),
.B(n_2),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_165),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_173),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_204),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_167),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_204),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_212),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_170),
.B(n_3),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_293),
.B(n_3),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_172),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_173),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_178),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_215),
.B(n_166),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_181),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_182),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_185),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_191),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_174),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_261),
.B(n_4),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_246),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_192),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_195),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_196),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_172),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_219),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_219),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_239),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_215),
.B(n_166),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_242),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_197),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_198),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_246),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_210),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_222),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_323),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_323),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_168),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_319),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_244),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_224),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_226),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_168),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_179),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_179),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_230),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_175),
.B(n_4),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_186),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_175),
.B(n_6),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_186),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_176),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_189),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_252),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_174),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_267),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_193),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_189),
.B(n_6),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_203),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_180),
.B(n_8),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_180),
.B(n_13),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_231),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_203),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_206),
.B(n_16),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_233),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_235),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_237),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_206),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_214),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_214),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_229),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_240),
.Y(n_402)
);

BUFx6f_ASAP7_75t_SL g403 ( 
.A(n_171),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_229),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_236),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_236),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_253),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_335),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_369),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_331),
.B(n_243),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_331),
.B(n_243),
.Y(n_412)
);

BUFx8_ASAP7_75t_L g413 ( 
.A(n_403),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_330),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_385),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_333),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_339),
.B(n_269),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_R g419 ( 
.A(n_341),
.B(n_292),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_343),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_339),
.B(n_269),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_374),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_387),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_376),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_R g427 ( 
.A(n_344),
.B(n_247),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_328),
.Y(n_428)
);

OR2x6_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_281),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_261),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_345),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_346),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_328),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_342),
.B(n_275),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_356),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_350),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_328),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_379),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_351),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_332),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_379),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_381),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_383),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_352),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_348),
.B(n_169),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_332),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_337),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_332),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_357),
.B(n_275),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_337),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_334),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

BUFx8_ASAP7_75t_L g457 ( 
.A(n_403),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_393),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_334),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_371),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_347),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_334),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_393),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_363),
.B(n_234),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_384),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_349),
.B(n_200),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_338),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_360),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_386),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_R g470 ( 
.A(n_358),
.B(n_329),
.Y(n_470)
);

CKINVDCx8_ASAP7_75t_R g471 ( 
.A(n_347),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_349),
.B(n_234),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_362),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_365),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_366),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_338),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_353),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_428),
.Y(n_479)
);

INVx6_ASAP7_75t_L g480 ( 
.A(n_413),
.Y(n_480)
);

INVx4_ASAP7_75t_SL g481 ( 
.A(n_447),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_431),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_372),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_435),
.B(n_373),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_441),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_452),
.B(n_296),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_409),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_414),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_452),
.B(n_296),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_450),
.B(n_454),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_447),
.B(n_169),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_447),
.B(n_377),
.Y(n_493)
);

BUFx4f_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_423),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_450),
.B(n_392),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_423),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_447),
.A2(n_380),
.B1(n_390),
.B2(n_378),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_447),
.B(n_395),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_454),
.B(n_396),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_397),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_429),
.A2(n_391),
.B1(n_388),
.B2(n_394),
.Y(n_502)
);

CKINVDCx8_ASAP7_75t_R g503 ( 
.A(n_461),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_402),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

AND2x6_ASAP7_75t_L g506 ( 
.A(n_466),
.B(n_234),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_349),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_434),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_464),
.B(n_177),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_434),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_429),
.B(n_327),
.Y(n_511)
);

AND2x6_ASAP7_75t_L g512 ( 
.A(n_466),
.B(n_234),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_461),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_427),
.B(n_193),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_414),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_419),
.Y(n_516)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_466),
.B(n_201),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_414),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_434),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_L g522 ( 
.A(n_410),
.B(n_220),
.C(n_336),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_470),
.A2(n_370),
.B1(n_403),
.B2(n_340),
.Y(n_523)
);

BUFx10_ASAP7_75t_L g524 ( 
.A(n_415),
.Y(n_524)
);

AND2x2_ASAP7_75t_SL g525 ( 
.A(n_431),
.B(n_177),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_470),
.A2(n_403),
.B1(n_382),
.B2(n_211),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_408),
.Y(n_528)
);

AND2x2_ASAP7_75t_SL g529 ( 
.A(n_431),
.B(n_245),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_429),
.B(n_412),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_429),
.B(n_398),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_434),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_451),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_429),
.B(n_399),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_425),
.Y(n_536)
);

OAI22xp33_ASAP7_75t_L g537 ( 
.A1(n_471),
.A2(n_394),
.B1(n_293),
.B2(n_284),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_426),
.B(n_399),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_451),
.B(n_200),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_418),
.B(n_404),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_426),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_451),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_428),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_451),
.B(n_251),
.Y(n_545)
);

AND3x2_ASAP7_75t_L g546 ( 
.A(n_416),
.B(n_223),
.C(n_253),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_430),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_436),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_430),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_439),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_416),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_459),
.B(n_262),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_460),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_439),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_428),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_417),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_459),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_459),
.B(n_266),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_459),
.B(n_268),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_438),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_442),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_419),
.B(n_245),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_442),
.Y(n_565)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_459),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_443),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_459),
.B(n_213),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_438),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_413),
.B(n_290),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_441),
.B(n_270),
.Y(n_574)
);

AND2x6_ASAP7_75t_L g575 ( 
.A(n_448),
.B(n_213),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_445),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_441),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_441),
.B(n_285),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_421),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_413),
.B(n_290),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_462),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_449),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_462),
.B(n_287),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_462),
.B(n_295),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_420),
.B(n_400),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_453),
.A2(n_263),
.B1(n_264),
.B2(n_322),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_413),
.A2(n_308),
.B1(n_311),
.B2(n_183),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

OAI21xp33_ASAP7_75t_SL g591 ( 
.A1(n_453),
.A2(n_225),
.B(n_221),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_411),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_456),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_456),
.A2(n_314),
.B1(n_302),
.B2(n_305),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_457),
.B(n_291),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_411),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_465),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_458),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_448),
.B(n_297),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_422),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_458),
.B(n_400),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_457),
.B(n_291),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_448),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_455),
.B(n_463),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_432),
.B(n_401),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_463),
.Y(n_606)
);

INVx5_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_476),
.B(n_401),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_422),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_476),
.Y(n_610)
);

INVxp33_ASAP7_75t_L g611 ( 
.A(n_427),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_478),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_455),
.B(n_221),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_433),
.B(n_405),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_422),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_437),
.B(n_405),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_440),
.B(n_407),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_455),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_457),
.B(n_193),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_477),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_480),
.B(n_281),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_531),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_525),
.A2(n_288),
.B1(n_298),
.B2(n_286),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_486),
.B(n_468),
.C(n_446),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_525),
.B(n_473),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_558),
.B(n_471),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_527),
.B(n_474),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_529),
.B(n_475),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_593),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_486),
.B(n_490),
.C(n_502),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_593),
.Y(n_631)
);

NOR2xp67_ASAP7_75t_L g632 ( 
.A(n_552),
.B(n_580),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_529),
.A2(n_249),
.B1(n_325),
.B2(n_318),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_504),
.B(n_477),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_531),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_504),
.B(n_485),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_535),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_485),
.B(n_477),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_502),
.B(n_204),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_524),
.B(n_471),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_494),
.B(n_193),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_480),
.B(n_225),
.Y(n_642)
);

OAI221xp5_ASAP7_75t_L g643 ( 
.A1(n_498),
.A2(n_314),
.B1(n_279),
.B2(n_302),
.C(n_274),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_507),
.B(n_478),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_498),
.A2(n_286),
.B1(n_273),
.B2(n_288),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_603),
.B(n_478),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_590),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_603),
.B(n_478),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_227),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_487),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_483),
.B(n_457),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_482),
.B(n_467),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_513),
.B(n_406),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_545),
.A2(n_424),
.B(n_467),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_481),
.B(n_193),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_530),
.A2(n_312),
.B1(n_306),
.B2(n_316),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_481),
.B(n_204),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_479),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_481),
.B(n_204),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_530),
.A2(n_260),
.B1(n_257),
.B2(n_249),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_483),
.B(n_484),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_484),
.B(n_227),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_491),
.B(n_467),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_611),
.B(n_587),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_535),
.B(n_605),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_590),
.Y(n_666)
);

O2A1O1Ixp5_ASAP7_75t_L g667 ( 
.A1(n_492),
.A2(n_315),
.B(n_273),
.C(n_260),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_490),
.A2(n_298),
.B1(n_313),
.B2(n_315),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_616),
.B(n_406),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_495),
.B(n_497),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_479),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_536),
.B(n_542),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_424),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_617),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_550),
.B(n_424),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_544),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_587),
.B(n_204),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_488),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_SL g679 ( 
.A(n_573),
.B(n_190),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_511),
.A2(n_317),
.B1(n_321),
.B2(n_320),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_551),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_555),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_505),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_544),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_597),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_614),
.B(n_204),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_556),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_511),
.A2(n_283),
.B1(n_272),
.B2(n_258),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_556),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_563),
.B(n_204),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_614),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_524),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_565),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_567),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_568),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_571),
.B(n_407),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_576),
.B(n_184),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_611),
.B(n_469),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_577),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_583),
.B(n_187),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_584),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_598),
.B(n_188),
.Y(n_702)
);

AO22x1_ASAP7_75t_L g703 ( 
.A1(n_522),
.A2(n_263),
.B1(n_264),
.B2(n_274),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_606),
.B(n_194),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_493),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_539),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_492),
.A2(n_279),
.B1(n_322),
.B2(n_305),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_562),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_501),
.B(n_199),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_570),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_518),
.B(n_202),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_570),
.Y(n_712)
);

O2A1O1Ixp5_ASAP7_75t_L g713 ( 
.A1(n_509),
.A2(n_368),
.B(n_367),
.C(n_364),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_499),
.B(n_205),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_539),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_541),
.B(n_309),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_496),
.B(n_207),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_572),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_500),
.B(n_171),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_572),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_509),
.B(n_208),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_601),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_601),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_599),
.B(n_209),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_522),
.A2(n_309),
.B1(n_171),
.B2(n_259),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_608),
.Y(n_726)
);

OAI221xp5_ASAP7_75t_L g727 ( 
.A1(n_588),
.A2(n_289),
.B1(n_216),
.B2(n_217),
.C(n_218),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_480),
.B(n_353),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_SL g729 ( 
.A1(n_541),
.A2(n_368),
.B(n_367),
.C(n_364),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_612),
.B(n_232),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_608),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_588),
.B(n_354),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_489),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_515),
.B(n_171),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_620),
.B(n_238),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_519),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_564),
.A2(n_228),
.B1(n_294),
.B2(n_282),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_574),
.B(n_241),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_523),
.B(n_248),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_579),
.B(n_250),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_540),
.B(n_254),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_585),
.B(n_255),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_SL g743 ( 
.A1(n_516),
.A2(n_303),
.B1(n_265),
.B2(n_276),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_586),
.B(n_256),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_604),
.B(n_310),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_594),
.B(n_361),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_594),
.B(n_361),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_618),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_610),
.B(n_359),
.Y(n_749)
);

NOR3xp33_ASAP7_75t_L g750 ( 
.A(n_537),
.B(n_304),
.C(n_277),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_618),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_592),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_578),
.B(n_301),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_506),
.B(n_324),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_564),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_SL g756 ( 
.A(n_619),
.B(n_299),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_506),
.B(n_326),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_537),
.B(n_278),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_512),
.B(n_280),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_540),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_619),
.A2(n_573),
.B1(n_595),
.B2(n_602),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_592),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_578),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_609),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_503),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_516),
.B(n_259),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_609),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_528),
.Y(n_768)
);

NAND2xp33_ASAP7_75t_L g769 ( 
.A(n_540),
.B(n_569),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_581),
.A2(n_355),
.B1(n_354),
.B2(n_259),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_512),
.B(n_72),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_553),
.A2(n_63),
.B(n_164),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_512),
.B(n_104),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_591),
.B(n_526),
.Y(n_774)
);

NOR3x1_ASAP7_75t_L g775 ( 
.A(n_581),
.B(n_259),
.C(n_20),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_635),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_646),
.A2(n_560),
.B(n_561),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_648),
.A2(n_532),
.B(n_557),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_661),
.B(n_505),
.Y(n_779)
);

NOR3xp33_ASAP7_75t_L g780 ( 
.A(n_664),
.B(n_589),
.C(n_548),
.Y(n_780)
);

AO22x1_ASAP7_75t_L g781 ( 
.A1(n_758),
.A2(n_554),
.B1(n_569),
.B2(n_540),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_636),
.A2(n_543),
.B(n_520),
.Y(n_782)
);

NOR3xp33_ASAP7_75t_L g783 ( 
.A(n_625),
.B(n_602),
.C(n_595),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_634),
.A2(n_557),
.B(n_549),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_644),
.A2(n_755),
.B(n_638),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_705),
.B(n_520),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_658),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_630),
.A2(n_543),
.B1(n_508),
.B2(n_559),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_683),
.A2(n_549),
.B(n_517),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_683),
.A2(n_705),
.B(n_641),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_683),
.A2(n_517),
.B(n_534),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_645),
.A2(n_505),
.B1(n_508),
.B2(n_559),
.Y(n_792)
);

NOR3xp33_ASAP7_75t_L g793 ( 
.A(n_628),
.B(n_514),
.C(n_546),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_691),
.B(n_546),
.Y(n_794)
);

AOI21x1_ASAP7_75t_L g795 ( 
.A1(n_657),
.A2(n_600),
.B(n_532),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_635),
.B(n_559),
.Y(n_796)
);

AOI21x1_ASAP7_75t_L g797 ( 
.A1(n_657),
.A2(n_534),
.B(n_505),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_662),
.B(n_582),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_SL g799 ( 
.A(n_626),
.B(n_640),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_653),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_623),
.A2(n_508),
.B1(n_533),
.B2(n_559),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_633),
.A2(n_508),
.B1(n_533),
.B2(n_578),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_652),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_774),
.A2(n_613),
.B(n_575),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_663),
.B(n_582),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_643),
.A2(n_607),
.B(n_582),
.C(n_578),
.Y(n_806)
);

O2A1O1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_639),
.A2(n_575),
.B(n_613),
.C(n_540),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_663),
.B(n_669),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_669),
.B(n_533),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_683),
.A2(n_510),
.B(n_521),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_641),
.A2(n_510),
.B(n_521),
.Y(n_811)
);

AOI22xp5_ASAP7_75t_L g812 ( 
.A1(n_665),
.A2(n_569),
.B1(n_613),
.B2(n_575),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_639),
.A2(n_739),
.B(n_679),
.C(n_716),
.Y(n_813)
);

OAI21xp5_ASAP7_75t_L g814 ( 
.A1(n_774),
.A2(n_686),
.B(n_677),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_650),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_622),
.A2(n_637),
.B1(n_635),
.B2(n_665),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_653),
.B(n_674),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_635),
.Y(n_818)
);

NOR2xp67_ASAP7_75t_L g819 ( 
.A(n_624),
.B(n_607),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_674),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_760),
.Y(n_821)
);

NOR2x1_ASAP7_75t_L g822 ( 
.A(n_692),
.B(n_615),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_677),
.A2(n_575),
.B(n_613),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_670),
.A2(n_510),
.B(n_538),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_632),
.B(n_615),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_716),
.A2(n_607),
.B(n_596),
.C(n_21),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_647),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_717),
.B(n_596),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_622),
.B(n_607),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_637),
.A2(n_566),
.B1(n_538),
.B2(n_613),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_719),
.B(n_19),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_761),
.B(n_566),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_681),
.B(n_575),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_SL g835 ( 
.A(n_651),
.B(n_20),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_682),
.B(n_569),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_686),
.A2(n_569),
.B(n_566),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_760),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_685),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_672),
.A2(n_659),
.B(n_647),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_694),
.B(n_566),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_659),
.A2(n_538),
.B(n_74),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_695),
.B(n_538),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_719),
.B(n_21),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_647),
.B(n_158),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_711),
.B(n_22),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_679),
.A2(n_24),
.B(n_26),
.C(n_28),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_655),
.A2(n_82),
.B(n_153),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_666),
.A2(n_155),
.B(n_150),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_654),
.A2(n_144),
.B(n_142),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_666),
.B(n_715),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_768),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_655),
.A2(n_138),
.B(n_131),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_699),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_671),
.A2(n_116),
.B(n_102),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_666),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_673),
.A2(n_101),
.B(n_94),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_760),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_675),
.A2(n_90),
.B(n_87),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_701),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_709),
.B(n_24),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_629),
.Y(n_863)
);

OAI321xp33_ASAP7_75t_L g864 ( 
.A1(n_668),
.A2(n_26),
.A3(n_29),
.B1(n_32),
.B2(n_33),
.C(n_35),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_631),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_732),
.A2(n_747),
.B(n_746),
.C(n_660),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_676),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_649),
.A2(n_39),
.B(n_42),
.Y(n_868)
);

O2A1O1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_729),
.A2(n_39),
.B(n_42),
.C(n_45),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_738),
.B(n_46),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_715),
.A2(n_83),
.B1(n_51),
.B2(n_53),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_684),
.A2(n_49),
.B(n_51),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_740),
.B(n_53),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_742),
.B(n_56),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_714),
.B(n_62),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_684),
.A2(n_59),
.B(n_60),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_744),
.B(n_59),
.Y(n_877)
);

NOR3xp33_ASAP7_75t_L g878 ( 
.A(n_766),
.B(n_698),
.C(n_703),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_765),
.Y(n_879)
);

AO21x1_ASAP7_75t_L g880 ( 
.A1(n_649),
.A2(n_62),
.B(n_771),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_692),
.B(n_737),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_706),
.A2(n_722),
.B1(n_723),
.B2(n_726),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_773),
.A2(n_724),
.B(n_763),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_731),
.B(n_732),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_688),
.B(n_745),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_725),
.A2(n_750),
.B(n_727),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_697),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_745),
.B(n_700),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_687),
.A2(n_708),
.B(n_751),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_763),
.A2(n_764),
.B(n_752),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_702),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_696),
.B(n_735),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_721),
.A2(n_656),
.B(n_730),
.C(n_733),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_704),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_753),
.B(n_680),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_752),
.B(n_762),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_763),
.A2(n_764),
.B(n_762),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_689),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_689),
.A2(n_718),
.B(n_720),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_767),
.A2(n_736),
.B(n_754),
.Y(n_900)
);

OAI321xp33_ASAP7_75t_L g901 ( 
.A1(n_770),
.A2(n_707),
.A3(n_734),
.B1(n_753),
.B2(n_690),
.C(n_757),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_621),
.A2(n_759),
.B1(n_627),
.B2(n_728),
.Y(n_902)
);

INVx3_ASAP7_75t_SL g903 ( 
.A(n_685),
.Y(n_903)
);

INVx11_ASAP7_75t_L g904 ( 
.A(n_775),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_710),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_769),
.A2(n_678),
.B(n_751),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_756),
.A2(n_713),
.B(n_667),
.C(n_678),
.Y(n_907)
);

INVx1_ASAP7_75t_SL g908 ( 
.A(n_743),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_678),
.B(n_748),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_769),
.A2(n_710),
.B(n_712),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_712),
.A2(n_720),
.B(n_748),
.Y(n_911)
);

INVxp67_ASAP7_75t_L g912 ( 
.A(n_734),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_756),
.A2(n_749),
.B1(n_741),
.B2(n_621),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_749),
.B(n_729),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_772),
.A2(n_741),
.B(n_642),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_642),
.B(n_661),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_646),
.A2(n_648),
.B(n_634),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_661),
.B(n_635),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_646),
.A2(n_648),
.B(n_634),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_661),
.B(n_636),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_653),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_661),
.A2(n_636),
.B1(n_630),
.B2(n_645),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_646),
.A2(n_648),
.B(n_634),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_661),
.B(n_636),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_646),
.A2(n_648),
.B(n_634),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_635),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_636),
.A2(n_634),
.B(n_644),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_646),
.A2(n_648),
.B(n_634),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_661),
.B(n_636),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_L g930 ( 
.A(n_661),
.B(n_691),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_661),
.A2(n_636),
.B1(n_630),
.B2(n_645),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_661),
.B(n_636),
.Y(n_932)
);

NAND3xp33_ASAP7_75t_SL g933 ( 
.A(n_661),
.B(n_688),
.C(n_452),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_646),
.A2(n_648),
.B(n_634),
.Y(n_934)
);

BUFx12f_ASAP7_75t_L g935 ( 
.A(n_653),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_SL g936 ( 
.A(n_651),
.B(n_611),
.Y(n_936)
);

NAND2x1p5_ASAP7_75t_L g937 ( 
.A(n_635),
.B(n_622),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_661),
.B(n_636),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_653),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_661),
.A2(n_636),
.B1(n_630),
.B2(n_645),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_653),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_920),
.A2(n_924),
.B(n_932),
.C(n_929),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_817),
.B(n_800),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_853),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_815),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_800),
.B(n_939),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_938),
.B(n_930),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_917),
.A2(n_923),
.B(n_919),
.Y(n_948)
);

AOI21x1_ASAP7_75t_L g949 ( 
.A1(n_779),
.A2(n_900),
.B(n_833),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_939),
.B(n_921),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_925),
.A2(n_934),
.B(n_928),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_930),
.B(n_808),
.Y(n_952)
);

NOR2xp67_ASAP7_75t_L g953 ( 
.A(n_887),
.B(n_891),
.Y(n_953)
);

BUFx2_ASAP7_75t_L g954 ( 
.A(n_935),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_795),
.A2(n_797),
.B(n_883),
.Y(n_955)
);

AO21x2_ASAP7_75t_L g956 ( 
.A1(n_782),
.A2(n_927),
.B(n_915),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_777),
.A2(n_790),
.B(n_784),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_776),
.B(n_818),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_776),
.B(n_818),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_837),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_821),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_829),
.A2(n_814),
.B(n_798),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_803),
.B(n_894),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_829),
.A2(n_809),
.B(n_805),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_910),
.A2(n_899),
.B(n_889),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_922),
.A2(n_940),
.B(n_931),
.Y(n_966)
);

OAI21x1_ASAP7_75t_L g967 ( 
.A1(n_841),
.A2(n_906),
.B(n_897),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_890),
.A2(n_788),
.B(n_804),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_888),
.B(n_892),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_888),
.B(n_884),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_778),
.A2(n_911),
.B(n_791),
.Y(n_971)
);

NOR2xp67_ASAP7_75t_L g972 ( 
.A(n_879),
.B(n_912),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_789),
.A2(n_807),
.B(n_823),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_903),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_785),
.A2(n_918),
.B(n_801),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_821),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_866),
.B1(n_916),
.B2(n_895),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_895),
.B(n_799),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_847),
.B(n_875),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_787),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_903),
.Y(n_981)
);

BUFx2_ASAP7_75t_L g982 ( 
.A(n_941),
.Y(n_982)
);

AOI21x1_ASAP7_75t_L g983 ( 
.A1(n_914),
.A2(n_918),
.B(n_896),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_802),
.A2(n_792),
.B(n_893),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_847),
.B(n_875),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_866),
.B(n_885),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_796),
.A2(n_786),
.B(n_852),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_933),
.A2(n_885),
.B(n_845),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_840),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_855),
.B(n_861),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_826),
.B(n_862),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_870),
.A2(n_873),
.B(n_877),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_867),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_SL g994 ( 
.A(n_821),
.B(n_825),
.Y(n_994)
);

NAND2x1_ASAP7_75t_L g995 ( 
.A(n_821),
.B(n_825),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_874),
.B(n_783),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_811),
.A2(n_838),
.B(n_851),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_810),
.A2(n_824),
.B(n_849),
.Y(n_998)
);

AO21x1_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_845),
.B(n_936),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_832),
.A2(n_886),
.B(n_876),
.C(n_872),
.Y(n_1000)
);

AND2x4_ASAP7_75t_L g1001 ( 
.A(n_926),
.B(n_863),
.Y(n_1001)
);

AOI221xp5_ASAP7_75t_SL g1002 ( 
.A1(n_848),
.A2(n_882),
.B1(n_827),
.B2(n_865),
.C(n_794),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_825),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_825),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_913),
.A2(n_828),
.B1(n_857),
.B2(n_926),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_839),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_854),
.A2(n_834),
.B(n_856),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_864),
.A2(n_848),
.B(n_827),
.C(n_794),
.Y(n_1008)
);

OAI21x1_ASAP7_75t_L g1009 ( 
.A1(n_909),
.A2(n_846),
.B(n_831),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_881),
.B(n_780),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_820),
.B(n_904),
.Y(n_1011)
);

BUFx8_ASAP7_75t_SL g1012 ( 
.A(n_839),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_905),
.Y(n_1013)
);

OAI21x1_ASAP7_75t_L g1014 ( 
.A1(n_846),
.A2(n_836),
.B(n_844),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_869),
.A2(n_871),
.B(n_835),
.C(n_901),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_907),
.A2(n_806),
.B(n_898),
.Y(n_1016)
);

NAND2x1_ASAP7_75t_L g1017 ( 
.A(n_839),
.B(n_859),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_830),
.A2(n_902),
.B(n_816),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_839),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_793),
.B(n_878),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_842),
.A2(n_843),
.B(n_937),
.Y(n_1021)
);

AO21x2_ASAP7_75t_L g1022 ( 
.A1(n_880),
.A2(n_812),
.B(n_830),
.Y(n_1022)
);

OAI22x1_ASAP7_75t_L g1023 ( 
.A1(n_908),
.A2(n_822),
.B1(n_868),
.B2(n_781),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_850),
.A2(n_858),
.B(n_860),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_859),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_819),
.B(n_859),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_859),
.B(n_817),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_920),
.A2(n_661),
.B(n_929),
.C(n_924),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_930),
.A2(n_661),
.B(n_452),
.Y(n_1029)
);

AOI21x1_ASAP7_75t_L g1030 ( 
.A1(n_779),
.A2(n_900),
.B(n_833),
.Y(n_1030)
);

AO31x2_ASAP7_75t_L g1031 ( 
.A1(n_922),
.A2(n_940),
.A3(n_931),
.B(n_880),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_821),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_903),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_795),
.A2(n_797),
.B(n_910),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_903),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_903),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_917),
.A2(n_923),
.B(n_919),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_920),
.B(n_661),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_922),
.B(n_661),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_917),
.A2(n_923),
.B(n_919),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_920),
.A2(n_661),
.B(n_929),
.C(n_924),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_920),
.A2(n_661),
.B(n_929),
.C(n_924),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_787),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_814),
.A2(n_661),
.B(n_922),
.Y(n_1047)
);

OAI21x1_ASAP7_75t_L g1048 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_815),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_930),
.B(n_661),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1051)
);

INVx3_ASAP7_75t_SL g1052 ( 
.A(n_840),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_L g1053 ( 
.A(n_885),
.B(n_661),
.C(n_664),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_920),
.B(n_661),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_920),
.B(n_661),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_920),
.A2(n_661),
.B1(n_929),
.B2(n_924),
.Y(n_1057)
);

OAI21x1_ASAP7_75t_L g1058 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_920),
.B(n_661),
.Y(n_1060)
);

NOR2xp67_ASAP7_75t_L g1061 ( 
.A(n_921),
.B(n_624),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1062)
);

NOR2x1_ASAP7_75t_SL g1063 ( 
.A(n_821),
.B(n_825),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_900),
.A2(n_795),
.B(n_797),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_795),
.A2(n_797),
.B(n_910),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_920),
.B(n_661),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_920),
.B(n_661),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_787),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_920),
.B(n_661),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_821),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_922),
.B(n_661),
.Y(n_1071)
);

AOI21x1_ASAP7_75t_L g1072 ( 
.A1(n_779),
.A2(n_900),
.B(n_833),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_981),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1050),
.A2(n_1067),
.B1(n_1066),
.B2(n_1055),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_988),
.A2(n_1000),
.B(n_1029),
.C(n_1050),
.Y(n_1075)
);

BUFx10_ASAP7_75t_L g1076 ( 
.A(n_989),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_980),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_943),
.B(n_1010),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_959),
.B(n_1027),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_950),
.B(n_947),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_945),
.Y(n_1082)
);

O2A1O1Ixp5_ASAP7_75t_L g1083 ( 
.A1(n_979),
.A2(n_985),
.B(n_966),
.C(n_1071),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1060),
.B(n_1069),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_944),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_981),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_SL g1087 ( 
.A1(n_992),
.A2(n_1047),
.B(n_1016),
.C(n_1011),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_1034),
.A2(n_1065),
.B(n_1041),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_953),
.B(n_989),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_946),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1057),
.B(n_1028),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_986),
.A2(n_1053),
.B1(n_1044),
.B2(n_1045),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_1033),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_1011),
.A2(n_984),
.B(n_996),
.C(n_1020),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_959),
.B(n_1001),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_1000),
.A2(n_969),
.B(n_963),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1012),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1035),
.Y(n_1098)
);

INVx4_ASAP7_75t_L g1099 ( 
.A(n_1035),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1036),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1028),
.A2(n_1044),
.B(n_1045),
.C(n_978),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_959),
.B(n_1001),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_952),
.B(n_942),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1033),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_1036),
.Y(n_1105)
);

INVx5_ASAP7_75t_L g1106 ( 
.A(n_1012),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_942),
.B(n_970),
.Y(n_1107)
);

OAI321xp33_ASAP7_75t_L g1108 ( 
.A1(n_1040),
.A2(n_1071),
.A3(n_977),
.B1(n_978),
.B2(n_1008),
.C(n_1015),
.Y(n_1108)
);

INVx3_ASAP7_75t_L g1109 ( 
.A(n_961),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_990),
.B(n_982),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1040),
.A2(n_1008),
.B1(n_1015),
.B2(n_1049),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_991),
.B(n_960),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_1052),
.B(n_1001),
.Y(n_1113)
);

CKINVDCx16_ASAP7_75t_R g1114 ( 
.A(n_954),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_999),
.A2(n_1061),
.B1(n_1023),
.B2(n_972),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_974),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_976),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1052),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1031),
.B(n_964),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1002),
.B(n_1031),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_993),
.A2(n_1013),
.B1(n_975),
.B2(n_962),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1031),
.B(n_1046),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1031),
.B(n_1068),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_958),
.B(n_1025),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1005),
.A2(n_1026),
.B1(n_1018),
.B2(n_1022),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_958),
.B(n_1019),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_961),
.A2(n_1019),
.B1(n_976),
.B2(n_1004),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1003),
.Y(n_1128)
);

OR2x6_ASAP7_75t_SL g1129 ( 
.A(n_1063),
.B(n_994),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_983),
.B(n_1070),
.Y(n_1130)
);

BUFx2_ASAP7_75t_SL g1131 ( 
.A(n_976),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_956),
.A2(n_1022),
.B1(n_997),
.B2(n_1024),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_976),
.B(n_1004),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1006),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1004),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_994),
.A2(n_987),
.B1(n_1042),
.B2(n_1037),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_L g1137 ( 
.A(n_1004),
.B(n_1032),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_957),
.A2(n_997),
.B(n_971),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1032),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_1032),
.B(n_1017),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1032),
.B(n_995),
.Y(n_1141)
);

AO22x1_ASAP7_75t_L g1142 ( 
.A1(n_949),
.A2(n_1072),
.B1(n_1030),
.B2(n_1009),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_968),
.A2(n_973),
.B1(n_965),
.B2(n_1009),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_L g1144 ( 
.A1(n_968),
.A2(n_1014),
.B(n_973),
.Y(n_1144)
);

NOR2xp67_ASAP7_75t_L g1145 ( 
.A(n_1021),
.B(n_998),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_967),
.A2(n_1007),
.B1(n_1021),
.B2(n_957),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_971),
.A2(n_967),
.B(n_955),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_1007),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1038),
.A2(n_1051),
.B1(n_1062),
.B2(n_1059),
.Y(n_1149)
);

INVx6_ASAP7_75t_L g1150 ( 
.A(n_998),
.Y(n_1150)
);

AO21x1_ASAP7_75t_L g1151 ( 
.A1(n_1043),
.A2(n_1058),
.B(n_1062),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1043),
.B(n_1056),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_955),
.A2(n_1048),
.B(n_1051),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1064),
.A2(n_951),
.B(n_948),
.Y(n_1154)
);

BUFx2_ASAP7_75t_R g1155 ( 
.A(n_989),
.Y(n_1155)
);

BUFx2_ASAP7_75t_SL g1156 ( 
.A(n_1033),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_945),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_988),
.A2(n_661),
.B(n_1000),
.C(n_1029),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_981),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1160)
);

INVxp67_ASAP7_75t_SL g1161 ( 
.A(n_1063),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_959),
.B(n_1027),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_981),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1050),
.A2(n_1054),
.B1(n_1055),
.B2(n_1039),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_L g1166 ( 
.A(n_1053),
.B(n_661),
.C(n_452),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_945),
.Y(n_1167)
);

OA21x2_ASAP7_75t_L g1168 ( 
.A1(n_1016),
.A2(n_966),
.B(n_951),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_953),
.B(n_661),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_943),
.B(n_817),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1050),
.A2(n_1054),
.B1(n_1055),
.B2(n_1039),
.Y(n_1172)
);

CKINVDCx20_ASAP7_75t_R g1173 ( 
.A(n_1033),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_943),
.B(n_817),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_981),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_945),
.Y(n_1177)
);

AND2x2_ASAP7_75t_SL g1178 ( 
.A(n_979),
.B(n_661),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_988),
.A2(n_661),
.B1(n_933),
.B2(n_1053),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_959),
.B(n_1027),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_944),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_979),
.A2(n_661),
.B(n_933),
.C(n_985),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_979),
.A2(n_661),
.B(n_933),
.C(n_985),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_988),
.A2(n_661),
.B1(n_933),
.B2(n_1053),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_946),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_945),
.Y(n_1186)
);

BUFx2_ASAP7_75t_SL g1187 ( 
.A(n_1033),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_959),
.B(n_1027),
.Y(n_1188)
);

OR2x2_ASAP7_75t_L g1189 ( 
.A(n_950),
.B(n_800),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1039),
.B(n_1054),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1050),
.A2(n_1054),
.B1(n_1055),
.B2(n_1039),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1050),
.A2(n_1054),
.B1(n_1055),
.B2(n_1039),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_944),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1012),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_959),
.B(n_1027),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1050),
.B(n_661),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_959),
.B(n_1027),
.Y(n_1198)
);

OR2x2_ASAP7_75t_L g1199 ( 
.A(n_950),
.B(n_800),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1150),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1197),
.A2(n_1178),
.B1(n_1166),
.B2(n_1164),
.Y(n_1201)
);

INVx2_ASAP7_75t_SL g1202 ( 
.A(n_1113),
.Y(n_1202)
);

BUFx12f_ASAP7_75t_L g1203 ( 
.A(n_1118),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1077),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1150),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_1085),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1079),
.A2(n_1084),
.B1(n_1176),
.B2(n_1171),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1160),
.A2(n_1176),
.B1(n_1171),
.B2(n_1191),
.Y(n_1208)
);

OAI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1165),
.A2(n_1190),
.B1(n_1160),
.B2(n_1172),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1123),
.Y(n_1210)
);

CKINVDCx11_ASAP7_75t_R g1211 ( 
.A(n_1173),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1090),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1179),
.A2(n_1184),
.B1(n_1169),
.B2(n_1074),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1074),
.A2(n_1193),
.B1(n_1172),
.B2(n_1164),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1121),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1192),
.A2(n_1193),
.B1(n_1111),
.B2(n_1096),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1153),
.A2(n_1088),
.B(n_1146),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1120),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1192),
.A2(n_1111),
.B1(n_1115),
.B2(n_1078),
.Y(n_1219)
);

BUFx8_ASAP7_75t_L g1220 ( 
.A(n_1195),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1106),
.A2(n_1156),
.B1(n_1187),
.B2(n_1092),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1130),
.Y(n_1222)
);

INVx8_ASAP7_75t_L g1223 ( 
.A(n_1126),
.Y(n_1223)
);

INVx6_ASAP7_75t_L g1224 ( 
.A(n_1102),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_1106),
.Y(n_1225)
);

CKINVDCx6p67_ASAP7_75t_R g1226 ( 
.A(n_1106),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1185),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1086),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1092),
.A2(n_1091),
.B1(n_1103),
.B2(n_1162),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1091),
.A2(n_1196),
.B1(n_1198),
.B2(n_1162),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1149),
.A2(n_1152),
.B(n_1143),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1149),
.A2(n_1152),
.B(n_1143),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1075),
.B(n_1158),
.Y(n_1233)
);

CKINVDCx11_ASAP7_75t_R g1234 ( 
.A(n_1076),
.Y(n_1234)
);

INVx1_ASAP7_75t_SL g1235 ( 
.A(n_1181),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1093),
.Y(n_1236)
);

INVxp33_ASAP7_75t_L g1237 ( 
.A(n_1116),
.Y(n_1237)
);

HB1xp67_ASAP7_75t_L g1238 ( 
.A(n_1185),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1106),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1080),
.A2(n_1180),
.B1(n_1198),
.B2(n_1196),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1080),
.A2(n_1180),
.B1(n_1188),
.B2(n_1174),
.Y(n_1241)
);

INVx2_ASAP7_75t_SL g1242 ( 
.A(n_1100),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1081),
.B(n_1188),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1170),
.A2(n_1112),
.B1(n_1107),
.B2(n_1089),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1144),
.A2(n_1119),
.B(n_1101),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1182),
.B(n_1183),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1126),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1168),
.A2(n_1110),
.B1(n_1194),
.B2(n_1125),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1099),
.Y(n_1249)
);

INVx2_ASAP7_75t_SL g1250 ( 
.A(n_1099),
.Y(n_1250)
);

INVx2_ASAP7_75t_SL g1251 ( 
.A(n_1105),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1083),
.B(n_1124),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1189),
.A2(n_1199),
.B1(n_1186),
.B2(n_1082),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1157),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1167),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1177),
.Y(n_1256)
);

HB1xp67_ASAP7_75t_L g1257 ( 
.A(n_1073),
.Y(n_1257)
);

CKINVDCx6p67_ASAP7_75t_R g1258 ( 
.A(n_1076),
.Y(n_1258)
);

OA21x2_ASAP7_75t_L g1259 ( 
.A1(n_1136),
.A2(n_1108),
.B(n_1151),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1148),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1161),
.A2(n_1098),
.B1(n_1159),
.B2(n_1163),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1108),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1104),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1132),
.Y(n_1264)
);

AO21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1141),
.A2(n_1139),
.B(n_1129),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1105),
.A2(n_1163),
.B1(n_1175),
.B2(n_1114),
.Y(n_1266)
);

HB1xp67_ASAP7_75t_L g1267 ( 
.A(n_1134),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1175),
.A2(n_1097),
.B1(n_1195),
.B2(n_1128),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1117),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1133),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1127),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1127),
.A2(n_1141),
.B(n_1109),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1097),
.A2(n_1195),
.B1(n_1094),
.B2(n_1140),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1087),
.A2(n_1137),
.B(n_1140),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1117),
.Y(n_1275)
);

NAND2x1p5_ASAP7_75t_L g1276 ( 
.A(n_1117),
.B(n_1135),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1135),
.Y(n_1277)
);

AOI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1131),
.A2(n_1135),
.B(n_1155),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1197),
.A2(n_661),
.B1(n_1050),
.B2(n_1039),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_SL g1280 ( 
.A1(n_1197),
.A2(n_661),
.B1(n_1050),
.B2(n_885),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1075),
.B(n_1179),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1122),
.Y(n_1282)
);

BUFx8_ASAP7_75t_L g1283 ( 
.A(n_1195),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1079),
.B(n_1084),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1095),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1197),
.A2(n_661),
.B1(n_933),
.B2(n_988),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1090),
.Y(n_1287)
);

BUFx4f_ASAP7_75t_SL g1288 ( 
.A(n_1173),
.Y(n_1288)
);

INVx6_ASAP7_75t_L g1289 ( 
.A(n_1095),
.Y(n_1289)
);

INVx4_ASAP7_75t_L g1290 ( 
.A(n_1126),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1090),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1122),
.Y(n_1292)
);

NOR2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1165),
.B(n_1020),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1142),
.A2(n_1145),
.B(n_1147),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1197),
.A2(n_661),
.B1(n_1050),
.B2(n_1039),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1075),
.B(n_1179),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1122),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1153),
.A2(n_1147),
.B(n_1088),
.Y(n_1298)
);

AO21x2_ASAP7_75t_L g1299 ( 
.A1(n_1138),
.A2(n_966),
.B(n_1147),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1075),
.B(n_1179),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1090),
.Y(n_1301)
);

OA21x2_ASAP7_75t_L g1302 ( 
.A1(n_1154),
.A2(n_966),
.B(n_1138),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1122),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1090),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1142),
.A2(n_1145),
.B(n_1147),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1075),
.B(n_1179),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1260),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1231),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1260),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1284),
.B(n_1243),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1209),
.B(n_1214),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1200),
.B(n_1205),
.Y(n_1312)
);

BUFx2_ASAP7_75t_L g1313 ( 
.A(n_1252),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1207),
.B(n_1208),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1252),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1216),
.B(n_1246),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1217),
.A2(n_1232),
.B(n_1231),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1210),
.B(n_1245),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1225),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1271),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1210),
.B(n_1245),
.Y(n_1321)
);

INVx4_ASAP7_75t_L g1322 ( 
.A(n_1223),
.Y(n_1322)
);

BUFx5_ASAP7_75t_L g1323 ( 
.A(n_1215),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1271),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1225),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1245),
.B(n_1282),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1298),
.A2(n_1305),
.B(n_1294),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1292),
.B(n_1297),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1292),
.B(n_1297),
.Y(n_1329)
);

CKINVDCx6p67_ASAP7_75t_R g1330 ( 
.A(n_1226),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1223),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1303),
.B(n_1264),
.Y(n_1332)
);

OR2x2_ASAP7_75t_L g1333 ( 
.A(n_1299),
.B(n_1259),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1218),
.Y(n_1334)
);

BUFx6f_ASAP7_75t_L g1335 ( 
.A(n_1223),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1222),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1262),
.B(n_1233),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1218),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1227),
.B(n_1248),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1227),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1254),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1259),
.B(n_1233),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1259),
.B(n_1281),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1254),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1302),
.A2(n_1272),
.B(n_1205),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1255),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1287),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1255),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1256),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1256),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1223),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1204),
.Y(n_1352)
);

BUFx2_ASAP7_75t_R g1353 ( 
.A(n_1239),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1204),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1280),
.B(n_1286),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1238),
.Y(n_1356)
);

INVx3_ASAP7_75t_L g1357 ( 
.A(n_1247),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1310),
.B(n_1288),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1307),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1314),
.B(n_1336),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1355),
.A2(n_1295),
.B1(n_1279),
.B2(n_1219),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1313),
.B(n_1306),
.Y(n_1362)
);

INVxp67_ASAP7_75t_SL g1363 ( 
.A(n_1336),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1313),
.B(n_1287),
.Y(n_1364)
);

OR2x2_ASAP7_75t_L g1365 ( 
.A(n_1315),
.B(n_1304),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1315),
.B(n_1281),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1340),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1326),
.B(n_1318),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1326),
.B(n_1306),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1314),
.B(n_1262),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1326),
.B(n_1296),
.Y(n_1371)
);

INVxp67_ASAP7_75t_L g1372 ( 
.A(n_1347),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_R g1373 ( 
.A(n_1330),
.B(n_1236),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1308),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1311),
.A2(n_1201),
.B1(n_1300),
.B2(n_1296),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1307),
.B(n_1304),
.Y(n_1376)
);

OAI222xp33_ASAP7_75t_L g1377 ( 
.A1(n_1311),
.A2(n_1300),
.B1(n_1213),
.B2(n_1244),
.C1(n_1221),
.C2(n_1229),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1316),
.A2(n_1293),
.B1(n_1244),
.B2(n_1230),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1318),
.B(n_1274),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1332),
.B(n_1293),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1316),
.A2(n_1253),
.B1(n_1291),
.B2(n_1212),
.C(n_1301),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1357),
.B(n_1290),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1318),
.B(n_1274),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1332),
.B(n_1270),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1357),
.B(n_1290),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1339),
.A2(n_1202),
.B1(n_1289),
.B2(n_1285),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1308),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1309),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1357),
.B(n_1247),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1340),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1337),
.B(n_1211),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1321),
.B(n_1274),
.Y(n_1392)
);

OAI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1337),
.A2(n_1241),
.B1(n_1273),
.B2(n_1268),
.C(n_1240),
.Y(n_1393)
);

OR2x2_ASAP7_75t_L g1394 ( 
.A(n_1339),
.B(n_1267),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1335),
.A2(n_1224),
.B1(n_1285),
.B2(n_1289),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1321),
.B(n_1274),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1321),
.B(n_1265),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1342),
.B(n_1265),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1343),
.B(n_1239),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1343),
.B(n_1290),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1358),
.B(n_1237),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_1361),
.B(n_1356),
.C(n_1266),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1361),
.B(n_1356),
.C(n_1347),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1381),
.B(n_1312),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1377),
.A2(n_1261),
.B(n_1345),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1380),
.B(n_1341),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1381),
.B(n_1206),
.C(n_1257),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1380),
.B(n_1341),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1393),
.A2(n_1323),
.B1(n_1343),
.B2(n_1342),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1410)
);

NAND3xp33_ASAP7_75t_L g1411 ( 
.A(n_1375),
.B(n_1346),
.C(n_1344),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1360),
.B(n_1344),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1369),
.B(n_1342),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1360),
.B(n_1346),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1394),
.B(n_1348),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1394),
.B(n_1348),
.Y(n_1416)
);

OAI221xp5_ASAP7_75t_SL g1417 ( 
.A1(n_1378),
.A2(n_1333),
.B1(n_1235),
.B2(n_1226),
.C(n_1330),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1370),
.B(n_1350),
.C(n_1349),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1370),
.B(n_1349),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1367),
.B(n_1350),
.Y(n_1420)
);

OA211x2_ASAP7_75t_L g1421 ( 
.A1(n_1391),
.A2(n_1353),
.B(n_1330),
.C(n_1278),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1369),
.B(n_1323),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1379),
.A2(n_1317),
.B(n_1327),
.Y(n_1423)
);

OAI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1393),
.A2(n_1242),
.B1(n_1250),
.B2(n_1251),
.C(n_1249),
.Y(n_1424)
);

NAND3xp33_ASAP7_75t_L g1425 ( 
.A(n_1386),
.B(n_1352),
.C(n_1354),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1367),
.B(n_1334),
.Y(n_1426)
);

OAI221xp5_ASAP7_75t_L g1427 ( 
.A1(n_1395),
.A2(n_1242),
.B1(n_1250),
.B2(n_1251),
.C(n_1249),
.Y(n_1427)
);

NAND4xp25_ASAP7_75t_L g1428 ( 
.A(n_1384),
.B(n_1320),
.C(n_1324),
.D(n_1333),
.Y(n_1428)
);

OAI21xp33_ASAP7_75t_L g1429 ( 
.A1(n_1362),
.A2(n_1353),
.B(n_1333),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.B(n_1323),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1371),
.B(n_1323),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1368),
.B(n_1323),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1362),
.A2(n_1289),
.B1(n_1285),
.B2(n_1224),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1377),
.A2(n_1278),
.B(n_1351),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1364),
.B(n_1334),
.Y(n_1435)
);

OAI21xp33_ASAP7_75t_L g1436 ( 
.A1(n_1362),
.A2(n_1338),
.B(n_1329),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1368),
.B(n_1397),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1364),
.B(n_1338),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1368),
.B(n_1397),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1365),
.B(n_1328),
.Y(n_1440)
);

AOI21xp5_ASAP7_75t_SL g1441 ( 
.A1(n_1363),
.A2(n_1331),
.B(n_1335),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1398),
.A2(n_1351),
.B(n_1335),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1365),
.B(n_1328),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1366),
.A2(n_1285),
.B1(n_1289),
.B2(n_1224),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1397),
.B(n_1323),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1398),
.B(n_1323),
.Y(n_1446)
);

NAND3xp33_ASAP7_75t_L g1447 ( 
.A(n_1372),
.B(n_1352),
.C(n_1354),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1398),
.B(n_1323),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1366),
.B(n_1328),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1366),
.B(n_1323),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1372),
.B(n_1329),
.Y(n_1451)
);

AND2x2_ASAP7_75t_SL g1452 ( 
.A(n_1422),
.B(n_1387),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1423),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1410),
.B(n_1379),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1434),
.A2(n_1390),
.B1(n_1400),
.B2(n_1384),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1413),
.B(n_1390),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1420),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1410),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1437),
.B(n_1379),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1432),
.B(n_1374),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1423),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1423),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1412),
.B(n_1363),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1414),
.B(n_1406),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1447),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1447),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1437),
.B(n_1383),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1428),
.B(n_1383),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1415),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1428),
.B(n_1413),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1416),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1423),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1439),
.B(n_1383),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1451),
.B(n_1392),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1439),
.B(n_1392),
.Y(n_1475)
);

OR2x2_ASAP7_75t_L g1476 ( 
.A(n_1440),
.B(n_1399),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1432),
.B(n_1392),
.Y(n_1477)
);

INVxp67_ASAP7_75t_SL g1478 ( 
.A(n_1418),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1435),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1399),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1422),
.B(n_1374),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1430),
.B(n_1396),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1438),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1430),
.B(n_1374),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1446),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1426),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1431),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1418),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1403),
.A2(n_1351),
.B1(n_1335),
.B2(n_1322),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1408),
.B(n_1396),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1419),
.B(n_1396),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1436),
.B(n_1388),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1431),
.B(n_1387),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1401),
.B(n_1234),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1449),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1450),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1479),
.B(n_1403),
.Y(n_1497)
);

OAI21xp33_ASAP7_75t_L g1498 ( 
.A1(n_1478),
.A2(n_1409),
.B(n_1429),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1458),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1452),
.B(n_1446),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1470),
.B(n_1468),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_L g1502 ( 
.A(n_1494),
.B(n_1258),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1458),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1479),
.B(n_1436),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1487),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1452),
.B(n_1448),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1483),
.B(n_1450),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1470),
.B(n_1359),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1452),
.B(n_1448),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1485),
.B(n_1459),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1487),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1487),
.Y(n_1513)
);

OAI21xp33_ASAP7_75t_L g1514 ( 
.A1(n_1455),
.A2(n_1429),
.B(n_1402),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1470),
.B(n_1359),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1488),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_R g1517 ( 
.A(n_1493),
.B(n_1421),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1485),
.B(n_1445),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1488),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1489),
.A2(n_1417),
.B1(n_1402),
.B2(n_1421),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1483),
.B(n_1404),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1465),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1469),
.B(n_1376),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1459),
.B(n_1445),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1459),
.B(n_1442),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1486),
.Y(n_1526)
);

OAI211xp5_ASAP7_75t_L g1527 ( 
.A1(n_1465),
.A2(n_1405),
.B(n_1407),
.C(n_1411),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1466),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1466),
.B(n_1407),
.C(n_1455),
.Y(n_1529)
);

INVxp67_ASAP7_75t_SL g1530 ( 
.A(n_1486),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1464),
.B(n_1258),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1495),
.A2(n_1411),
.B1(n_1424),
.B2(n_1442),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1468),
.B(n_1376),
.Y(n_1533)
);

OR2x6_ASAP7_75t_L g1534 ( 
.A(n_1468),
.B(n_1441),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1463),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1525),
.B(n_1467),
.Y(n_1536)
);

AO21x1_ASAP7_75t_SL g1537 ( 
.A1(n_1514),
.A2(n_1492),
.B(n_1456),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1532),
.B(n_1469),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1529),
.B(n_1471),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1525),
.B(n_1467),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1521),
.B(n_1471),
.Y(n_1542)
);

OAI21xp33_ASAP7_75t_L g1543 ( 
.A1(n_1498),
.A2(n_1464),
.B(n_1492),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1516),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1516),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1527),
.A2(n_1425),
.B(n_1441),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1519),
.Y(n_1547)
);

INVxp67_ASAP7_75t_SL g1548 ( 
.A(n_1497),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1522),
.B(n_1457),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1501),
.B(n_1474),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1519),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1512),
.B(n_1387),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1500),
.B(n_1467),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1534),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1528),
.B(n_1474),
.Y(n_1555)
);

OR2x2_ASAP7_75t_L g1556 ( 
.A(n_1535),
.B(n_1491),
.Y(n_1556)
);

AOI21xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1520),
.A2(n_1534),
.B(n_1531),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1499),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1499),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1503),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1530),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1510),
.B(n_1473),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1523),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1526),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1500),
.B(n_1473),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1504),
.B(n_1457),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1535),
.B(n_1491),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1508),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1506),
.B(n_1473),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1508),
.Y(n_1570)
);

NOR2x1p5_ASAP7_75t_SL g1571 ( 
.A(n_1512),
.B(n_1453),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1515),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1507),
.B(n_1495),
.Y(n_1573)
);

INVxp67_ASAP7_75t_L g1574 ( 
.A(n_1515),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1533),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1510),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1533),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1505),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1548),
.B(n_1524),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1553),
.B(n_1506),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1539),
.B(n_1524),
.Y(n_1581)
);

INVx3_ASAP7_75t_SL g1582 ( 
.A(n_1554),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1572),
.B(n_1505),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1546),
.A2(n_1534),
.B1(n_1518),
.B2(n_1509),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1552),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1553),
.B(n_1509),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1565),
.B(n_1534),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1545),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1557),
.B(n_1502),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1565),
.B(n_1518),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1552),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1566),
.B(n_1496),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1547),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1551),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1543),
.B(n_1540),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1555),
.B(n_1511),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1552),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1564),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1566),
.B(n_1561),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1569),
.B(n_1511),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1558),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1559),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1574),
.A2(n_1425),
.B(n_1427),
.Y(n_1604)
);

INVx1_ASAP7_75t_SL g1605 ( 
.A(n_1554),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1542),
.B(n_1496),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1560),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1569),
.B(n_1513),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1549),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1576),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1537),
.A2(n_1335),
.B1(n_1351),
.B2(n_1513),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1555),
.B(n_1463),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1537),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1554),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1580),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1596),
.A2(n_1570),
.B1(n_1568),
.B2(n_1577),
.C(n_1575),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1613),
.A2(n_1563),
.B(n_1576),
.Y(n_1617)
);

OAI31xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1585),
.A2(n_1536),
.A3(n_1541),
.B(n_1562),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1599),
.B(n_1536),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1591),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1590),
.A2(n_1562),
.B1(n_1541),
.B2(n_1573),
.Y(n_1621)
);

AOI211xp5_ASAP7_75t_L g1622 ( 
.A1(n_1585),
.A2(n_1538),
.B(n_1550),
.C(n_1373),
.Y(n_1622)
);

NOR4xp25_ASAP7_75t_SL g1623 ( 
.A(n_1607),
.B(n_1571),
.C(n_1517),
.D(n_1578),
.Y(n_1623)
);

OAI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1599),
.A2(n_1550),
.B1(n_1538),
.B2(n_1517),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1584),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1600),
.B(n_1562),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1605),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_L g1628 ( 
.A1(n_1605),
.A2(n_1567),
.B(n_1556),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1584),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1589),
.Y(n_1630)
);

AOI21xp33_ASAP7_75t_SL g1631 ( 
.A1(n_1604),
.A2(n_1567),
.B(n_1556),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1614),
.Y(n_1632)
);

AOI221xp5_ASAP7_75t_L g1633 ( 
.A1(n_1604),
.A2(n_1462),
.B1(n_1453),
.B2(n_1461),
.C(n_1472),
.Y(n_1633)
);

AOI322xp5_ASAP7_75t_L g1634 ( 
.A1(n_1581),
.A2(n_1454),
.A3(n_1475),
.B1(n_1496),
.B2(n_1477),
.C1(n_1482),
.C2(n_1462),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1580),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1582),
.A2(n_1571),
.B(n_1461),
.C(n_1462),
.Y(n_1636)
);

AOI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1588),
.A2(n_1385),
.B1(n_1389),
.B2(n_1382),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_SL g1638 ( 
.A1(n_1588),
.A2(n_1323),
.B1(n_1263),
.B2(n_1220),
.Y(n_1638)
);

OAI322xp33_ASAP7_75t_L g1639 ( 
.A1(n_1609),
.A2(n_1607),
.A3(n_1614),
.B1(n_1579),
.B2(n_1583),
.C1(n_1602),
.C2(n_1603),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1587),
.B(n_1477),
.Y(n_1640)
);

NAND2xp33_ASAP7_75t_R g1641 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1627),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1616),
.B(n_1582),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1627),
.B(n_1591),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1624),
.A2(n_1582),
.B1(n_1609),
.B2(n_1610),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1626),
.B(n_1203),
.Y(n_1646)
);

AND2x2_ASAP7_75t_SL g1647 ( 
.A(n_1618),
.B(n_1611),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1632),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1619),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1589),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1615),
.B(n_1593),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1631),
.B(n_1203),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1583),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1622),
.A2(n_1612),
.B1(n_1606),
.B2(n_1602),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1612),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1632),
.B(n_1594),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1635),
.B(n_1594),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1620),
.B(n_1595),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1633),
.A2(n_1608),
.B1(n_1601),
.B2(n_1603),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1617),
.B(n_1621),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_SL g1661 ( 
.A(n_1645),
.B(n_1638),
.C(n_1636),
.Y(n_1661)
);

AOI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1650),
.A2(n_1637),
.B1(n_1628),
.B2(n_1625),
.Y(n_1662)
);

AOI221xp5_ASAP7_75t_L g1663 ( 
.A1(n_1642),
.A2(n_1639),
.B1(n_1630),
.B2(n_1629),
.C(n_1595),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_L g1664 ( 
.A(n_1643),
.B(n_1640),
.C(n_1592),
.Y(n_1664)
);

XOR2x2_ASAP7_75t_L g1665 ( 
.A(n_1646),
.B(n_1220),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1660),
.A2(n_1592),
.B(n_1586),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1649),
.B(n_1601),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1649),
.B(n_1608),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1653),
.Y(n_1669)
);

OAI221xp5_ASAP7_75t_L g1670 ( 
.A1(n_1641),
.A2(n_1634),
.B1(n_1597),
.B2(n_1586),
.C(n_1592),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1648),
.B(n_1597),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1647),
.A2(n_1598),
.B(n_1586),
.C(n_1453),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_SL g1673 ( 
.A(n_1653),
.B(n_1598),
.C(n_1444),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1671),
.B(n_1652),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1669),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1667),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1668),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1661),
.B(n_1644),
.Y(n_1678)
);

AOI211x1_ASAP7_75t_L g1679 ( 
.A1(n_1670),
.A2(n_1656),
.B(n_1654),
.C(n_1658),
.Y(n_1679)
);

NOR2xp67_ASAP7_75t_L g1680 ( 
.A(n_1673),
.B(n_1655),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1663),
.B(n_1657),
.C(n_1659),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1666),
.Y(n_1682)
);

OAI211xp5_ASAP7_75t_L g1683 ( 
.A1(n_1662),
.A2(n_1651),
.B(n_1598),
.C(n_1472),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1675),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1679),
.B(n_1664),
.C(n_1672),
.Y(n_1685)
);

OAI211xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1678),
.A2(n_1665),
.B(n_1263),
.C(n_1433),
.Y(n_1686)
);

AND4x1_ASAP7_75t_L g1687 ( 
.A(n_1681),
.B(n_1674),
.C(n_1682),
.D(n_1677),
.Y(n_1687)
);

OAI311xp33_ASAP7_75t_L g1688 ( 
.A1(n_1676),
.A2(n_1480),
.A3(n_1476),
.B1(n_1456),
.C1(n_1490),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1684),
.Y(n_1689)
);

NOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1685),
.B(n_1680),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_L g1691 ( 
.A(n_1686),
.B(n_1683),
.C(n_1283),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1687),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1688),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1493),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1690),
.A2(n_1472),
.B(n_1461),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1693),
.A2(n_1220),
.B1(n_1283),
.B2(n_1228),
.Y(n_1696)
);

OR5x1_ASAP7_75t_L g1697 ( 
.A(n_1691),
.B(n_1283),
.C(n_1220),
.D(n_1493),
.E(n_1477),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1694),
.B(n_1476),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1692),
.A2(n_1283),
.B1(n_1460),
.B2(n_1484),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1696),
.Y(n_1700)
);

NOR3xp33_ASAP7_75t_L g1701 ( 
.A(n_1698),
.B(n_1689),
.C(n_1322),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1699),
.A2(n_1460),
.B1(n_1484),
.B2(n_1481),
.Y(n_1702)
);

OR3x1_ASAP7_75t_L g1703 ( 
.A(n_1700),
.B(n_1697),
.C(n_1701),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1703),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1704),
.B(n_1695),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1704),
.A2(n_1702),
.B1(n_1460),
.B2(n_1484),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1705),
.Y(n_1707)
);

OAI32xp33_ASAP7_75t_L g1708 ( 
.A1(n_1706),
.A2(n_1276),
.A3(n_1269),
.B1(n_1490),
.B2(n_1480),
.Y(n_1708)
);

AOI221xp5_ASAP7_75t_L g1709 ( 
.A1(n_1707),
.A2(n_1460),
.B1(n_1484),
.B2(n_1481),
.C(n_1482),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1708),
.A2(n_1482),
.B(n_1460),
.Y(n_1710)
);

AOI21xp5_ASAP7_75t_L g1711 ( 
.A1(n_1710),
.A2(n_1484),
.B(n_1481),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1711),
.A2(n_1709),
.B1(n_1277),
.B2(n_1275),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1712),
.A2(n_1481),
.B1(n_1475),
.B2(n_1454),
.Y(n_1713)
);

AOI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1713),
.A2(n_1319),
.B(n_1325),
.C(n_1275),
.Y(n_1714)
);


endmodule