module real_aes_8532_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_666;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g184 ( .A1(n_0), .A2(n_185), .B(n_188), .C(n_192), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_1), .B(n_176), .Y(n_195) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_3), .B(n_186), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g541 ( .A1(n_4), .A2(n_149), .B(n_152), .C(n_542), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_5), .A2(n_144), .B(n_566), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_6), .A2(n_144), .B(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_7), .B(n_176), .Y(n_572) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_8), .A2(n_178), .B(n_250), .Y(n_249) );
AND2x6_ASAP7_75t_L g149 ( .A(n_9), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_10), .A2(n_149), .B(n_152), .C(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g533 ( .A(n_11), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_12), .B(n_39), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_12), .B(n_39), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_13), .B(n_191), .Y(n_544) );
INVx1_ASAP7_75t_L g170 ( .A(n_14), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_15), .B(n_186), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_16), .A2(n_187), .B(n_552), .C(n_554), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_17), .B(n_176), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_18), .B(n_164), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g151 ( .A1(n_19), .A2(n_152), .B(n_155), .C(n_163), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_20), .A2(n_190), .B(n_258), .C(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_21), .B(n_191), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g495 ( .A(n_22), .B(n_191), .Y(n_495) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_23), .Y(n_514) );
INVx1_ASAP7_75t_L g494 ( .A(n_24), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_25), .A2(n_152), .B(n_163), .C(n_253), .Y(n_252) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_26), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_27), .Y(n_540) );
INVx1_ASAP7_75t_L g508 ( .A(n_28), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_29), .A2(n_144), .B(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g147 ( .A(n_30), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_31), .A2(n_202), .B(n_203), .C(n_207), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_32), .A2(n_33), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_32), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_33), .Y(n_124) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_34), .A2(n_190), .B(n_569), .C(n_571), .Y(n_568) );
INVxp67_ASAP7_75t_L g509 ( .A(n_35), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_36), .B(n_255), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_37), .A2(n_152), .B(n_163), .C(n_493), .Y(n_492) );
CKINVDCx14_ASAP7_75t_R g567 ( .A(n_38), .Y(n_567) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_40), .A2(n_192), .B(n_531), .C(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_41), .B(n_143), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_42), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_43), .B(n_186), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_44), .B(n_144), .Y(n_251) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_45), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_46), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_47), .A2(n_202), .B(n_207), .C(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g189 ( .A(n_48), .Y(n_189) );
INVx1_ASAP7_75t_L g233 ( .A(n_49), .Y(n_233) );
INVx1_ASAP7_75t_L g580 ( .A(n_50), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_51), .B(n_144), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_52), .Y(n_172) );
CKINVDCx14_ASAP7_75t_R g529 ( .A(n_53), .Y(n_529) );
AOI22xp5_ASAP7_75t_SL g465 ( .A1(n_54), .A2(n_457), .B1(n_466), .B2(n_763), .Y(n_465) );
INVx1_ASAP7_75t_L g150 ( .A(n_55), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_56), .B(n_144), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_57), .B(n_176), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_58), .A2(n_162), .B(n_218), .C(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g169 ( .A(n_59), .Y(n_169) );
INVx1_ASAP7_75t_SL g570 ( .A(n_60), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_61), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_62), .B(n_186), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_63), .B(n_176), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_64), .B(n_187), .Y(n_268) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_65), .A2(n_105), .B1(n_113), .B2(n_768), .Y(n_104) );
INVx1_ASAP7_75t_L g517 ( .A(n_66), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g182 ( .A(n_67), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_68), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_69), .A2(n_152), .B(n_207), .C(n_216), .Y(n_215) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_70), .Y(n_242) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_72), .A2(n_144), .B(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_73), .A2(n_95), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_73), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_74), .Y(n_521) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_75), .A2(n_103), .B1(n_476), .B2(n_477), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_75), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_76), .A2(n_144), .B(n_549), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_77), .A2(n_143), .B(n_504), .Y(n_503) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_78), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_79), .A2(n_473), .B1(n_474), .B2(n_475), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_79), .Y(n_473) );
INVx1_ASAP7_75t_L g550 ( .A(n_80), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_81), .B(n_160), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_82), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_83), .A2(n_144), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g553 ( .A(n_84), .Y(n_553) );
INVx2_ASAP7_75t_L g167 ( .A(n_85), .Y(n_167) );
INVx1_ASAP7_75t_L g543 ( .A(n_86), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_87), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_88), .B(n_191), .Y(n_269) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_89), .B(n_109), .C(n_110), .Y(n_108) );
OR2x2_ASAP7_75t_L g456 ( .A(n_89), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g468 ( .A(n_89), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_90), .A2(n_152), .B(n_207), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_91), .B(n_144), .Y(n_200) );
INVx1_ASAP7_75t_L g204 ( .A(n_92), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_93), .B(n_461), .Y(n_460) );
INVxp67_ASAP7_75t_L g245 ( .A(n_94), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_95), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_96), .A2(n_472), .B1(n_478), .B2(n_479), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_96), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_97), .B(n_178), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_98), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g217 ( .A(n_99), .Y(n_217) );
INVx1_ASAP7_75t_L g264 ( .A(n_100), .Y(n_264) );
INVx2_ASAP7_75t_L g583 ( .A(n_101), .Y(n_583) );
AND2x2_ASAP7_75t_L g235 ( .A(n_102), .B(n_166), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_103), .Y(n_476) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g769 ( .A(n_106), .Y(n_769) );
OR2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x2_ASAP7_75t_L g458 ( .A(n_109), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
AO21x2_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_464), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g767 ( .A(n_118), .Y(n_767) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_454), .B(n_460), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_126), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_123), .B(n_177), .Y(n_545) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_128), .B1(n_131), .B2(n_132), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_131), .A2(n_132), .B1(n_470), .B2(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_SL g132 ( .A(n_133), .B(n_409), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_344), .Y(n_133) );
NAND4xp25_ASAP7_75t_SL g134 ( .A(n_135), .B(n_289), .C(n_313), .D(n_336), .Y(n_134) );
AOI221xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_226), .B1(n_260), .B2(n_273), .C(n_276), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_196), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_138), .A2(n_174), .B1(n_227), .B2(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_138), .B(n_197), .Y(n_347) );
AND2x2_ASAP7_75t_L g366 ( .A(n_138), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_138), .B(n_350), .Y(n_436) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_174), .Y(n_138) );
AND2x2_ASAP7_75t_L g304 ( .A(n_139), .B(n_197), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_139), .B(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g327 ( .A(n_139), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g332 ( .A(n_139), .B(n_175), .Y(n_332) );
INVx2_ASAP7_75t_L g364 ( .A(n_139), .Y(n_364) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_139), .Y(n_408) );
AND2x2_ASAP7_75t_L g425 ( .A(n_139), .B(n_302), .Y(n_425) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g343 ( .A(n_140), .B(n_302), .Y(n_343) );
AND2x4_ASAP7_75t_L g357 ( .A(n_140), .B(n_174), .Y(n_357) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_140), .Y(n_361) );
AND2x2_ASAP7_75t_L g381 ( .A(n_140), .B(n_296), .Y(n_381) );
AND2x2_ASAP7_75t_L g431 ( .A(n_140), .B(n_198), .Y(n_431) );
AND2x2_ASAP7_75t_L g441 ( .A(n_140), .B(n_175), .Y(n_441) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_171), .Y(n_140) );
AOI21xp5_ASAP7_75t_SL g141 ( .A1(n_142), .A2(n_151), .B(n_164), .Y(n_141) );
BUFx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g265 ( .A(n_145), .B(n_149), .Y(n_265) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g153 ( .A(n_147), .Y(n_153) );
INVx1_ASAP7_75t_L g259 ( .A(n_147), .Y(n_259) );
INVx1_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
INVx3_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_148), .Y(n_191) );
INVx1_ASAP7_75t_L g255 ( .A(n_148), .Y(n_255) );
BUFx3_ASAP7_75t_L g163 ( .A(n_149), .Y(n_163) );
INVx4_ASAP7_75t_SL g194 ( .A(n_149), .Y(n_194) );
INVx5_ASAP7_75t_L g183 ( .A(n_152), .Y(n_183) );
AND2x6_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
BUFx3_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_153), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_161), .Y(n_155) );
INVx2_ASAP7_75t_L g160 ( .A(n_157), .Y(n_160) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_160), .A2(n_204), .B(n_205), .C(n_206), .Y(n_203) );
O2A1O1Ixp33_ASAP7_75t_L g232 ( .A1(n_160), .A2(n_206), .B(n_233), .C(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_160), .A2(n_517), .B(n_518), .C(n_519), .Y(n_516) );
O2A1O1Ixp5_ASAP7_75t_L g542 ( .A1(n_160), .A2(n_519), .B(n_543), .C(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_161), .A2(n_186), .B(n_494), .C(n_495), .Y(n_493) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_162), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_165), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g173 ( .A(n_166), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_166), .A2(n_230), .B(n_231), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_166), .A2(n_265), .B(n_491), .C(n_492), .Y(n_490) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_166), .A2(n_527), .B(n_534), .Y(n_526) );
AND2x2_ASAP7_75t_SL g166 ( .A(n_167), .B(n_168), .Y(n_166) );
AND2x2_ASAP7_75t_L g179 ( .A(n_167), .B(n_168), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_173), .A2(n_539), .B(n_545), .Y(n_538) );
AND2x2_ASAP7_75t_L g297 ( .A(n_174), .B(n_197), .Y(n_297) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_174), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_174), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g387 ( .A(n_174), .Y(n_387) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g275 ( .A(n_175), .B(n_212), .Y(n_275) );
AND2x2_ASAP7_75t_L g302 ( .A(n_175), .B(n_213), .Y(n_302) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_180), .B(n_195), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_177), .B(n_209), .Y(n_208) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_177), .A2(n_214), .B(n_224), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_177), .B(n_225), .Y(n_224) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_177), .A2(n_263), .B(n_270), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_177), .B(n_497), .Y(n_496) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_177), .A2(n_513), .B(n_520), .Y(n_512) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_178), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_178), .A2(n_251), .B(n_252), .Y(n_250) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g272 ( .A(n_179), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_SL g181 ( .A1(n_182), .A2(n_183), .B(n_184), .C(n_194), .Y(n_181) );
INVx2_ASAP7_75t_L g202 ( .A(n_183), .Y(n_202) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_183), .A2(n_194), .B(n_242), .C(n_243), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_SL g504 ( .A1(n_183), .A2(n_194), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_SL g528 ( .A1(n_183), .A2(n_194), .B(n_529), .C(n_530), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_183), .A2(n_194), .B(n_550), .C(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_183), .A2(n_194), .B(n_567), .C(n_568), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_SL g579 ( .A1(n_183), .A2(n_194), .B(n_580), .C(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_186), .B(n_245), .Y(n_244) );
OAI22xp33_ASAP7_75t_L g507 ( .A1(n_186), .A2(n_219), .B1(n_508), .B2(n_509), .Y(n_507) );
INVx5_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_187), .B(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_190), .B(n_570), .Y(n_569) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g531 ( .A(n_191), .Y(n_531) );
INVx2_ASAP7_75t_L g519 ( .A(n_192), .Y(n_519) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_193), .Y(n_206) );
INVx1_ASAP7_75t_L g554 ( .A(n_193), .Y(n_554) );
INVx1_ASAP7_75t_L g207 ( .A(n_194), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_196), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_210), .Y(n_196) );
OR2x2_ASAP7_75t_L g328 ( .A(n_197), .B(n_211), .Y(n_328) );
AND2x2_ASAP7_75t_L g365 ( .A(n_197), .B(n_275), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_197), .B(n_296), .Y(n_376) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_197), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_197), .B(n_332), .Y(n_449) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
BUFx2_ASAP7_75t_L g274 ( .A(n_198), .Y(n_274) );
AND2x2_ASAP7_75t_L g283 ( .A(n_198), .B(n_211), .Y(n_283) );
AND2x2_ASAP7_75t_L g399 ( .A(n_198), .B(n_294), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_198), .B(n_332), .Y(n_421) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_208), .Y(n_198) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_211), .Y(n_367) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_212), .Y(n_319) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx2_ASAP7_75t_L g296 ( .A(n_213), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_223), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_220), .C(n_221), .Y(n_216) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_219), .B(n_553), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_219), .B(n_583), .Y(n_582) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g571 ( .A(n_222), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_227), .B(n_236), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_227), .B(n_309), .Y(n_428) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_228), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g280 ( .A(n_228), .B(n_281), .Y(n_280) );
INVx5_ASAP7_75t_SL g288 ( .A(n_228), .Y(n_288) );
OR2x2_ASAP7_75t_L g311 ( .A(n_228), .B(n_281), .Y(n_311) );
OR2x2_ASAP7_75t_L g321 ( .A(n_228), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g384 ( .A(n_228), .B(n_238), .Y(n_384) );
AND2x2_ASAP7_75t_SL g422 ( .A(n_228), .B(n_237), .Y(n_422) );
NOR4xp25_ASAP7_75t_L g443 ( .A(n_228), .B(n_364), .C(n_444), .D(n_445), .Y(n_443) );
AND2x2_ASAP7_75t_L g453 ( .A(n_228), .B(n_285), .Y(n_453) );
OR2x6_ASAP7_75t_L g228 ( .A(n_229), .B(n_235), .Y(n_228) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g278 ( .A(n_237), .B(n_274), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_237), .B(n_280), .Y(n_447) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_247), .Y(n_237) );
OR2x2_ASAP7_75t_L g287 ( .A(n_238), .B(n_288), .Y(n_287) );
INVx3_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_238), .B(n_262), .Y(n_306) );
INVxp67_ASAP7_75t_L g309 ( .A(n_238), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_238), .B(n_281), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_238), .B(n_248), .Y(n_375) );
AND2x2_ASAP7_75t_L g390 ( .A(n_238), .B(n_285), .Y(n_390) );
OR2x2_ASAP7_75t_L g419 ( .A(n_238), .B(n_248), .Y(n_419) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_246), .Y(n_238) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_239), .A2(n_548), .B(n_555), .Y(n_547) );
OA21x2_ASAP7_75t_L g564 ( .A1(n_239), .A2(n_565), .B(n_572), .Y(n_564) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_239), .A2(n_578), .B(n_584), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_247), .B(n_324), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_247), .B(n_288), .Y(n_427) );
OR2x2_ASAP7_75t_L g448 ( .A(n_247), .B(n_325), .Y(n_448) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g261 ( .A(n_248), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g285 ( .A(n_248), .B(n_281), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_248), .B(n_262), .Y(n_300) );
AND2x2_ASAP7_75t_L g370 ( .A(n_248), .B(n_294), .Y(n_370) );
AND2x2_ASAP7_75t_L g404 ( .A(n_248), .B(n_288), .Y(n_404) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_249), .B(n_288), .Y(n_307) );
AND2x2_ASAP7_75t_L g335 ( .A(n_249), .B(n_262), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_256), .B(n_257), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_257), .A2(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_260), .B(n_343), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_261), .A2(n_350), .B1(n_386), .B2(n_403), .C(n_405), .Y(n_402) );
INVx5_ASAP7_75t_SL g281 ( .A(n_262), .Y(n_281) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_265), .B(n_266), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_265), .A2(n_514), .B(n_515), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g539 ( .A1(n_265), .A2(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g502 ( .A(n_272), .Y(n_502) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
OAI33xp33_ASAP7_75t_L g301 ( .A1(n_274), .A2(n_302), .A3(n_303), .B1(n_305), .B2(n_308), .B3(n_312), .Y(n_301) );
OR2x2_ASAP7_75t_L g317 ( .A(n_274), .B(n_318), .Y(n_317) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_274), .A2(n_343), .A3(n_350), .B1(n_427), .B2(n_428), .C1(n_429), .C2(n_432), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_274), .B(n_302), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_SL g450 ( .A1(n_274), .A2(n_302), .B(n_451), .C(n_453), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_275), .A2(n_290), .B1(n_295), .B2(n_298), .C(n_301), .Y(n_289) );
INVx1_ASAP7_75t_L g382 ( .A(n_275), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_275), .B(n_431), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B1(n_282), .B2(n_284), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g359 ( .A(n_280), .B(n_294), .Y(n_359) );
AND2x2_ASAP7_75t_L g417 ( .A(n_280), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g325 ( .A(n_281), .B(n_288), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_281), .B(n_294), .Y(n_353) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_283), .B(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_283), .B(n_361), .Y(n_415) );
OAI321xp33_ASAP7_75t_L g434 ( .A1(n_283), .A2(n_356), .A3(n_435), .B1(n_436), .B2(n_437), .C(n_438), .Y(n_434) );
INVx1_ASAP7_75t_L g401 ( .A(n_284), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_285), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g340 ( .A(n_285), .B(n_288), .Y(n_340) );
AOI321xp33_ASAP7_75t_L g398 ( .A1(n_285), .A2(n_302), .A3(n_399), .B1(n_400), .B2(n_401), .C(n_402), .Y(n_398) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g315 ( .A(n_287), .B(n_300), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_288), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_288), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_288), .B(n_374), .Y(n_411) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g334 ( .A(n_292), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OR2x2_ASAP7_75t_L g299 ( .A(n_293), .B(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g407 ( .A(n_294), .Y(n_407) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_297), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g330 ( .A(n_302), .Y(n_330) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_304), .B(n_339), .Y(n_388) );
OR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
OR2x2_ASAP7_75t_L g352 ( .A(n_307), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_SL g397 ( .A(n_307), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_308), .A2(n_355), .B1(n_358), .B2(n_360), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx1_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g452 ( .A(n_311), .B(n_375), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B1(n_320), .B2(n_326), .C(n_329), .Y(n_313) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx2_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
INVx1_ASAP7_75t_SL g396 ( .A(n_322), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_324), .B(n_374), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_324), .A2(n_392), .B(n_394), .Y(n_391) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g437 ( .A(n_325), .B(n_419), .Y(n_437) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_SL g339 ( .A(n_328), .Y(n_339) );
AOI21xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B(n_333), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g383 ( .A(n_335), .B(n_384), .Y(n_383) );
INVxp67_ASAP7_75t_L g445 ( .A(n_335), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B(n_341), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_339), .B(n_357), .Y(n_393) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g414 ( .A(n_343), .Y(n_414) );
NAND5xp2_ASAP7_75t_L g344 ( .A(n_345), .B(n_362), .C(n_371), .D(n_391), .E(n_398), .Y(n_344) );
O2A1O1Ixp33_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_348), .B(n_351), .C(n_354), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g386 ( .A(n_350), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_358), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
OAI21xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_366), .B(n_368), .Y(n_362) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_363), .A2(n_417), .B1(n_420), .B2(n_422), .C(n_423), .Y(n_416) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AOI321xp33_ASAP7_75t_L g371 ( .A1(n_364), .A2(n_372), .A3(n_376), .B1(n_377), .B2(n_383), .C(n_385), .Y(n_371) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g442 ( .A(n_376), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_378), .B(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g394 ( .A(n_379), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
NOR2xp67_ASAP7_75t_SL g406 ( .A(n_380), .B(n_387), .Y(n_406) );
AOI321xp33_ASAP7_75t_SL g438 ( .A1(n_383), .A2(n_439), .A3(n_440), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_396), .B(n_404), .Y(n_433) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .C(n_408), .Y(n_405) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_434), .C(n_446), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g410 ( .A1(n_411), .A2(n_412), .B(n_416), .C(n_426), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_415), .Y(n_413) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_415), .A2(n_447), .B1(n_448), .B2(n_449), .C(n_450), .Y(n_446) );
INVx1_ASAP7_75t_L g435 ( .A(n_417), .Y(n_435) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g439 ( .A(n_437), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
CKINVDCx14_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g463 ( .A(n_456), .Y(n_463) );
NOR2x2_ASAP7_75t_L g765 ( .A(n_457), .B(n_468), .Y(n_765) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_460), .A2(n_465), .B(n_766), .Y(n_464) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_469), .B1(n_480), .B2(n_482), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g481 ( .A(n_468), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_470), .A2(n_471), .B1(n_483), .B2(n_484), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g479 ( .A(n_472), .Y(n_479) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OR4x2_ASAP7_75t_L g484 ( .A(n_485), .B(n_653), .C(n_700), .D(n_740), .Y(n_484) );
NAND3xp33_ASAP7_75t_SL g485 ( .A(n_486), .B(n_599), .C(n_628), .Y(n_485) );
AOI211xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_522), .B(n_556), .C(n_592), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_487), .A2(n_612), .B(n_629), .C(n_633), .Y(n_628) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_498), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g590 ( .A(n_489), .B(n_591), .Y(n_590) );
INVx3_ASAP7_75t_SL g595 ( .A(n_489), .Y(n_595) );
HB1xp67_ASAP7_75t_L g607 ( .A(n_489), .Y(n_607) );
AND2x4_ASAP7_75t_L g611 ( .A(n_489), .B(n_563), .Y(n_611) );
AND2x2_ASAP7_75t_L g622 ( .A(n_489), .B(n_512), .Y(n_622) );
OR2x2_ASAP7_75t_L g646 ( .A(n_489), .B(n_559), .Y(n_646) );
AND2x2_ASAP7_75t_L g659 ( .A(n_489), .B(n_564), .Y(n_659) );
AND2x2_ASAP7_75t_L g699 ( .A(n_489), .B(n_685), .Y(n_699) );
AND2x2_ASAP7_75t_L g706 ( .A(n_489), .B(n_669), .Y(n_706) );
AND2x2_ASAP7_75t_L g736 ( .A(n_489), .B(n_499), .Y(n_736) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_496), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_498), .B(n_663), .Y(n_675) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_511), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_499), .B(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g613 ( .A(n_499), .B(n_511), .Y(n_613) );
BUFx3_ASAP7_75t_L g621 ( .A(n_499), .Y(n_621) );
OR2x2_ASAP7_75t_L g642 ( .A(n_499), .B(n_525), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_499), .B(n_663), .Y(n_753) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B(n_510), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AO21x2_ASAP7_75t_L g559 ( .A1(n_501), .A2(n_560), .B(n_561), .Y(n_559) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g560 ( .A(n_503), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_510), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_511), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g606 ( .A(n_511), .Y(n_606) );
AND2x2_ASAP7_75t_L g669 ( .A(n_511), .B(n_564), .Y(n_669) );
AOI221xp5_ASAP7_75t_L g671 ( .A1(n_511), .A2(n_672), .B1(n_674), .B2(n_676), .C(n_677), .Y(n_671) );
AND2x2_ASAP7_75t_L g685 ( .A(n_511), .B(n_559), .Y(n_685) );
AND2x2_ASAP7_75t_L g711 ( .A(n_511), .B(n_595), .Y(n_711) );
INVx2_ASAP7_75t_SL g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g591 ( .A(n_512), .B(n_564), .Y(n_591) );
BUFx2_ASAP7_75t_L g725 ( .A(n_512), .Y(n_725) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
OAI32xp33_ASAP7_75t_L g691 ( .A1(n_523), .A2(n_652), .A3(n_666), .B1(n_692), .B2(n_693), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
AND2x2_ASAP7_75t_L g632 ( .A(n_524), .B(n_576), .Y(n_632) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g614 ( .A(n_525), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_525), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g686 ( .A(n_525), .B(n_576), .Y(n_686) );
AND2x2_ASAP7_75t_L g697 ( .A(n_525), .B(n_589), .Y(n_697) );
BUFx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g598 ( .A(n_526), .B(n_577), .Y(n_598) );
AND2x2_ASAP7_75t_L g602 ( .A(n_526), .B(n_577), .Y(n_602) );
AND2x2_ASAP7_75t_L g637 ( .A(n_526), .B(n_588), .Y(n_637) );
AND2x2_ASAP7_75t_L g644 ( .A(n_526), .B(n_546), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_526), .A2(n_595), .B(n_606), .C(n_650), .Y(n_649) );
INVx2_ASAP7_75t_L g703 ( .A(n_526), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_526), .B(n_537), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_535), .B(n_586), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_535), .B(n_602), .Y(n_692) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g597 ( .A(n_536), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_546), .Y(n_536) );
AND2x2_ASAP7_75t_L g589 ( .A(n_537), .B(n_547), .Y(n_589) );
OR2x2_ASAP7_75t_L g604 ( .A(n_537), .B(n_547), .Y(n_604) );
AND2x2_ASAP7_75t_L g627 ( .A(n_537), .B(n_588), .Y(n_627) );
INVx1_ASAP7_75t_L g631 ( .A(n_537), .Y(n_631) );
AND2x2_ASAP7_75t_L g650 ( .A(n_537), .B(n_587), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g660 ( .A1(n_537), .A2(n_615), .B1(n_661), .B2(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_537), .B(n_703), .Y(n_727) );
AND2x2_ASAP7_75t_L g742 ( .A(n_537), .B(n_602), .Y(n_742) );
INVx4_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g574 ( .A(n_538), .Y(n_574) );
AND2x2_ASAP7_75t_L g616 ( .A(n_538), .B(n_547), .Y(n_616) );
AND2x2_ASAP7_75t_L g618 ( .A(n_538), .B(n_576), .Y(n_618) );
AND3x2_ASAP7_75t_L g680 ( .A(n_538), .B(n_644), .C(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g715 ( .A(n_546), .B(n_587), .Y(n_715) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g576 ( .A(n_547), .B(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_547), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_547), .B(n_586), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g755 ( .A(n_547), .B(n_627), .C(n_703), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_573), .B1(n_585), .B2(n_590), .Y(n_556) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_559), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g667 ( .A(n_559), .Y(n_667) );
OAI31xp33_ASAP7_75t_L g683 ( .A1(n_562), .A2(n_684), .A3(n_685), .B(n_686), .Y(n_683) );
AND2x2_ASAP7_75t_L g708 ( .A(n_562), .B(n_595), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_562), .B(n_621), .Y(n_754) );
AND2x2_ASAP7_75t_L g663 ( .A(n_563), .B(n_595), .Y(n_663) );
AND2x2_ASAP7_75t_L g724 ( .A(n_563), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g594 ( .A(n_564), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g652 ( .A(n_564), .Y(n_652) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
CKINVDCx16_ASAP7_75t_R g673 ( .A(n_574), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_575), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
AOI221x1_ASAP7_75t_SL g640 ( .A1(n_576), .A2(n_641), .B1(n_643), .B2(n_645), .C(n_647), .Y(n_640) );
INVx2_ASAP7_75t_L g588 ( .A(n_577), .Y(n_588) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_577), .Y(n_682) );
INVx1_ASAP7_75t_L g670 ( .A(n_585), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_586), .B(n_603), .Y(n_695) );
INVx1_ASAP7_75t_SL g758 ( .A(n_586), .Y(n_758) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g676 ( .A(n_589), .B(n_602), .Y(n_676) );
INVx1_ASAP7_75t_L g744 ( .A(n_590), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_590), .B(n_673), .Y(n_757) );
INVx2_ASAP7_75t_SL g596 ( .A(n_591), .Y(n_596) );
AND2x2_ASAP7_75t_L g639 ( .A(n_591), .B(n_595), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_591), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_591), .B(n_666), .Y(n_693) );
AOI21xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_596), .B(n_597), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_594), .B(n_666), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_594), .B(n_621), .Y(n_762) );
OR2x2_ASAP7_75t_L g634 ( .A(n_595), .B(n_613), .Y(n_634) );
AND2x2_ASAP7_75t_L g733 ( .A(n_595), .B(n_724), .Y(n_733) );
OAI22xp5_ASAP7_75t_SL g608 ( .A1(n_596), .A2(n_609), .B1(n_614), .B2(n_617), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_596), .B(n_642), .Y(n_641) );
OR2x2_ASAP7_75t_L g656 ( .A(n_598), .B(n_604), .Y(n_656) );
INVx1_ASAP7_75t_L g720 ( .A(n_598), .Y(n_720) );
AOI311xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_605), .A3(n_607), .B(n_608), .C(n_619), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_603), .A2(n_735), .B1(n_747), .B2(n_750), .C(n_752), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_603), .B(n_758), .Y(n_760) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g657 ( .A(n_605), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g647 ( .A1(n_606), .A2(n_648), .B(n_649), .C(n_651), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_SL g716 ( .A1(n_610), .A2(n_612), .B(n_717), .C(n_718), .Y(n_716) );
INVx3_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_611), .B(n_685), .Y(n_751) );
INVx1_ASAP7_75t_SL g612 ( .A(n_613), .Y(n_612) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_614), .A2(n_634), .B1(n_635), .B2(n_638), .C(n_640), .Y(n_633) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g636 ( .A(n_616), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g719 ( .A(n_616), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_620), .A2(n_678), .B(n_679), .C(n_683), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_621), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_621), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVxp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g643 ( .A(n_627), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_631), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g745 ( .A(n_634), .Y(n_745) );
INVx1_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_637), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g672 ( .A(n_637), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g749 ( .A(n_637), .Y(n_749) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g690 ( .A(n_639), .B(n_666), .Y(n_690) );
INVx1_ASAP7_75t_SL g684 ( .A(n_646), .Y(n_684) );
INVx1_ASAP7_75t_L g661 ( .A(n_652), .Y(n_661) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_654), .B(n_671), .C(n_687), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .A3(n_658), .B1(n_660), .B2(n_664), .C1(n_668), .C2(n_670), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g707 ( .A1(n_655), .A2(n_708), .B(n_709), .C(n_716), .Y(n_707) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_658), .A2(n_679), .B1(n_710), .B2(n_712), .Y(n_709) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_666), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g705 ( .A(n_666), .B(n_706), .Y(n_705) );
AOI32xp33_ASAP7_75t_L g756 ( .A1(n_666), .A2(n_757), .A3(n_758), .B1(n_759), .B2(n_761), .Y(n_756) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g678 ( .A(n_669), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_669), .A2(n_722), .B1(n_726), .B2(n_728), .C(n_731), .Y(n_721) );
AND2x2_ASAP7_75t_L g735 ( .A(n_669), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g738 ( .A(n_673), .B(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g748 ( .A(n_673), .B(n_749), .Y(n_748) );
INVxp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g739 ( .A(n_682), .B(n_703), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B(n_691), .C(n_694), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B(n_698), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_SL g700 ( .A1(n_701), .A2(n_704), .B(n_707), .C(n_721), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_715), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g730 ( .A(n_727), .Y(n_730) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_734), .B(n_737), .Y(n_731) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI211xp5_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_743), .B(n_746), .C(n_756), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_745), .Y(n_743) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
INVx3_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
endmodule