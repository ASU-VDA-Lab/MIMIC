module fake_jpeg_10202_n_321 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_19),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_17),
.B1(n_22),
.B2(n_33),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_50),
.B1(n_62),
.B2(n_22),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_53),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_23),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_28),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_18),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_17),
.B1(n_22),
.B2(n_33),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_63),
.B(n_65),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_20),
.Y(n_65)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_88),
.CI(n_27),
.CON(n_96),
.SN(n_96)
);

XOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_85),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_69),
.B(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_90),
.B1(n_24),
.B2(n_31),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_75),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_82),
.Y(n_109)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_46),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_34),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_87),
.C(n_89),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_48),
.A2(n_26),
.B(n_20),
.C(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_34),
.Y(n_87)
);

AOI222xp33_ASAP7_75t_L g88 ( 
.A1(n_45),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.C1(n_29),
.C2(n_35),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_35),
.C(n_38),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_24),
.B1(n_31),
.B2(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_67),
.B(n_88),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_97),
.B(n_108),
.Y(n_145)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_101),
.Y(n_121)
);

NOR2xp67_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_60),
.Y(n_100)
);

AOI31xp33_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_95),
.A3(n_94),
.B(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_107),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_49),
.B1(n_35),
.B2(n_39),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_106),
.A2(n_118),
.B1(n_119),
.B2(n_76),
.Y(n_149)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_64),
.B(n_35),
.C(n_38),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_35),
.Y(n_128)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_38),
.B1(n_29),
.B2(n_25),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_64),
.B1(n_70),
.B2(n_85),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_131),
.B1(n_147),
.B2(n_95),
.Y(n_154)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_124),
.Y(n_160)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_99),
.C(n_35),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_27),
.C(n_77),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_82),
.B1(n_80),
.B2(n_71),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_71),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_149),
.B1(n_46),
.B2(n_93),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_68),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_138),
.B(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_141),
.A2(n_27),
.B(n_19),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_75),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_142),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_115),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_144),
.B(n_146),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_99),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_112),
.A2(n_49),
.B1(n_91),
.B2(n_76),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_163),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_154),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_143),
.A2(n_96),
.B1(n_106),
.B2(n_92),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_171),
.B1(n_174),
.B2(n_183),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_140),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_162),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_182),
.C(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_16),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_123),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_93),
.B1(n_103),
.B2(n_39),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_103),
.B1(n_39),
.B2(n_84),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_117),
.B1(n_110),
.B2(n_30),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_175),
.A2(n_181),
.B1(n_149),
.B2(n_120),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_36),
.B(n_47),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_148),
.Y(n_179)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_139),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_130),
.B(n_36),
.C(n_27),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_170),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_203),
.Y(n_225)
);

NAND3xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_142),
.C(n_120),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_7),
.C(n_13),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_192),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_125),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_194),
.A2(n_195),
.B(n_200),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_172),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_156),
.A2(n_134),
.B1(n_133),
.B2(n_129),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_196),
.A2(n_208),
.B1(n_166),
.B2(n_159),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_133),
.B1(n_129),
.B2(n_30),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_202),
.B1(n_191),
.B2(n_185),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_9),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_177),
.A2(n_153),
.B1(n_176),
.B2(n_165),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_148),
.C(n_36),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_161),
.B(n_36),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_168),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_148),
.B1(n_30),
.B2(n_16),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_168),
.A2(n_30),
.B1(n_16),
.B2(n_27),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_174),
.B1(n_171),
.B2(n_152),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_212),
.B(n_183),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_214),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_215),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_157),
.Y(n_216)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_231),
.B1(n_235),
.B2(n_237),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_220),
.B(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_208),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_223),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_212),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_211),
.B1(n_222),
.B2(n_213),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_195),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_230),
.A2(n_232),
.B(n_234),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_197),
.A2(n_152),
.B1(n_158),
.B2(n_182),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_194),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_186),
.A2(n_7),
.B(n_13),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_186),
.A2(n_0),
.B(n_1),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_187),
.C(n_207),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_238),
.B(n_243),
.C(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_196),
.C(n_191),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_244),
.B(n_239),
.Y(n_265)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_216),
.B(n_188),
.CI(n_204),
.CON(n_246),
.SN(n_246)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_233),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_188),
.C(n_201),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_209),
.C(n_200),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_235),
.C(n_236),
.Y(n_264)
);

XOR2x2_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_6),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_253),
.B(n_7),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_215),
.Y(n_259)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_248),
.A2(n_214),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_260),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_221),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_270),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_233),
.B(n_229),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_262),
.A2(n_271),
.B(n_253),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_265),
.C(n_269),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_228),
.B1(n_217),
.B2(n_2),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_266),
.A2(n_245),
.B1(n_249),
.B2(n_242),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_241),
.B(n_242),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_6),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_252),
.B(n_8),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_257),
.A2(n_5),
.B(n_12),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_9),
.Y(n_273)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_287),
.B1(n_11),
.B2(n_12),
.Y(n_297)
);

FAx1_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_246),
.CI(n_243),
.CON(n_280),
.SN(n_280)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_4),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_238),
.C(n_251),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_283),
.C(n_264),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_250),
.C(n_247),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_284),
.B(n_11),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_246),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_285),
.A2(n_273),
.B(n_269),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_267),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_290),
.C(n_293),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_266),
.B(n_268),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_295),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_3),
.B(n_4),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_292),
.A2(n_297),
.B1(n_298),
.B2(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_0),
.C(n_1),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_281),
.C(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_296),
.Y(n_300)
);

INVxp67_ASAP7_75t_SL g295 ( 
.A(n_279),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_4),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_15),
.B(n_0),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_284),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_302),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_278),
.C(n_281),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_306),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_290),
.B(n_276),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_280),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_286),
.B1(n_280),
.B2(n_274),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_307),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_312),
.A2(n_301),
.B(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_309),
.C(n_310),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_316),
.B(n_315),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_300),
.C(n_277),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_297),
.B(n_15),
.Y(n_321)
);


endmodule