module fake_jpeg_5354_n_232 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_232);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_232;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_19),
.A2(n_12),
.B(n_11),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_18),
.B1(n_27),
.B2(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_20),
.B1(n_17),
.B2(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_13),
.B(n_12),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_23),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_47),
.B(n_37),
.C(n_26),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_20),
.B1(n_17),
.B2(n_25),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_52),
.B1(n_16),
.B2(n_15),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_45),
.B1(n_14),
.B2(n_15),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_24),
.B1(n_27),
.B2(n_14),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_60),
.B(n_51),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_56),
.B(n_0),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_34),
.B1(n_29),
.B2(n_38),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_73),
.B(n_48),
.C(n_43),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_46),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_14),
.B1(n_21),
.B2(n_16),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_61),
.A2(n_67),
.B1(n_51),
.B2(n_9),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_13),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_38),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_70),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_13),
.B1(n_28),
.B2(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_45),
.A2(n_22),
.B1(n_26),
.B2(n_2),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_44),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_39),
.A2(n_22),
.B1(n_1),
.B2(n_2),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_82),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_44),
.B1(n_40),
.B2(n_48),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_72),
.B1(n_70),
.B2(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_80),
.B(n_88),
.Y(n_118)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_59),
.B1(n_49),
.B2(n_42),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_94),
.Y(n_110)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_60),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_91),
.A2(n_95),
.B(n_10),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_73),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_106),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_94),
.A2(n_69),
.B1(n_73),
.B2(n_71),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_100),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_73),
.B1(n_58),
.B2(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_42),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_107),
.A2(n_87),
.B1(n_86),
.B2(n_93),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_95),
.Y(n_130)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_114),
.B(n_76),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_59),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_R g134 ( 
.A(n_115),
.B(n_89),
.Y(n_134)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_42),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_81),
.B1(n_104),
.B2(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_91),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_130),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_128),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_78),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_80),
.B(n_84),
.C(n_96),
.D(n_81),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_115),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_112),
.B(n_101),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_103),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_82),
.A3(n_96),
.B1(n_99),
.B2(n_114),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_102),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_80),
.C(n_76),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_42),
.C(n_63),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_144),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_108),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_156),
.C(n_158),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_100),
.B1(n_111),
.B2(n_77),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_149),
.B(n_119),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_118),
.B1(n_110),
.B2(n_80),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_122),
.A2(n_118),
.B1(n_112),
.B2(n_115),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_159),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_89),
.B1(n_116),
.B2(n_49),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_127),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_137),
.A2(n_85),
.B1(n_68),
.B2(n_63),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_119),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_127),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_140),
.B(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_165),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_130),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_120),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_168),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_133),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_150),
.B(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_135),
.C(n_129),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_176),
.B(n_157),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_176),
.C(n_172),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_160),
.B1(n_159),
.B2(n_146),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_183),
.A2(n_189),
.B1(n_145),
.B2(n_161),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_170),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_184),
.Y(n_199)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_187),
.A2(n_188),
.B(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_155),
.B1(n_144),
.B2(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_194),
.B(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_161),
.B1(n_168),
.B2(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_172),
.C(n_167),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_195),
.B(n_185),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_166),
.B(n_153),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_153),
.B1(n_139),
.B2(n_121),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_177),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_121),
.B1(n_68),
.B2(n_65),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_198),
.B(n_179),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_65),
.B1(n_42),
.B2(n_3),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_200),
.A2(n_8),
.B1(n_12),
.B2(n_11),
.Y(n_205)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_181),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_203),
.B(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_204),
.B(n_190),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_200),
.B1(n_197),
.B2(n_192),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_185),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_208),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_207),
.C(n_202),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_213),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_196),
.B1(n_194),
.B2(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_215),
.B(n_216),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_219),
.C(n_0),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_216),
.A2(n_207),
.B(n_186),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_10),
.B(n_9),
.Y(n_220)
);

A2O1A1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_1),
.B(n_4),
.C(n_5),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_211),
.A2(n_213),
.A3(n_214),
.B1(n_3),
.B2(n_4),
.C1(n_0),
.C2(n_6),
.Y(n_221)
);

OAI21x1_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_1),
.B(n_5),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_223)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_223),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_225),
.C(n_226),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_228),
.A2(n_222),
.B(n_220),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_227),
.C(n_6),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_6),
.C(n_7),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_231),
.B(n_7),
.Y(n_232)
);


endmodule