module real_jpeg_21017_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_0),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_0),
.B(n_24),
.Y(n_192)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_0),
.A2(n_14),
.B(n_48),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_165),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_0),
.A2(n_79),
.B1(n_152),
.B2(n_222),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_0),
.B(n_196),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_0),
.B(n_27),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g250 ( 
.A1(n_0),
.A2(n_27),
.B(n_246),
.Y(n_250)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_2),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_161),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_161),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_161),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_63),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_63),
.Y(n_149)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_5),
.B(n_47),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_52),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_7),
.A2(n_25),
.B1(n_27),
.B2(n_52),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_8),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_8),
.A2(n_25),
.B1(n_27),
.B2(n_134),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_134),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_134),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_9),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_167),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_167),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_167),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_11),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_11),
.A2(n_31),
.B1(n_47),
.B2(n_48),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_12),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_12),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_12),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_45),
.C(n_46),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_112),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_110),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_93),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_19),
.B(n_93),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_66),
.C(n_75),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g138 ( 
.A(n_20),
.B(n_66),
.CI(n_75),
.CON(n_138),
.SN(n_138)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_21),
.A2(n_22),
.B1(n_95),
.B2(n_108),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_22),
.B(n_39),
.C(n_54),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_23),
.A2(n_28),
.B1(n_89),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_23),
.A2(n_89),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_23),
.A2(n_89),
.B1(n_133),
.B2(n_178),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_24),
.B(n_33),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_24),
.B(n_91),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_24),
.A2(n_35),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_25),
.A2(n_36),
.B1(n_164),
.B2(n_171),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_25),
.A2(n_42),
.A3(n_58),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_26),
.B(n_27),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_27),
.A2(n_57),
.B(n_59),
.C(n_60),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_27),
.B(n_57),
.Y(n_59)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g164 ( 
.A(n_30),
.B(n_165),
.CON(n_164),
.SN(n_164)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_53),
.B2(n_54),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_39),
.A2(n_40),
.B1(n_100),
.B2(n_106),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_46),
.B(n_50),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_41),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_41),
.A2(n_46),
.B1(n_85),
.B2(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_41),
.A2(n_50),
.B(n_86),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_41),
.A2(n_46),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_41),
.A2(n_46),
.B1(n_217),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_41),
.A2(n_46),
.B1(n_237),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_41),
.A2(n_70),
.B(n_253),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_43),
.B1(n_57),
.B2(n_58),
.Y(n_60)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_43),
.A2(n_49),
.B(n_165),
.C(n_213),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g247 ( 
.A(n_43),
.B(n_57),
.Y(n_247)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_46),
.A2(n_72),
.B(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_46),
.B(n_165),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_47),
.B(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_61),
.B(n_64),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_55),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_55),
.A2(n_102),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_55),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_55),
.A2(n_64),
.B(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_56),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_56),
.A2(n_60),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_56),
.A2(n_60),
.B1(n_195),
.B2(n_250),
.Y(n_249)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_60),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_60),
.A2(n_68),
.B(n_104),
.Y(n_137)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_60),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_73),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_87),
.B(n_88),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_77),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_87),
.B1(n_88),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_78),
.A2(n_84),
.B1(n_87),
.B2(n_306),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_82),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_79),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_79),
.A2(n_149),
.B1(n_152),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_79),
.A2(n_81),
.B1(n_207),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_79),
.A2(n_127),
.B(n_209),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_80),
.A2(n_128),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_80),
.A2(n_83),
.B(n_151),
.Y(n_244)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_81),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_84),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_88),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_90),
.B(n_92),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_89),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_109),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_107),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_103),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_139),
.B(n_315),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_138),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_114),
.B(n_138),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_120),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_115),
.B(n_119),
.Y(n_313)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_120),
.A2(n_121),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_131),
.C(n_136),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_122),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_123),
.B(n_129),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

OAI21x1_ASAP7_75t_SL g191 ( 
.A1(n_124),
.A2(n_152),
.B(n_173),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_138),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_309),
.B(n_314),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_297),
.B(n_308),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_198),
.B(n_276),
.C(n_296),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_183),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_143),
.B(n_183),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B1(n_168),
.B2(n_182),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_146),
.B(n_155),
.C(n_182),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_153),
.B2(n_154),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_147),
.B(n_154),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_165),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_153),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_163),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_160),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_168),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_169),
.B(n_175),
.C(n_180),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_179),
.B2(n_180),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_184),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_193),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_192),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_193),
.B(n_263),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_275),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_270),
.B(n_274),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_258),
.B(n_269),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_240),
.B(n_257),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_229),
.B(n_239),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_218),
.B(n_228),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_210),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_210),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_214),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_223),
.B(n_227),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_238),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_236),
.C(n_238),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_242),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_248),
.B1(n_255),
.B2(n_256),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_243),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_251),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_249),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_266),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_267),
.C(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_278),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_294),
.B2(n_295),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_281),
.B(n_284),
.C(n_295),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_291),
.C(n_293),
.Y(n_307)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_294),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_307),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_305),
.C(n_307),
.Y(n_310)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);


endmodule