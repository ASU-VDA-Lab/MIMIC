module fake_jpeg_23948_n_139 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_34),
.Y(n_51)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_0),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_23),
.A2(n_1),
.B(n_2),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_29),
.C(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_19),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_22),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_44),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_45),
.Y(n_61)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_33),
.A2(n_38),
.B1(n_32),
.B2(n_30),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_16),
.B1(n_40),
.B2(n_18),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_14),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_30),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_58),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_40),
.C(n_37),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_47),
.C(n_56),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B1(n_71),
.B2(n_72),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_65),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_28),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_27),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_26),
.B1(n_17),
.B2(n_24),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_40),
.B1(n_4),
.B2(n_18),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_4),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_78),
.B(n_69),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_85),
.C(n_86),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_43),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_63),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_48),
.C(n_54),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_43),
.B(n_4),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_46),
.C(n_50),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_52),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_68),
.C(n_62),
.Y(n_103)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_78),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_61),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_103),
.C(n_90),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_68),
.B1(n_73),
.B2(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_101),
.B(n_102),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_80),
.C(n_77),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_103),
.C(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_113),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_111),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_116),
.Y(n_127)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_106),
.A2(n_94),
.B(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_80),
.B(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_113),
.B(n_59),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_59),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_112),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_72),
.C(n_112),
.Y(n_126)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_126),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_74),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_128),
.B(n_125),
.C(n_99),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_116),
.B(n_52),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_131),
.A2(n_126),
.B(n_50),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NAND4xp25_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_134),
.C(n_6),
.D(n_10),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_121),
.Y(n_133)
);

AOI332xp33_ASAP7_75t_SL g136 ( 
.A1(n_133),
.A2(n_135),
.A3(n_72),
.B1(n_7),
.B2(n_8),
.B3(n_10),
.C1(n_12),
.C2(n_13),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_136),
.B(n_137),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_13),
.Y(n_139)
);


endmodule