module fake_ibex_1458_n_1091 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1091);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1091;

wire n_1084;
wire n_599;
wire n_778;
wire n_822;
wire n_1042;
wire n_507;
wire n_743;
wire n_1060;
wire n_540;
wire n_754;
wire n_395;
wire n_1011;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_1041;
wire n_688;
wire n_1090;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_1079;
wire n_1031;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_1067;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_1080;
wire n_957;
wire n_1015;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_1034;
wire n_371;
wire n_974;
wire n_1036;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_1018;
wire n_1044;
wire n_449;
wire n_547;
wire n_727;
wire n_1077;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_1045;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_1061;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_1056;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_1010;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_1029;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_243;
wire n_287;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_1051;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_1053;
wire n_343;
wire n_310;
wire n_714;
wire n_1076;
wire n_1032;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_928;
wire n_655;
wire n_333;
wire n_898;
wire n_967;
wire n_400;
wire n_306;
wire n_550;
wire n_736;
wire n_1055;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_1025;
wire n_465;
wire n_1057;
wire n_1068;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_1013;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_1024;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_1075;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_1081;
wire n_215;
wire n_279;
wire n_1037;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_1021;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_1052;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_1083;
wire n_656;
wire n_1014;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_1023;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_1001;
wire n_570;
wire n_623;
wire n_585;
wire n_1030;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_543;
wire n_580;
wire n_483;
wire n_487;
wire n_769;
wire n_1082;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_1070;
wire n_1074;
wire n_777;
wire n_1017;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_1089;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_1064;
wire n_1071;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_1012;
wire n_1028;
wire n_689;
wire n_960;
wire n_1022;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_1038;
wire n_999;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_1009;
wire n_635;
wire n_979;
wire n_844;
wire n_1066;
wire n_245;
wire n_648;
wire n_589;
wire n_229;
wire n_209;
wire n_472;
wire n_571;
wire n_783;
wire n_347;
wire n_1020;
wire n_847;
wire n_830;
wire n_1062;
wire n_1004;
wire n_473;
wire n_1027;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_1072;
wire n_263;
wire n_1069;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_1063;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_1054;
wire n_672;
wire n_1039;
wire n_722;
wire n_401;
wire n_1046;
wire n_554;
wire n_553;
wire n_1078;
wire n_1043;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_566;
wire n_484;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_516;
wire n_567;
wire n_548;
wire n_943;
wire n_1049;
wire n_1086;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_564;
wire n_444;
wire n_562;
wire n_506;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_1065;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_1026;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_1033;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_1087;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_1019;
wire n_1059;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_1073;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_288;
wire n_379;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_385;
wire n_233;
wire n_414;
wire n_342;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_1016;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_1047;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_1040;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_1085;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_1048;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_1088;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_897;
wire n_889;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_921;
wire n_912;
wire n_890;
wire n_1058;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_1035;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_855;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;
wire n_1050;

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_88),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_183),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_6),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_1),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_22),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_38),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_105),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_55),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_5),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_117),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_134),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_60),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_15),
.B(n_57),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_137),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_124),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_140),
.B(n_135),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_38),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_40),
.Y(n_217)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_120),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_89),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g223 ( 
.A(n_51),
.B(n_14),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_59),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_23),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_103),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_28),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_115),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_171),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_172),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_21),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_151),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_40),
.B(n_10),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_106),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_139),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_76),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_164),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_93),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_161),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_30),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_144),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_24),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_80),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_101),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_32),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_75),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_61),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_110),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_148),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_35),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_53),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_64),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_114),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_98),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_86),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_74),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_123),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_145),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_112),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_78),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_21),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_67),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_165),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_87),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_174),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_81),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_119),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_0),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_8),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_3),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_96),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_62),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_46),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_69),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_104),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_77),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_118),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_158),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_9),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_170),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_94),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_63),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_35),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_45),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_99),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_22),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_90),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_154),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_43),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_155),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_178),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_82),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_14),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_54),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_25),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_42),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_163),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_128),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_130),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_43),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_85),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_133),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_149),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_46),
.Y(n_311)
);

INVxp67_ASAP7_75t_SL g312 ( 
.A(n_131),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_122),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_173),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_50),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_136),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_126),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_31),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_2),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_27),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_66),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_34),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_27),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_184),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_13),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_20),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_15),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_116),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_157),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_12),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_73),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_8),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_13),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_138),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_18),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_218),
.B(n_0),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_187),
.Y(n_337)
);

OAI21x1_ASAP7_75t_L g338 ( 
.A1(n_253),
.A2(n_91),
.B(n_182),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_218),
.B(n_3),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_253),
.B(n_4),
.Y(n_340)
);

BUFx8_ASAP7_75t_L g341 ( 
.A(n_262),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_189),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_268),
.B(n_4),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_195),
.A2(n_7),
.B1(n_9),
.B2(n_11),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_189),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_191),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_259),
.Y(n_347)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_7),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

CKINVDCx8_ASAP7_75t_R g351 ( 
.A(n_188),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_217),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_272),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_273),
.B(n_11),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_217),
.Y(n_355)
);

OA21x2_ASAP7_75t_L g356 ( 
.A1(n_272),
.A2(n_97),
.B(n_181),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_294),
.Y(n_357)
);

AND2x4_ASAP7_75t_L g358 ( 
.A(n_291),
.B(n_12),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_191),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_280),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_194),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_187),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_294),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_282),
.B(n_16),
.Y(n_365)
);

OA21x2_ASAP7_75t_L g366 ( 
.A1(n_196),
.A2(n_100),
.B(n_179),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_198),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_232),
.Y(n_368)
);

AND2x4_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_17),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_195),
.A2(n_19),
.B1(n_20),
.B2(n_23),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_299),
.B(n_24),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_187),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_280),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_232),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_250),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g376 ( 
.A1(n_224),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_200),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_245),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_187),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_261),
.B(n_26),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_192),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_192),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_245),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_197),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_29),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_192),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_251),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_250),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_304),
.B(n_29),
.Y(n_389)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_201),
.A2(n_107),
.B(n_177),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_204),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_303),
.B(n_31),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_205),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_300),
.B(n_32),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_246),
.B(n_33),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_251),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_190),
.B(n_34),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_197),
.Y(n_398)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_208),
.A2(n_111),
.B(n_176),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_256),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_214),
.A2(n_266),
.B1(n_292),
.B2(n_243),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_209),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_212),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_192),
.Y(n_404)
);

BUFx8_ASAP7_75t_L g405 ( 
.A(n_199),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_220),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_289),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_256),
.B(n_39),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_222),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_197),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_199),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_199),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g413 ( 
.A(n_307),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_219),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_199),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_226),
.B(n_185),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_289),
.B(n_335),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_307),
.B(n_41),
.Y(n_418)
);

OAI21x1_ASAP7_75t_L g419 ( 
.A1(n_229),
.A2(n_113),
.B(n_166),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_230),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_236),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_238),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_193),
.B(n_41),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_203),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_210),
.B(n_42),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_219),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_239),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_224),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_214),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_429)
);

NAND2x1p5_ASAP7_75t_L g430 ( 
.A(n_237),
.B(n_121),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_240),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_242),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_213),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_213),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_248),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_249),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_252),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_216),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_254),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_255),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_258),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_234),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_260),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_213),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_340),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_L g447 ( 
.A1(n_358),
.A2(n_327),
.B1(n_333),
.B2(n_332),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_202),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_346),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_337),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_221),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_340),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_358),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_228),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_368),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_368),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_417),
.B(n_263),
.Y(n_459)
);

BUFx8_ASAP7_75t_SL g460 ( 
.A(n_428),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_416),
.A2(n_324),
.B1(n_243),
.B2(n_234),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g463 ( 
.A(n_416),
.B(n_244),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_206),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_349),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_371),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_398),
.B(n_321),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_417),
.B(n_264),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_362),
.B(n_265),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

CKINVDCx6p67_ASAP7_75t_R g473 ( 
.A(n_395),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_410),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_385),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_438),
.B(n_206),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_416),
.A2(n_315),
.B1(n_293),
.B2(n_330),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_361),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_362),
.A2(n_275),
.B1(n_286),
.B2(n_302),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_348),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_388),
.B(n_247),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_410),
.B(n_267),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_336),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_378),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_269),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_367),
.B(n_270),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_347),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_337),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_413),
.B(n_426),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_383),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_348),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_281),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_337),
.Y(n_498)
);

INVxp67_ASAP7_75t_SL g499 ( 
.A(n_336),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_395),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_426),
.B(n_284),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_337),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_414),
.B(n_207),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_367),
.A2(n_421),
.B1(n_391),
.B2(n_441),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_384),
.B(n_207),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_337),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_383),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_424),
.B(n_276),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_350),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_377),
.B(n_285),
.Y(n_510)
);

INVx6_ASAP7_75t_L g511 ( 
.A(n_405),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_SL g512 ( 
.A(n_339),
.B(n_266),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_339),
.Y(n_513)
);

BUFx2_ASAP7_75t_L g514 ( 
.A(n_341),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_353),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_341),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_369),
.A2(n_324),
.B1(n_309),
.B2(n_292),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_387),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_396),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_353),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_369),
.B(n_320),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_363),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_357),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_364),
.Y(n_525)
);

INVx4_ASAP7_75t_SL g526 ( 
.A(n_384),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_369),
.B(n_287),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_377),
.B(n_288),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_341),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_364),
.Y(n_530)
);

OR2x2_ASAP7_75t_SL g531 ( 
.A(n_397),
.B(n_325),
.Y(n_531)
);

AND2x6_ASAP7_75t_L g532 ( 
.A(n_369),
.B(n_295),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_391),
.B(n_393),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_341),
.Y(n_534)
);

NAND3x1_ASAP7_75t_L g535 ( 
.A(n_400),
.B(n_235),
.C(n_311),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_430),
.B(n_225),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_402),
.B(n_298),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_403),
.A2(n_244),
.B1(n_328),
.B2(n_313),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_365),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_403),
.B(n_329),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_406),
.B(n_331),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_392),
.A2(n_309),
.B1(n_310),
.B2(n_227),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_354),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_392),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_406),
.A2(n_244),
.B1(n_233),
.B2(n_334),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_361),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_409),
.B(n_308),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_396),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_407),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_409),
.B(n_308),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_421),
.B(n_312),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_407),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_431),
.B(n_213),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_431),
.B(n_241),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_397),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_355),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_432),
.B(n_223),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_420),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_432),
.B(n_271),
.Y(n_559)
);

INVx6_ASAP7_75t_L g560 ( 
.A(n_405),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_420),
.Y(n_561)
);

AND3x2_ASAP7_75t_L g562 ( 
.A(n_376),
.B(n_211),
.C(n_310),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_343),
.B(n_231),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_422),
.Y(n_565)
);

BUFx10_ASAP7_75t_L g566 ( 
.A(n_373),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_355),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_351),
.B(n_274),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_427),
.Y(n_569)
);

INVx4_ASAP7_75t_L g570 ( 
.A(n_356),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_363),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_427),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_461),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_461),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_380),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_543),
.B(n_547),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_514),
.B(n_401),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_516),
.B(n_344),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_470),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g582 ( 
.A1(n_462),
.A2(n_400),
.B1(n_487),
.B2(n_442),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_474),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_563),
.B(n_394),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_533),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_529),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_547),
.B(n_435),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_463),
.A2(n_455),
.B1(n_457),
.B2(n_453),
.Y(n_591)
);

AOI21xp5_ASAP7_75t_L g592 ( 
.A1(n_446),
.A2(n_356),
.B(n_390),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_464),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_463),
.A2(n_418),
.B1(n_408),
.B2(n_442),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_550),
.B(n_435),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_550),
.B(n_436),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_542),
.A2(n_344),
.B1(n_370),
.B2(n_311),
.Y(n_597)
);

BUFx12f_ASAP7_75t_SL g598 ( 
.A(n_476),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_445),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_522),
.A2(n_429),
.B1(n_376),
.B2(n_370),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_556),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_534),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_452),
.A2(n_437),
.B1(n_443),
.B2(n_440),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_465),
.B(n_436),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_558),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_559),
.B(n_439),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_478),
.A2(n_555),
.B1(n_466),
.B2(n_467),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_468),
.B(n_503),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_505),
.B(n_423),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_564),
.B(n_425),
.Y(n_612)
);

NOR2xp67_ASAP7_75t_L g613 ( 
.A(n_479),
.B(n_359),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g614 ( 
.A1(n_478),
.A2(n_277),
.B1(n_257),
.B2(n_326),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_535),
.B(n_338),
.Y(n_615)
);

OAI22x1_ASAP7_75t_L g616 ( 
.A1(n_517),
.A2(n_323),
.B1(n_290),
.B2(n_296),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_565),
.Y(n_617)
);

AND2x2_ASAP7_75t_SL g618 ( 
.A(n_448),
.B(n_451),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_567),
.Y(n_619)
);

AND2x2_ASAP7_75t_SL g620 ( 
.A(n_536),
.B(n_356),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_472),
.B(n_360),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_475),
.B(n_278),
.Y(n_622)
);

BUFx5_ASAP7_75t_L g623 ( 
.A(n_527),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_480),
.B(n_481),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_449),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_527),
.A2(n_342),
.B1(n_345),
.B2(n_352),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_504),
.B(n_360),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_570),
.A2(n_356),
.B(n_390),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_569),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_531),
.A2(n_318),
.B1(n_319),
.B2(n_322),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_456),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_527),
.A2(n_345),
.B1(n_352),
.B2(n_342),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_572),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_566),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_449),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_522),
.B(n_279),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_527),
.A2(n_366),
.B1(n_390),
.B2(n_338),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_460),
.Y(n_639)
);

OR2x6_ASAP7_75t_L g640 ( 
.A(n_494),
.B(n_399),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_468),
.B(n_297),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_515),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_544),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_513),
.B(n_283),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_447),
.B(n_539),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_500),
.A2(n_366),
.B1(n_390),
.B2(n_301),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_454),
.B(n_485),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_473),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_551),
.B(n_306),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_511),
.B(n_399),
.Y(n_650)
);

NOR2x2_ASAP7_75t_L g651 ( 
.A(n_512),
.B(n_419),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_486),
.B(n_366),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_490),
.B(n_366),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_546),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_527),
.A2(n_532),
.B1(n_530),
.B2(n_525),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_532),
.A2(n_419),
.B1(n_314),
.B2(n_316),
.Y(n_656)
);

AND2x6_ASAP7_75t_SL g657 ( 
.A(n_557),
.B(n_215),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_490),
.B(n_305),
.Y(n_658)
);

O2A1O1Ixp5_ASAP7_75t_L g659 ( 
.A1(n_570),
.A2(n_305),
.B(n_314),
.C(n_316),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_521),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_532),
.A2(n_305),
.B1(n_314),
.B2(n_316),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_497),
.B(n_305),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_477),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_SL g664 ( 
.A(n_508),
.B(n_314),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_497),
.B(n_316),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_501),
.A2(n_444),
.B(n_434),
.C(n_433),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_492),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_L g668 ( 
.A1(n_532),
.A2(n_444),
.B1(n_434),
.B2(n_433),
.Y(n_668)
);

O2A1O1Ixp5_ASAP7_75t_L g669 ( 
.A1(n_528),
.A2(n_444),
.B(n_434),
.C(n_433),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_501),
.B(n_404),
.Y(n_670)
);

AND2x6_ASAP7_75t_SL g671 ( 
.A(n_557),
.B(n_444),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_532),
.A2(n_444),
.B1(n_434),
.B2(n_433),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_568),
.A2(n_434),
.B1(n_433),
.B2(n_415),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_545),
.A2(n_415),
.B1(n_412),
.B2(n_411),
.Y(n_674)
);

AND3x1_ASAP7_75t_L g675 ( 
.A(n_482),
.B(n_56),
.C(n_58),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_566),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_654),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_588),
.B(n_459),
.Y(n_678)
);

O2A1O1Ixp33_ASAP7_75t_L g679 ( 
.A1(n_582),
.A2(n_469),
.B(n_528),
.C(n_471),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_634),
.Y(n_680)
);

AO21x2_ASAP7_75t_L g681 ( 
.A1(n_628),
.A2(n_537),
.B(n_491),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_604),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_R g683 ( 
.A(n_639),
.B(n_539),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_578),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_579),
.B(n_648),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_676),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_577),
.B(n_471),
.Y(n_687)
);

NOR2xp67_ASAP7_75t_SL g688 ( 
.A(n_589),
.B(n_511),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_587),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_643),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_635),
.B(n_554),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_625),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_625),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_642),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_573),
.Y(n_695)
);

XNOR2xp5_ASAP7_75t_L g696 ( 
.A(n_582),
.B(n_562),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_642),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_647),
.B(n_482),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_573),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_577),
.B(n_526),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_602),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_653),
.A2(n_592),
.B(n_576),
.Y(n_702)
);

BUFx12f_ASAP7_75t_L g703 ( 
.A(n_580),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_575),
.B(n_612),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_608),
.A2(n_510),
.B1(n_541),
.B2(n_540),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_587),
.Y(n_706)
);

A2O1A1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_610),
.A2(n_510),
.B(n_537),
.C(n_541),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_599),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_590),
.B(n_540),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_579),
.B(n_560),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_620),
.A2(n_552),
.B(n_548),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_579),
.A2(n_560),
.B1(n_524),
.B2(n_509),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_605),
.Y(n_713)
);

O2A1O1Ixp33_ASAP7_75t_L g714 ( 
.A1(n_645),
.A2(n_518),
.B(n_484),
.C(n_549),
.Y(n_714)
);

INVx3_ASAP7_75t_L g715 ( 
.A(n_660),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_607),
.A2(n_483),
.B(n_496),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_599),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_660),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_671),
.Y(n_719)
);

CKINVDCx8_ASAP7_75t_R g720 ( 
.A(n_657),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_621),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_593),
.B(n_560),
.Y(n_722)
);

OAI22xp5_ASAP7_75t_L g723 ( 
.A1(n_591),
.A2(n_545),
.B1(n_538),
.B2(n_488),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_605),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_591),
.A2(n_655),
.B1(n_626),
.B2(n_632),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_659),
.A2(n_519),
.B(n_495),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_624),
.A2(n_520),
.B(n_507),
.C(n_489),
.Y(n_727)
);

OR2x6_ASAP7_75t_L g728 ( 
.A(n_580),
.B(n_496),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_594),
.B(n_622),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_574),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_623),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_610),
.B(n_553),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_627),
.A2(n_553),
.B(n_65),
.C(n_68),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_623),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_623),
.B(n_571),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_580),
.B(n_616),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_615),
.A2(n_553),
.B1(n_412),
.B2(n_411),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_646),
.A2(n_450),
.B(n_523),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_606),
.Y(n_739)
);

O2A1O1Ixp33_ASAP7_75t_L g740 ( 
.A1(n_630),
.A2(n_553),
.B(n_71),
.C(n_72),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_581),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_611),
.A2(n_411),
.B(n_372),
.C(n_379),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_595),
.B(n_382),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_596),
.B(n_382),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_618),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_586),
.A2(n_523),
.B(n_506),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_615),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_655),
.B(n_571),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_650),
.A2(n_506),
.B(n_502),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_626),
.B(n_404),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_609),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_615),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_659),
.A2(n_502),
.B(n_498),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_632),
.A2(n_404),
.B1(n_372),
.B2(n_379),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_603),
.B(n_412),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_600),
.B(n_411),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_583),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_600),
.B(n_404),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_618),
.B(n_386),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_603),
.B(n_404),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_SL g761 ( 
.A1(n_597),
.A2(n_386),
.B1(n_382),
.B2(n_381),
.Y(n_761)
);

NOR2x1_ASAP7_75t_L g762 ( 
.A(n_637),
.B(n_382),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_650),
.A2(n_498),
.B(n_493),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_617),
.Y(n_764)
);

BUFx4f_ASAP7_75t_L g765 ( 
.A(n_584),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_670),
.A2(n_493),
.B(n_450),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_656),
.A2(n_381),
.B1(n_372),
.B2(n_386),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_649),
.B(n_381),
.Y(n_768)
);

O2A1O1Ixp5_ASAP7_75t_L g769 ( 
.A1(n_664),
.A2(n_493),
.B(n_450),
.C(n_95),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_601),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_658),
.A2(n_386),
.B(n_382),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_613),
.A2(n_386),
.B1(n_381),
.B2(n_379),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_629),
.B(n_379),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_614),
.A2(n_83),
.B(n_92),
.C(n_102),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_638),
.A2(n_363),
.B(n_372),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_644),
.B(n_363),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_633),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_675),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_641),
.B(n_125),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_682),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_738),
.A2(n_666),
.A3(n_662),
.B(n_665),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_696),
.A2(n_692),
.B1(n_698),
.B2(n_704),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_775),
.A2(n_638),
.B(n_669),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_775),
.A2(n_669),
.B(n_656),
.Y(n_784)
);

INVxp33_ASAP7_75t_L g785 ( 
.A(n_683),
.Y(n_785)
);

O2A1O1Ixp5_ASAP7_75t_L g786 ( 
.A1(n_759),
.A2(n_779),
.B(n_702),
.C(n_763),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_677),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_SL g788 ( 
.A1(n_685),
.A2(n_640),
.B1(n_585),
.B2(n_651),
.Y(n_788)
);

OA21x2_ASAP7_75t_L g789 ( 
.A1(n_753),
.A2(n_661),
.B(n_673),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_684),
.Y(n_790)
);

OAI21xp5_ASAP7_75t_L g791 ( 
.A1(n_711),
.A2(n_667),
.B(n_674),
.Y(n_791)
);

AO32x2_ASAP7_75t_L g792 ( 
.A1(n_761),
.A2(n_705),
.A3(n_725),
.B1(n_767),
.B2(n_754),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_739),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_679),
.A2(n_619),
.B(n_601),
.C(n_636),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_751),
.Y(n_795)
);

AO31x2_ASAP7_75t_L g796 ( 
.A1(n_767),
.A2(n_663),
.A3(n_631),
.B(n_668),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_749),
.A2(n_672),
.B(n_668),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_705),
.A2(n_127),
.B(n_129),
.C(n_132),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_690),
.B(n_162),
.Y(n_799)
);

INVx1_ASAP7_75t_SL g800 ( 
.A(n_701),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_694),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_764),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_686),
.Y(n_803)
);

A2O1A1Ixp33_ASAP7_75t_L g804 ( 
.A1(n_729),
.A2(n_141),
.B(n_143),
.C(n_146),
.Y(n_804)
);

HB1xp67_ASAP7_75t_L g805 ( 
.A(n_693),
.Y(n_805)
);

BUFx4f_ASAP7_75t_SL g806 ( 
.A(n_680),
.Y(n_806)
);

OAI222xp33_ASAP7_75t_L g807 ( 
.A1(n_685),
.A2(n_728),
.B1(n_778),
.B2(n_736),
.C1(n_719),
.C2(n_720),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_687),
.B(n_715),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_732),
.A2(n_150),
.B(n_153),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_777),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_743),
.A2(n_744),
.B(n_687),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_774),
.B(n_160),
.C(n_772),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_744),
.A2(n_681),
.B(n_768),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_681),
.A2(n_716),
.B(n_746),
.Y(n_814)
);

AO31x2_ASAP7_75t_L g815 ( 
.A1(n_742),
.A2(n_755),
.A3(n_760),
.B(n_754),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_688),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_713),
.A2(n_745),
.B1(n_685),
.B2(n_725),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_721),
.B(n_728),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_703),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_724),
.Y(n_820)
);

O2A1O1Ixp33_ASAP7_75t_SL g821 ( 
.A1(n_750),
.A2(n_760),
.B(n_755),
.C(n_773),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_756),
.Y(n_822)
);

OAI21x1_ASAP7_75t_L g823 ( 
.A1(n_726),
.A2(n_766),
.B(n_771),
.Y(n_823)
);

BUFx8_ASAP7_75t_L g824 ( 
.A(n_758),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_714),
.A2(n_691),
.B(n_727),
.C(n_740),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_728),
.B(n_747),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_735),
.A2(n_748),
.B(n_730),
.Y(n_827)
);

AOI22xp5_ASAP7_75t_L g828 ( 
.A1(n_710),
.A2(n_752),
.B1(n_712),
.B2(n_722),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_715),
.A2(n_776),
.B(n_733),
.C(n_757),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_695),
.A2(n_699),
.B(n_741),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_689),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_SL g832 ( 
.A1(n_723),
.A2(n_717),
.B(n_706),
.C(n_708),
.Y(n_832)
);

OAI21xp33_ASAP7_75t_L g833 ( 
.A1(n_723),
.A2(n_737),
.B(n_762),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_694),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_694),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_770),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_765),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_697),
.B(n_718),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_745),
.A2(n_718),
.B1(n_700),
.B2(n_731),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_718),
.A2(n_700),
.B1(n_731),
.B2(n_734),
.Y(n_840)
);

AO32x2_ASAP7_75t_L g841 ( 
.A1(n_734),
.A2(n_646),
.A3(n_761),
.B1(n_705),
.B2(n_725),
.Y(n_841)
);

AO31x2_ASAP7_75t_L g842 ( 
.A1(n_769),
.A2(n_738),
.A3(n_775),
.B(n_702),
.Y(n_842)
);

OR2x2_ASAP7_75t_L g843 ( 
.A(n_690),
.B(n_401),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_704),
.B(n_577),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_704),
.A2(n_707),
.B(n_582),
.C(n_705),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_698),
.A2(n_463),
.B1(n_582),
.B2(n_729),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_682),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_682),
.Y(n_848)
);

AO21x2_ASAP7_75t_L g849 ( 
.A1(n_738),
.A2(n_775),
.B(n_628),
.Y(n_849)
);

OAI221xp5_ASAP7_75t_L g850 ( 
.A1(n_704),
.A2(n_600),
.B1(n_696),
.B2(n_613),
.C(n_593),
.Y(n_850)
);

NAND2x1p5_ASAP7_75t_L g851 ( 
.A(n_690),
.B(n_680),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_682),
.Y(n_852)
);

AO31x2_ASAP7_75t_L g853 ( 
.A1(n_738),
.A2(n_775),
.A3(n_702),
.B(n_711),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_690),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_678),
.A2(n_463),
.B1(n_709),
.B2(n_478),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_704),
.B(n_598),
.Y(n_856)
);

OAI22x1_ASAP7_75t_L g857 ( 
.A1(n_677),
.A2(n_542),
.B1(n_462),
.B2(n_517),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_704),
.B(n_598),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_677),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_702),
.A2(n_653),
.B(n_652),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_707),
.A2(n_679),
.B(n_729),
.C(n_709),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_677),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_707),
.A2(n_679),
.B(n_729),
.C(n_709),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_704),
.B(n_647),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_680),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_707),
.A2(n_679),
.B(n_729),
.C(n_709),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_704),
.B(n_647),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_682),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_682),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_682),
.Y(n_870)
);

OAI22x1_ASAP7_75t_L g871 ( 
.A1(n_677),
.A2(n_542),
.B1(n_462),
.B2(n_517),
.Y(n_871)
);

OAI22xp33_ASAP7_75t_L g872 ( 
.A1(n_690),
.A2(n_401),
.B1(n_462),
.B2(n_542),
.Y(n_872)
);

AO31x2_ASAP7_75t_L g873 ( 
.A1(n_738),
.A2(n_775),
.A3(n_702),
.B(n_711),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_738),
.A2(n_775),
.A3(n_702),
.B(n_711),
.Y(n_874)
);

BUFx12f_ASAP7_75t_L g875 ( 
.A(n_677),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_682),
.Y(n_876)
);

AO32x2_ASAP7_75t_L g877 ( 
.A1(n_761),
.A2(n_646),
.A3(n_705),
.B1(n_725),
.B2(n_767),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_702),
.A2(n_653),
.B(n_652),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_707),
.A2(n_679),
.B(n_729),
.C(n_709),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_698),
.A2(n_463),
.B1(n_582),
.B2(n_729),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_696),
.A2(n_582),
.B1(n_597),
.B2(n_463),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_864),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_867),
.B(n_844),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_834),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_861),
.A2(n_866),
.B(n_863),
.C(n_879),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_834),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_843),
.B(n_800),
.Y(n_887)
);

AO31x2_ASAP7_75t_L g888 ( 
.A1(n_814),
.A2(n_813),
.A3(n_878),
.B(n_860),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_780),
.Y(n_889)
);

HB1xp67_ASAP7_75t_L g890 ( 
.A(n_808),
.Y(n_890)
);

CKINVDCx20_ASAP7_75t_R g891 ( 
.A(n_859),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_850),
.B(n_872),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_SL g893 ( 
.A1(n_881),
.A2(n_782),
.B1(n_862),
.B2(n_787),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_835),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_847),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_852),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_846),
.A2(n_880),
.B1(n_822),
.B2(n_871),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_869),
.B(n_870),
.Y(n_898)
);

OA21x2_ASAP7_75t_L g899 ( 
.A1(n_783),
.A2(n_823),
.B(n_784),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_SL g900 ( 
.A1(n_788),
.A2(n_803),
.B1(n_857),
.B2(n_856),
.Y(n_900)
);

OA21x2_ASAP7_75t_L g901 ( 
.A1(n_833),
.A2(n_786),
.B(n_829),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_855),
.A2(n_824),
.B1(n_817),
.B2(n_848),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_876),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_858),
.B(n_805),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_868),
.B(n_795),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_793),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_802),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_875),
.Y(n_908)
);

OAI222xp33_ASAP7_75t_L g909 ( 
.A1(n_828),
.A2(n_799),
.B1(n_798),
.B2(n_854),
.C1(n_818),
.C2(n_810),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_790),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_820),
.B(n_824),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_838),
.Y(n_912)
);

XOR2xp5_ASAP7_75t_L g913 ( 
.A(n_819),
.B(n_785),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_831),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_837),
.B(n_826),
.Y(n_915)
);

OA21x2_ASAP7_75t_L g916 ( 
.A1(n_833),
.A2(n_825),
.B(n_791),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_865),
.B(n_799),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_801),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_816),
.A2(n_840),
.B1(n_839),
.B2(n_794),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_806),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_836),
.B(n_830),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_827),
.B(n_815),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_807),
.B(n_812),
.Y(n_923)
);

OA21x2_ASAP7_75t_L g924 ( 
.A1(n_809),
.A2(n_797),
.B(n_804),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_781),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_SL g926 ( 
.A1(n_841),
.A2(n_792),
.B1(n_789),
.B2(n_877),
.Y(n_926)
);

AOI22xp33_ASAP7_75t_SL g927 ( 
.A1(n_792),
.A2(n_841),
.B1(n_877),
.B2(n_849),
.Y(n_927)
);

OA21x2_ASAP7_75t_L g928 ( 
.A1(n_842),
.A2(n_853),
.B(n_873),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_815),
.B(n_853),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_877),
.A2(n_853),
.B1(n_873),
.B2(n_874),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_796),
.B(n_864),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_SL g932 ( 
.A1(n_796),
.A2(n_401),
.B1(n_597),
.B2(n_778),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_864),
.B(n_867),
.Y(n_933)
);

AOI221xp5_ASAP7_75t_L g934 ( 
.A1(n_850),
.A2(n_582),
.B1(n_845),
.B2(n_872),
.C(n_704),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_864),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_881),
.A2(n_597),
.B1(n_850),
.B2(n_880),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_821),
.A2(n_832),
.B(n_878),
.Y(n_937)
);

CKINVDCx11_ASAP7_75t_R g938 ( 
.A(n_875),
.Y(n_938)
);

OR2x6_ASAP7_75t_L g939 ( 
.A(n_851),
.B(n_401),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_821),
.A2(n_832),
.B(n_878),
.Y(n_940)
);

AO31x2_ASAP7_75t_L g941 ( 
.A1(n_814),
.A2(n_813),
.A3(n_738),
.B(n_860),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_845),
.A2(n_863),
.B(n_866),
.C(n_861),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_821),
.A2(n_832),
.B(n_878),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_864),
.B(n_867),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_846),
.A2(n_462),
.B1(n_880),
.B2(n_855),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_881),
.A2(n_597),
.B1(n_850),
.B2(n_880),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_864),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_864),
.B(n_867),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_864),
.B(n_867),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_864),
.B(n_867),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_811),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_897),
.B(n_942),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_931),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_894),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_892),
.A2(n_934),
.B(n_923),
.C(n_946),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_891),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_921),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_925),
.Y(n_958)
);

BUFx2_ASAP7_75t_L g959 ( 
.A(n_951),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_951),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_897),
.B(n_942),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_889),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_944),
.B(n_933),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_937),
.A2(n_940),
.B(n_943),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_888),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_892),
.A2(n_936),
.B1(n_946),
.B2(n_945),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_885),
.B(n_930),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_895),
.Y(n_968)
);

OA21x2_ASAP7_75t_L g969 ( 
.A1(n_930),
.A2(n_929),
.B(n_922),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_885),
.B(n_926),
.Y(n_970)
);

OAI221xp5_ASAP7_75t_L g971 ( 
.A1(n_936),
.A2(n_932),
.B1(n_883),
.B2(n_949),
.C(n_948),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_896),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_950),
.B(n_912),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_927),
.B(n_928),
.Y(n_974)
);

AO21x2_ASAP7_75t_L g975 ( 
.A1(n_909),
.A2(n_919),
.B(n_923),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_912),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_927),
.B(n_928),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_916),
.B(n_907),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_903),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_884),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_932),
.B(n_882),
.Y(n_981)
);

OAI211xp5_ASAP7_75t_SL g982 ( 
.A1(n_935),
.A2(n_947),
.B(n_887),
.C(n_915),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_902),
.A2(n_939),
.B1(n_905),
.B2(n_890),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_L g984 ( 
.A1(n_917),
.A2(n_911),
.B(n_898),
.C(n_904),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_SL g985 ( 
.A1(n_900),
.A2(n_939),
.B1(n_893),
.B2(n_906),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_901),
.B(n_939),
.C(n_924),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_974),
.B(n_899),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_965),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_958),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_971),
.A2(n_910),
.B1(n_914),
.B2(n_920),
.C(n_913),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_974),
.B(n_941),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_960),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_977),
.B(n_941),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_977),
.B(n_941),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_977),
.B(n_924),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_953),
.B(n_918),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_957),
.Y(n_997)
);

INVxp67_ASAP7_75t_SL g998 ( 
.A(n_959),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_967),
.B(n_886),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_976),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_971),
.A2(n_908),
.B1(n_938),
.B2(n_966),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_952),
.B(n_961),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_978),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_952),
.B(n_961),
.Y(n_1004)
);

NOR2x1_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_984),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_989),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_988),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_R g1008 ( 
.A(n_1003),
.B(n_956),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_991),
.B(n_969),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_992),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_1002),
.B(n_967),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_993),
.B(n_970),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_993),
.B(n_969),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_993),
.B(n_969),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_992),
.B(n_973),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1002),
.B(n_970),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_1015),
.B(n_994),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1011),
.B(n_997),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_1016),
.B(n_984),
.Y(n_1019)
);

NOR2x1p5_ASAP7_75t_L g1020 ( 
.A(n_1015),
.B(n_998),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_1010),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_1005),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1006),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1009),
.B(n_987),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_1009),
.B(n_995),
.Y(n_1025)
);

INVxp67_ASAP7_75t_SL g1026 ( 
.A(n_1005),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_1007),
.Y(n_1027)
);

NOR2x1p5_ASAP7_75t_SL g1028 ( 
.A(n_1007),
.B(n_964),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_1009),
.B(n_987),
.Y(n_1029)
);

OR2x2_ASAP7_75t_L g1030 ( 
.A(n_1024),
.B(n_1013),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1024),
.B(n_1013),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_1027),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1019),
.B(n_1012),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1021),
.B(n_1012),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1029),
.B(n_1013),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1021),
.B(n_1014),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1023),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1027),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1029),
.B(n_1014),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1025),
.B(n_1014),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1025),
.B(n_1018),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1023),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_1026),
.A2(n_983),
.B(n_998),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_1031),
.B(n_1025),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1032),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_1043),
.B(n_1022),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_1032),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1038),
.Y(n_1048)
);

OAI31xp33_ASAP7_75t_L g1049 ( 
.A1(n_1033),
.A2(n_1020),
.A3(n_1022),
.B(n_1026),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_1034),
.Y(n_1050)
);

OAI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1036),
.A2(n_985),
.B(n_1001),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1038),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1037),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1041),
.B(n_1017),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1042),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_1051),
.A2(n_985),
.B1(n_1008),
.B2(n_1020),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_1046),
.A2(n_955),
.B(n_982),
.C(n_1001),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_SL g1058 ( 
.A(n_1049),
.B(n_1030),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1053),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1044),
.A2(n_1030),
.B1(n_1040),
.B2(n_1039),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1053),
.Y(n_1061)
);

NAND4xp75_ASAP7_75t_L g1062 ( 
.A(n_1044),
.B(n_990),
.C(n_981),
.D(n_1028),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1050),
.B(n_1031),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_1059),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1058),
.A2(n_990),
.B(n_1035),
.C(n_1054),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_SL g1066 ( 
.A1(n_1057),
.A2(n_982),
.B(n_980),
.C(n_954),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_1063),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_1056),
.A2(n_1035),
.B(n_1017),
.C(n_1055),
.Y(n_1068)
);

OAI311xp33_ASAP7_75t_L g1069 ( 
.A1(n_1062),
.A2(n_981),
.A3(n_1061),
.B1(n_1018),
.C1(n_1004),
.Y(n_1069)
);

NAND5xp2_ASAP7_75t_L g1070 ( 
.A(n_1060),
.B(n_961),
.C(n_970),
.D(n_999),
.E(n_1004),
.Y(n_1070)
);

AOI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1065),
.A2(n_1055),
.B1(n_983),
.B2(n_1048),
.C(n_1052),
.Y(n_1071)
);

NOR4xp25_ASAP7_75t_L g1072 ( 
.A(n_1069),
.B(n_979),
.C(n_968),
.D(n_972),
.Y(n_1072)
);

NOR3x1_ASAP7_75t_SL g1073 ( 
.A(n_1066),
.B(n_976),
.C(n_963),
.Y(n_1073)
);

NOR2x1p5_ASAP7_75t_L g1074 ( 
.A(n_1064),
.B(n_1047),
.Y(n_1074)
);

OAI211xp5_ASAP7_75t_SL g1075 ( 
.A1(n_1066),
.A2(n_963),
.B(n_1016),
.C(n_1000),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1075),
.B(n_1068),
.C(n_1070),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_L g1077 ( 
.A(n_1071),
.B(n_1067),
.C(n_986),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_L g1078 ( 
.A(n_1073),
.B(n_986),
.C(n_980),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_SL g1079 ( 
.A(n_1072),
.B(n_1011),
.C(n_968),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1079),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_1077),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1076),
.Y(n_1082)
);

OR4x2_ASAP7_75t_L g1083 ( 
.A(n_1078),
.B(n_1074),
.C(n_963),
.D(n_975),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1079),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1082),
.B(n_1045),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1080),
.A2(n_1084),
.B1(n_1081),
.B2(n_1083),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_1086),
.A2(n_1081),
.B(n_1083),
.Y(n_1087)
);

OAI222xp33_ASAP7_75t_L g1088 ( 
.A1(n_1087),
.A2(n_1085),
.B1(n_979),
.B2(n_972),
.C1(n_962),
.C2(n_1045),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1088),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_1089),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1090),
.A2(n_962),
.B(n_1047),
.Y(n_1091)
);


endmodule