module real_jpeg_2605_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_1),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_6),
.A2(n_26),
.B1(n_29),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_6),
.A2(n_45),
.B1(n_57),
.B2(n_59),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_6),
.B(n_17),
.C(n_38),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_6),
.B(n_24),
.C(n_26),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_17),
.B1(n_21),
.B2(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_6),
.B(n_46),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_6),
.B(n_67),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_7),
.A2(n_17),
.B1(n_21),
.B2(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_7),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_7),
.A2(n_34),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_78),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_76),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_52),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_12),
.B(n_52),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_35),
.C(n_40),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_13),
.A2(n_14),
.B1(n_35),
.B2(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_30),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_22),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_16),
.B(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_17),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_21),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NAND2x1_ASAP7_75t_SL g82 ( 
.A(n_17),
.B(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_29),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_39),
.B1(n_57),
.B2(n_59),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_40),
.A2(n_41),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_49),
.B(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_44),
.B(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_48),
.B(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_50),
.B(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_50),
.B(n_99),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_70),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_65),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_73),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_91),
.B(n_112),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_87),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_100),
.B(n_111),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_97),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_106),
.B(n_110),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_109),
.Y(n_110)
);


endmodule