module real_jpeg_11359_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_139;
wire n_33;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_1),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_2),
.A2(n_28),
.B1(n_31),
.B2(n_35),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_35),
.B1(n_86),
.B2(n_113),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_3),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_3),
.A2(n_11),
.B(n_24),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_4),
.A2(n_28),
.B1(n_31),
.B2(n_51),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_10),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_10),
.A2(n_23),
.B1(n_24),
.B2(n_63),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_10),
.A2(n_45),
.B1(n_46),
.B2(n_63),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_11),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_23),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_11),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_11),
.A2(n_84),
.B1(n_86),
.B2(n_113),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_11),
.A2(n_31),
.B(n_57),
.C(n_65),
.D(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_11),
.B(n_31),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_27),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_11),
.A2(n_91),
.B(n_139),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g165 ( 
.A1(n_11),
.A2(n_23),
.B(n_36),
.C(n_72),
.D(n_166),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_12),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_13),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_13),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_14),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_14),
.A2(n_25),
.B1(n_28),
.B2(n_31),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_14),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_119),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_117),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_18),
.B(n_79),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_55),
.C(n_68),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_19),
.B(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_38),
.B2(n_54),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_20),
.B(n_39),
.C(n_43),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_32),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_22),
.A2(n_26),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_SL g36 ( 
.A1(n_24),
.A2(n_27),
.B(n_29),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_26),
.B(n_34),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_28),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_28),
.B(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_28),
.A2(n_37),
.B1(n_71),
.B2(n_73),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_29),
.B(n_31),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_36),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_40),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_42),
.B(n_86),
.C(n_111),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_42),
.B(n_86),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_44),
.A2(n_49),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_45),
.B(n_58),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_45),
.B(n_155),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_46),
.A2(n_60),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_49),
.B(n_78),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_55),
.A2(n_68),
.B1(n_69),
.B2(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_55),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_64),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_56),
.A2(n_62),
.B1(n_66),
.B2(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_66),
.A2(n_101),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_66),
.B(n_84),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_74),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_70),
.B(n_74),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_76),
.B(n_77),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_76),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_76),
.A2(n_77),
.B(n_144),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_76),
.B(n_84),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_97),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_91),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_94),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_112),
.B(n_114),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_172),
.B(n_177),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_159),
.B(n_171),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_140),
.B(n_158),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_130),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_123),
.B(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_126),
.B1(n_127),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_135),
.C(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_138),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_148),
.B(n_157),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_146),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_152),
.B(n_156),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_151),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_160),
.B(n_161),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_169),
.B2(n_170),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_164),
.Y(n_168)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_165),
.B(n_168),
.C(n_170),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_169),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_173),
.B(n_174),
.Y(n_177)
);


endmodule