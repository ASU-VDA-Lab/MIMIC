module real_jpeg_15071_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_4),
.A2(n_32),
.B1(n_54),
.B2(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_73),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_5),
.A2(n_54),
.B1(n_56),
.B2(n_73),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_73),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_6),
.A2(n_34),
.B1(n_54),
.B2(n_56),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_8),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_54),
.B1(n_56),
.B2(n_62),
.Y(n_120)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_10),
.A2(n_36),
.B(n_37),
.C(n_42),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_10),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_10),
.B(n_113),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_39),
.B1(n_54),
.B2(n_56),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_10),
.A2(n_98),
.B1(n_102),
.B2(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_60),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_11),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_11),
.A2(n_40),
.B1(n_41),
.B2(n_70),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_70),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_70),
.Y(n_185)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_13),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_54),
.B1(n_56),
.B2(n_83),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_83),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_49),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_14),
.A2(n_49),
.B1(n_54),
.B2(n_56),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_49),
.Y(n_179)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_114),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_114),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_46),
.C(n_63),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_21),
.A2(n_22),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_35),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_23),
.A2(n_24),
.B1(n_35),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_25),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_25),
.A2(n_79),
.B(n_101),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_25),
.A2(n_29),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_26),
.A2(n_27),
.B1(n_89),
.B2(n_90),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_26),
.B(n_39),
.C(n_90),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_26),
.B(n_183),
.Y(n_182)
);

CKINVDCx6p67_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_29),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_31),
.A2(n_80),
.B(n_102),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_35),
.Y(n_211)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B(n_40),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g140 ( 
.A(n_39),
.B(n_41),
.CON(n_140),
.SN(n_140)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_39),
.B(n_102),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_39),
.B(n_91),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_41),
.B1(n_53),
.B2(n_57),
.Y(n_58)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_40),
.B(n_54),
.C(n_57),
.Y(n_141)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_46),
.B(n_63),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_59),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_48),
.A2(n_51),
.B1(n_60),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_50),
.A2(n_52),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_51),
.A2(n_61),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_51),
.A2(n_60),
.B1(n_140),
.B2(n_151),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_110),
.Y(n_109)
);

OA22x2_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_53),
.A2(n_56),
.B(n_139),
.C(n_141),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_54),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_56),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_56),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_72),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_65),
.A2(n_69),
.B1(n_113),
.B2(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_95),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_84),
.B2(n_94),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_78),
.A2(n_98),
.B(n_179),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_91),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_87),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_87),
.A2(n_92),
.B1(n_146),
.B2(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_87),
.A2(n_92),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_87),
.A2(n_92),
.B1(n_162),
.B2(n_172),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_89),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_91),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_120),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_103),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_97),
.B(n_103),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_98),
.A2(n_102),
.B1(n_177),
.B2(n_185),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_126),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_115),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_118),
.B(n_126),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_124),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_119),
.B(n_122),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_123),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_124),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_221),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_217),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_207),
.B(n_216),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_163),
.B(n_206),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_158),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_135),
.B(n_158),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_148),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_137),
.B(n_143),
.C(n_148),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_142),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_145),
.B(n_147),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_149),
.B(n_154),
.C(n_157),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.C(n_161),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_159),
.B(n_203),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_160),
.B(n_161),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_201),
.B(n_205),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_191),
.B(n_200),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_180),
.B(n_190),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_175),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_173),
.B2(n_174),
.Y(n_167)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_170),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_173),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_189),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.C(n_199),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_204),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_215),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_215),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_212),
.C(n_213),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_220),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);


endmodule