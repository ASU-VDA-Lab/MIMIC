module real_jpeg_30367_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_1),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_0),
.B(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_2),
.A2(n_7),
.B1(n_27),
.B2(n_31),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_3),
.B(n_12),
.Y(n_11)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

OAI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_9),
.B1(n_20),
.B2(n_22),
.C(n_26),
.Y(n_6)
);

INVx1_ASAP7_75t_SL g7 ( 
.A(n_8),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_14),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_13),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_24),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_17),
.B(n_18),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);


endmodule