module fake_jpeg_17133_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_45),
.B(n_38),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_65),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_57),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_19),
.B1(n_17),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_25),
.B1(n_31),
.B2(n_16),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_19),
.B1(n_17),
.B2(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_62),
.B1(n_28),
.B2(n_23),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_20),
.B1(n_30),
.B2(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_32),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_61),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_70),
.B(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_74),
.A2(n_49),
.B1(n_44),
.B2(n_40),
.Y(n_114)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_31),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_54),
.A2(n_17),
.B1(n_22),
.B2(n_24),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_65),
.B(n_31),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_53),
.B(n_52),
.Y(n_109)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_23),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_28),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_90),
.B(n_92),
.C(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_52),
.B1(n_44),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_103),
.A2(n_68),
.B1(n_70),
.B2(n_74),
.Y(n_140)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_89),
.A2(n_40),
.A3(n_55),
.B1(n_47),
.B2(n_50),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_109),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_76),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_115),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp33_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_59),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_118),
.B(n_119),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_80),
.C(n_92),
.Y(n_138)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_131),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_84),
.B1(n_87),
.B2(n_73),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_140),
.B1(n_95),
.B2(n_88),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_79),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_146),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_101),
.B(n_86),
.C(n_71),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_142),
.C(n_103),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_69),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_137),
.B(n_139),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_20),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_100),
.B(n_72),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_141),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_86),
.C(n_71),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_96),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_143),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_144),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_97),
.B1(n_87),
.B2(n_88),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_74),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_116),
.A2(n_77),
.B1(n_63),
.B2(n_73),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_83),
.B1(n_119),
.B2(n_106),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_SL g148 ( 
.A1(n_99),
.A2(n_82),
.B(n_93),
.C(n_85),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_94),
.B(n_102),
.Y(n_159)
);

AO22x1_ASAP7_75t_SL g150 ( 
.A1(n_135),
.A2(n_104),
.B1(n_112),
.B2(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_150),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_134),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_151),
.B(n_152),
.C(n_153),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_146),
.C(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_160),
.B1(n_168),
.B2(n_127),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_145),
.B1(n_125),
.B2(n_122),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_162),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_128),
.A2(n_97),
.B1(n_110),
.B2(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_67),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_98),
.C(n_110),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_165),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_67),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_66),
.B1(n_41),
.B2(n_25),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_147),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_98),
.B(n_18),
.C(n_66),
.D(n_27),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_174),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_98),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_130),
.B(n_148),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_126),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_192),
.B1(n_201),
.B2(n_171),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_123),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_177),
.B(n_183),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_185),
.B(n_187),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_132),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_144),
.Y(n_188)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_188),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_189),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_193),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_155),
.A2(n_148),
.B1(n_143),
.B2(n_129),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_127),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_163),
.B1(n_156),
.B2(n_170),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_196),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_148),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_197),
.Y(n_207)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_167),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_98),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_199),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_160),
.B(n_141),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_162),
.B(n_168),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_126),
.B1(n_123),
.B2(n_30),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_203),
.B1(n_216),
.B2(n_224),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_195),
.A2(n_159),
.B1(n_150),
.B2(n_154),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_151),
.C(n_191),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_213),
.C(n_222),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_226),
.B1(n_194),
.B2(n_187),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_152),
.Y(n_213)
);

AOI211xp5_ASAP7_75t_SL g216 ( 
.A1(n_197),
.A2(n_150),
.B(n_169),
.C(n_165),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_27),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_225),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_182),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_27),
.C(n_18),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_223),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_178),
.A2(n_29),
.B1(n_26),
.B2(n_24),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_18),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_179),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_229),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_208),
.B(n_196),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_211),
.A2(n_187),
.B1(n_178),
.B2(n_200),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_230),
.A2(n_209),
.B1(n_215),
.B2(n_226),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_186),
.C(n_193),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_237),
.C(n_247),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_180),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_234),
.B(n_235),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_180),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_185),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_241),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_186),
.C(n_201),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_190),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_243),
.B(n_246),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_176),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_203),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_192),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_175),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_198),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_208),
.B(n_202),
.C(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_233),
.A2(n_215),
.B(n_209),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_261),
.B(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_263),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_259),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_258),
.B(n_262),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_182),
.C(n_216),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_265),
.C(n_266),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_183),
.B(n_224),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_248),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_20),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_29),
.C(n_1),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_227),
.C(n_239),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_8),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_254),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_260),
.C(n_266),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_272),
.B(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_257),
.B(n_245),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_247),
.B1(n_229),
.B2(n_239),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_8),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_275),
.B(n_11),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_8),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_279),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_0),
.C(n_1),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_280),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_9),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_3),
.C(n_4),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_280),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_249),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_272),
.C(n_269),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_271),
.B(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_292),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_291),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_294),
.B(n_296),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_268),
.B(n_15),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_12),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_268),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_301),
.C(n_305),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_283),
.B(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_307),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_9),
.C(n_14),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_12),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_12),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_3),
.C(n_5),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_287),
.B(n_5),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_297),
.B(n_303),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_6),
.B1(n_7),
.B2(n_312),
.Y(n_324)
);

OAI21x1_ASAP7_75t_L g314 ( 
.A1(n_301),
.A2(n_294),
.B(n_15),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_314),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_15),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_3),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_6),
.B(n_7),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_5),
.B(n_6),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.C(n_324),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_6),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_311),
.C(n_7),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_326),
.A2(n_327),
.B1(n_323),
.B2(n_325),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_328),
.B(n_319),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_329),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_319),
.Y(n_331)
);


endmodule