module real_jpeg_15005_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_3),
.A2(n_33),
.B1(n_36),
.B2(n_92),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_52),
.B1(n_53),
.B2(n_92),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_45),
.B1(n_49),
.B2(n_92),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_4),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_4),
.A2(n_33),
.B1(n_36),
.B2(n_133),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_4),
.A2(n_52),
.B1(n_53),
.B2(n_133),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_4),
.A2(n_45),
.B1(n_49),
.B2(n_133),
.Y(n_259)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_6),
.A2(n_33),
.B1(n_36),
.B2(n_184),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_6),
.A2(n_52),
.B1(n_53),
.B2(n_184),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_6),
.A2(n_45),
.B1(n_49),
.B2(n_184),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_7),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_7),
.A2(n_30),
.B1(n_52),
.B2(n_53),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_30),
.B1(n_45),
.B2(n_49),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_9),
.A2(n_45),
.B1(n_49),
.B2(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_33),
.B1(n_36),
.B2(n_55),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_12),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_12),
.A2(n_33),
.B1(n_36),
.B2(n_157),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_157),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_12),
.A2(n_45),
.B1(n_49),
.B2(n_157),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_13),
.A2(n_33),
.B1(n_36),
.B2(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_13),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_13),
.A2(n_52),
.B1(n_53),
.B2(n_59),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_59),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_45),
.B1(n_49),
.B2(n_59),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_14),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_14),
.A2(n_27),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_14),
.B(n_187),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_14),
.B(n_36),
.Y(n_235)
);

OAI22xp33_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_176),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_14),
.A2(n_48),
.B(n_52),
.C(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_14),
.B(n_69),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_85),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_14),
.B(n_43),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_L g285 ( 
.A1(n_14),
.A2(n_36),
.B(n_235),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_15),
.A2(n_33),
.B1(n_36),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_15),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_15),
.A2(n_45),
.B1(n_49),
.B2(n_68),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_16),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_16),
.A2(n_33),
.B1(n_36),
.B2(n_39),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_16),
.A2(n_39),
.B1(n_52),
.B2(n_53),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_16),
.A2(n_39),
.B1(n_45),
.B2(n_49),
.Y(n_172)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_105),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_93),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_22),
.B(n_93),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_71),
.C(n_78),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_23),
.A2(n_71),
.B1(n_72),
.B2(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_24),
.A2(n_25),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_42),
.C(n_57),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_26),
.A2(n_31),
.B1(n_32),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g173 ( 
.A1(n_27),
.A2(n_33),
.A3(n_35),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_28),
.B(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_31),
.A2(n_32),
.B1(n_38),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_31),
.A2(n_32),
.B1(n_91),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_31),
.A2(n_32),
.B1(n_132),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_31),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_31),
.A2(n_32),
.B1(n_183),
.B2(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_37),
.Y(n_31)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_32),
.Y(n_187)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_33),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_34),
.B(n_36),
.Y(n_174)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI32xp33_ASAP7_75t_L g233 ( 
.A1(n_36),
.A2(n_53),
.A3(n_64),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_56),
.B1(n_57),
.B2(n_70),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_42),
.A2(n_70),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_50),
.B(n_54),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_43),
.A2(n_50),
.B1(n_54),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_50),
.B1(n_74),
.B2(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_43),
.A2(n_50),
.B1(n_89),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_43),
.A2(n_50),
.B1(n_151),
.B2(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_43),
.A2(n_50),
.B1(n_202),
.B2(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_43),
.A2(n_50),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_43),
.A2(n_50),
.B1(n_250),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_44),
.A2(n_128),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_44),
.A2(n_152),
.B1(n_229),
.B2(n_287),
.Y(n_286)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_44)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_45),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_45),
.B(n_273),
.Y(n_272)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_47),
.A2(n_49),
.B(n_176),
.Y(n_252)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_50),
.Y(n_152)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_52),
.B(n_63),
.Y(n_236)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_60),
.B1(n_66),
.B2(n_69),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_58),
.A2(n_60),
.B1(n_69),
.B2(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_60),
.A2(n_69),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_60),
.A2(n_69),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_62),
.B1(n_67),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_62),
.B1(n_77),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_61),
.A2(n_62),
.B1(n_130),
.B2(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_61),
.A2(n_62),
.B1(n_179),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_61),
.A2(n_62),
.B1(n_210),
.B2(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_62),
.Y(n_69)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_90),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_80),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_82),
.B1(n_90),
.B2(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_86),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_83),
.A2(n_85),
.B1(n_86),
.B2(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_83),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_83),
.A2(n_85),
.B1(n_148),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_83),
.A2(n_85),
.B1(n_172),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_83),
.A2(n_85),
.B1(n_214),
.B2(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_83),
.A2(n_85),
.B1(n_238),
.B2(n_259),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_83),
.A2(n_85),
.B1(n_176),
.B2(n_271),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_83),
.A2(n_85),
.B1(n_264),
.B2(n_271),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_84),
.A2(n_124),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_84),
.A2(n_146),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_90),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_134),
.B(n_307),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_107),
.B(n_110),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_118),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_129),
.C(n_131),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_120),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_121),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_160),
.B(n_306),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_158),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_137),
.B(n_158),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.C(n_142),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_141),
.Y(n_189)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_189),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.C(n_155),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_144),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_145),
.B(n_149),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_153),
.B(n_155),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_190),
.B(n_305),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_188),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_162),
.B(n_188),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.C(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_167),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_168),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_177),
.C(n_181),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_173),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_181),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_221),
.B(n_299),
.C(n_304),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_215),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_192),
.B(n_215),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_205),
.C(n_207),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_194),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_199),
.C(n_204),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_199),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_205),
.B(n_207),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_213),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_208),
.B(n_226),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_213),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_298),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_242),
.B(n_297),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_239),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_224),
.B(n_239),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.C(n_230),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_227),
.A2(n_230),
.B1(n_231),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_227),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_237),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_232),
.A2(n_233),
.B1(n_237),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_237),
.Y(n_289)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_291),
.B(n_296),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_244),
.A2(n_280),
.B(n_290),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_260),
.B(n_279),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_253),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_246),
.B(n_253),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_256),
.C(n_258),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_259),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_268),
.B(n_278),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_262),
.B(n_266),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B(n_277),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_281),
.B(n_282),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_288),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_286),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_286),
.C(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_293),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);


endmodule