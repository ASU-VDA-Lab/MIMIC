module fake_jpeg_8362_n_76 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_76);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_76;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_75;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_70;
wire n_15;
wire n_66;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_19),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_21),
.Y(n_23)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_13),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_20),
.B1(n_21),
.B2(n_12),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_21),
.C(n_17),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_17),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_12),
.B(n_18),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_9),
.B(n_10),
.C(n_8),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_20),
.B1(n_13),
.B2(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_24),
.B1(n_21),
.B2(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_8),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_10),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

OAI22x1_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_17),
.B1(n_9),
.B2(n_16),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_27),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_37),
.B1(n_24),
.B2(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_11),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_37),
.C(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_53),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_48),
.A2(n_50),
.B1(n_43),
.B2(n_11),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_35),
.C(n_28),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_52),
.C(n_41),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_35),
.C(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_17),
.C(n_16),
.Y(n_64)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_15),
.B1(n_14),
.B2(n_17),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_16),
.B1(n_1),
.B2(n_3),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_49),
.A2(n_14),
.B1(n_16),
.B2(n_3),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_5),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_56),
.B1(n_57),
.B2(n_6),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_62),
.A2(n_58),
.B(n_5),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_55),
.C(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_65),
.B(n_67),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_68),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_64),
.C(n_60),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_6),
.B(n_7),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_69),
.A2(n_62),
.B1(n_61),
.B2(n_7),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_73),
.C(n_70),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_6),
.B(n_0),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_0),
.Y(n_76)
);


endmodule