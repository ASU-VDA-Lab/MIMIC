module fake_jpeg_12926_n_158 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_27),
.B(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_21),
.Y(n_68)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_30),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_62),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_62),
.B1(n_72),
.B2(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_0),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_85),
.Y(n_86)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_65),
.B1(n_76),
.B2(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_76),
.B1(n_74),
.B2(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_81),
.A2(n_54),
.B1(n_75),
.B2(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_70),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_95),
.B(n_97),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_60),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_86),
.B(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_99),
.B(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_57),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_104),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_58),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_89),
.B(n_71),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_63),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_87),
.B(n_88),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_113),
.C(n_19),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_61),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_66),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_79),
.B1(n_68),
.B2(n_67),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_69),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_114),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_69),
.C(n_55),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_2),
.B(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_122),
.B(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_4),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_108),
.B(n_5),
.C(n_8),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_34),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_111),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_25),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_130),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_103),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_121),
.B(n_28),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_32),
.C(n_33),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_142),
.C(n_117),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_48),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_137),
.A2(n_42),
.B(n_45),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_38),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_117),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_40),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_134),
.C(n_132),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_150),
.A2(n_147),
.B(n_146),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_150),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_152),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_148),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_149),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_138),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_156),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_145),
.CI(n_139),
.CON(n_158),
.SN(n_158)
);


endmodule