module fake_netlist_5_2043_n_1928 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1928);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1928;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_87),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_72),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_103),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_83),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_43),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_60),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_69),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_35),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_100),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_109),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_53),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_31),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_65),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_146),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_95),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_23),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_5),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_38),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_23),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_52),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_159),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_27),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_31),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_19),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_74),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_94),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_30),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_2),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_136),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_39),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_0),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_99),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_137),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_92),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_178),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_45),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_182),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_73),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_56),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_54),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_67),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_70),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_143),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_8),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_53),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_11),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_30),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_122),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_59),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_163),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_66),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_106),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_88),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_165),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_7),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_34),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_6),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_12),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_18),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_78),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_26),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_149),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_66),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_120),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_180),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_79),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_114),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_81),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_144),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_184),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_130),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_24),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_89),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_157),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_35),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_152),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_189),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_147),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_179),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_90),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_9),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_42),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_62),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_176),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_164),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_126),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_15),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_2),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_68),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_39),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_140),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_17),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_50),
.Y(n_299)
);

BUFx5_ASAP7_75t_L g300 ( 
.A(n_183),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_141),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_86),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_118),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_71),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_128),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_127),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

BUFx10_ASAP7_75t_L g308 ( 
.A(n_139),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_167),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_187),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_138),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_82),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_47),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_20),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_26),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_62),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_52),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_42),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_47),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_29),
.Y(n_320)
);

INVx4_ASAP7_75t_R g321 ( 
.A(n_132),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_104),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_51),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_64),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_19),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_186),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_169),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_32),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_150),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_21),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_21),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_60),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_172),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_13),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_17),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_145),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_11),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_135),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_64),
.Y(n_340)
);

BUFx5_ASAP7_75t_L g341 ( 
.A(n_148),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_107),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_123),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_91),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_111),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_8),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_9),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_27),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_113),
.Y(n_349)
);

BUFx8_ASAP7_75t_SL g350 ( 
.A(n_0),
.Y(n_350)
);

BUFx5_ASAP7_75t_L g351 ( 
.A(n_162),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_5),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_133),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_59),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_63),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_57),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_48),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_45),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_171),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_119),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_10),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_44),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_51),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_112),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_108),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_134),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_117),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_4),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_96),
.Y(n_369)
);

BUFx10_ASAP7_75t_L g370 ( 
.A(n_84),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_28),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_16),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_7),
.Y(n_373)
);

BUFx10_ASAP7_75t_L g374 ( 
.A(n_4),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_57),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_76),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_158),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_12),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_43),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_38),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_350),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_270),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_191),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_312),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_270),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_312),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_258),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_266),
.Y(n_388)
);

INVxp33_ASAP7_75t_SL g389 ( 
.A(n_206),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_268),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_193),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_205),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_205),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_376),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_205),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_194),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_195),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_198),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_222),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_206),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_223),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_227),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_205),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_205),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_205),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_205),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_207),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g408 ( 
.A(n_293),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_359),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_359),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_207),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_207),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_207),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_233),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_207),
.Y(n_415)
);

INVxp33_ASAP7_75t_SL g416 ( 
.A(n_210),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_207),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_207),
.Y(n_418)
);

INVxp67_ASAP7_75t_SL g419 ( 
.A(n_365),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_356),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_365),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_356),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_248),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_332),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_235),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_248),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_293),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_281),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_300),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_293),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_281),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_301),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_374),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_238),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_239),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_358),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_240),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_358),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_263),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_263),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_264),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_264),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_288),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_247),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_288),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_300),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_318),
.Y(n_452)
);

INVxp33_ASAP7_75t_SL g453 ( 
.A(n_210),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_318),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_214),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_379),
.Y(n_457)
);

INVxp33_ASAP7_75t_SL g458 ( 
.A(n_214),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_379),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_203),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_202),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_257),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_216),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_220),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_221),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_374),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_224),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_225),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_374),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_259),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_243),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_267),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_250),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_251),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_261),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_392),
.B(n_342),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_392),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_383),
.B(n_360),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_460),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_393),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_420),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_420),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_393),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_422),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_423),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_395),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_391),
.B(n_360),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_403),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_403),
.B(n_342),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_387),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_404),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_423),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

AND2x2_ASAP7_75t_SL g498 ( 
.A(n_394),
.B(n_196),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_384),
.A2(n_197),
.B1(n_229),
.B2(n_213),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_396),
.B(n_196),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_426),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_386),
.A2(n_319),
.B1(n_213),
.B2(n_197),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_406),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_397),
.B(n_209),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_424),
.B(n_255),
.Y(n_506)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_406),
.A2(n_274),
.B(n_255),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_408),
.B(n_429),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_398),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_399),
.B(n_274),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_401),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_424),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_390),
.A2(n_368),
.B1(n_254),
.B2(n_319),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_402),
.B(n_192),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_382),
.B(n_237),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_407),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_407),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_427),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_439),
.B(n_192),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_389),
.A2(n_254),
.B1(n_229),
.B2(n_375),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_432),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_440),
.B(n_283),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_411),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_412),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_460),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_462),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_470),
.B(n_201),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_434),
.B(n_283),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_385),
.B(n_409),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_434),
.B(n_230),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_400),
.B(n_201),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_410),
.B(n_231),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_441),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_438),
.B(n_296),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_461),
.B(n_237),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_414),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_433),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_413),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_419),
.B(n_421),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_415),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_457),
.B(n_203),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_457),
.B(n_203),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_415),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_441),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_417),
.A2(n_244),
.B(n_232),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_442),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_435),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_417),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_456),
.B(n_246),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_520),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_544),
.B(n_505),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_498),
.A2(n_296),
.B1(n_375),
.B2(n_368),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_477),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_477),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_477),
.Y(n_561)
);

BUFx8_ASAP7_75t_SL g562 ( 
.A(n_493),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_SL g563 ( 
.A1(n_539),
.A2(n_469),
.B1(n_466),
.B2(n_453),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_480),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_480),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_544),
.B(n_436),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_480),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_487),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_484),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_478),
.B(n_416),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_484),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_500),
.B(n_443),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_486),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_486),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_486),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_517),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_517),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_517),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_490),
.B(n_458),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_543),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_476),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_543),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_545),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_533),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_553),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_533),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_553),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_514),
.B(n_449),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_532),
.A2(n_550),
.B(n_524),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_510),
.B(n_443),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_489),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_553),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_552),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_555),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_489),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_533),
.B(n_506),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_489),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_489),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_489),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_509),
.Y(n_607)
);

AND3x2_ASAP7_75t_L g608 ( 
.A(n_539),
.B(n_437),
.C(n_435),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_489),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_495),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_515),
.A2(n_287),
.B1(n_289),
.B2(n_262),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_521),
.B(n_472),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_491),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_495),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_541),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_552),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_381),
.Y(n_617)
);

INVxp67_ASAP7_75t_SL g618 ( 
.A(n_491),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_491),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_546),
.B(n_547),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_491),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_491),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_535),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_546),
.B(n_456),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_491),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_494),
.Y(n_627)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_498),
.A2(n_308),
.B1(n_370),
.B2(n_246),
.Y(n_628)
);

NOR2xp67_ASAP7_75t_L g629 ( 
.A(n_495),
.B(n_269),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_548),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_494),
.Y(n_631)
);

INVxp33_ASAP7_75t_L g632 ( 
.A(n_513),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_551),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_548),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_548),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_494),
.Y(n_636)
);

XOR2x2_ASAP7_75t_L g637 ( 
.A(n_499),
.B(n_234),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_548),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_513),
.A2(n_354),
.B1(n_355),
.B2(n_380),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_494),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_494),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_547),
.B(n_459),
.Y(n_642)
);

BUFx2_ASAP7_75t_L g643 ( 
.A(n_540),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_494),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_271),
.Y(n_645)
);

NAND2x1p5_ASAP7_75t_L g646 ( 
.A(n_550),
.B(n_245),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_540),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_497),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_497),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_522),
.A2(n_215),
.B1(n_219),
.B2(n_354),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_554),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_497),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_497),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_479),
.B(n_272),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_511),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_537),
.A2(n_324),
.B1(n_326),
.B2(n_329),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_497),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_497),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_533),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_501),
.B(n_273),
.Y(n_660)
);

INVx6_ASAP7_75t_L g661 ( 
.A(n_501),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_501),
.B(n_275),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_550),
.A2(n_314),
.B1(n_373),
.B2(n_299),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_501),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_528),
.B(n_437),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_504),
.B(n_276),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_504),
.Y(n_668)
);

OAI22xp33_ASAP7_75t_SL g669 ( 
.A1(n_540),
.A2(n_357),
.B1(n_347),
.B2(n_336),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_504),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_502),
.B(n_246),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_504),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_504),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_518),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_518),
.Y(n_676)
);

AND3x2_ASAP7_75t_L g677 ( 
.A(n_525),
.B(n_253),
.C(n_249),
.Y(n_677)
);

NOR2x1p5_ASAP7_75t_L g678 ( 
.A(n_554),
.B(n_215),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_518),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_518),
.Y(n_681)
);

AND2x6_ASAP7_75t_L g682 ( 
.A(n_506),
.B(n_342),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_518),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_519),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_519),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_476),
.B(n_342),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_519),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_550),
.A2(n_335),
.B1(n_320),
.B2(n_315),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_540),
.B(n_425),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_519),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_519),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_519),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_540),
.B(n_428),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_529),
.B(n_308),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_493),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_526),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_526),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_481),
.B(n_430),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_526),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_506),
.B(n_265),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_476),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_526),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_526),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_506),
.Y(n_704)
);

INVx4_ASAP7_75t_L g705 ( 
.A(n_587),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_557),
.B(n_508),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_704),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_651),
.B(n_598),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_570),
.B(n_522),
.Y(n_709)
);

O2A1O1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_566),
.A2(n_459),
.B(n_461),
.C(n_468),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_620),
.B(n_204),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_704),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_598),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_651),
.B(n_526),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_616),
.Y(n_715)
);

AOI22xp5_ASAP7_75t_L g716 ( 
.A1(n_580),
.A2(n_302),
.B1(n_278),
.B2(n_279),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_573),
.B(n_204),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_616),
.B(n_499),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_628),
.B(n_208),
.Y(n_719)
);

OAI221xp5_ASAP7_75t_L g720 ( 
.A1(n_656),
.A2(n_286),
.B1(n_290),
.B2(n_291),
.C(n_292),
.Y(n_720)
);

AND2x2_ASAP7_75t_SL g721 ( 
.A(n_558),
.B(n_643),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_607),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_587),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_595),
.B(n_527),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_666),
.B(n_208),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_689),
.B(n_211),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_559),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_625),
.B(n_527),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_678),
.A2(n_306),
.B1(n_280),
.B2(n_282),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_587),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_591),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_588),
.B(n_211),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_559),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_678),
.A2(n_344),
.B1(n_284),
.B2(n_285),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_558),
.A2(n_380),
.B1(n_355),
.B2(n_219),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_591),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_624),
.B(n_212),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_591),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_689),
.B(n_212),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_659),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_624),
.B(n_217),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_SL g742 ( 
.A(n_556),
.B(n_503),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_625),
.B(n_527),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_642),
.B(n_594),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_642),
.B(n_527),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_655),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_693),
.B(n_217),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_527),
.Y(n_748)
);

NAND3xp33_ASAP7_75t_L g749 ( 
.A(n_611),
.B(n_200),
.C(n_199),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_659),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_603),
.B(n_534),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_603),
.B(n_534),
.Y(n_752)
);

AND2x6_ASAP7_75t_L g753 ( 
.A(n_659),
.B(n_297),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_615),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_568),
.B(n_463),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_603),
.B(n_534),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_560),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_610),
.B(n_614),
.Y(n_758)
);

INVxp33_ASAP7_75t_L g759 ( 
.A(n_568),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_614),
.B(n_534),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_571),
.B(n_463),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_571),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_617),
.B(n_218),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_593),
.B(n_464),
.Y(n_764)
);

INVx4_ASAP7_75t_L g765 ( 
.A(n_657),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_622),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_622),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_630),
.B(n_534),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_698),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_693),
.B(n_218),
.Y(n_770)
);

O2A1O1Ixp33_ASAP7_75t_L g771 ( 
.A1(n_669),
.A2(n_464),
.B(n_465),
.C(n_475),
.Y(n_771)
);

OR2x2_ASAP7_75t_L g772 ( 
.A(n_695),
.B(n_503),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_630),
.B(n_534),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_634),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_634),
.B(n_536),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_663),
.A2(n_688),
.B(n_700),
.C(n_638),
.Y(n_776)
);

NAND2xp33_ASAP7_75t_L g777 ( 
.A(n_682),
.B(n_646),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_700),
.B(n_536),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_624),
.B(n_303),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_635),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_624),
.B(n_303),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_700),
.B(n_536),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_700),
.B(n_536),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_536),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_638),
.B(n_536),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_643),
.A2(n_309),
.B1(n_311),
.B2(n_322),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_694),
.B(n_304),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_629),
.B(n_531),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_657),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_612),
.B(n_304),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_629),
.B(n_531),
.Y(n_791)
);

INVx8_ASAP7_75t_L g792 ( 
.A(n_633),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_645),
.B(n_305),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_561),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_669),
.B(n_305),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_682),
.B(n_300),
.Y(n_796)
);

INVx8_ASAP7_75t_L g797 ( 
.A(n_562),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_654),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_661),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_564),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_647),
.B(n_295),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_608),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_672),
.B(n_226),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_677),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_618),
.B(n_531),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_647),
.B(n_328),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_565),
.A2(n_327),
.B(n_310),
.C(n_330),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_657),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_641),
.B(n_507),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_641),
.B(n_507),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_640),
.B(n_465),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_567),
.A2(n_337),
.B(n_377),
.C(n_353),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_660),
.A2(n_369),
.B1(n_364),
.B2(n_345),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_652),
.B(n_507),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_632),
.B(n_228),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_564),
.Y(n_817)
);

A2O1A1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_567),
.A2(n_334),
.B(n_339),
.C(n_343),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_662),
.B(n_236),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_564),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_563),
.B(n_467),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_652),
.B(n_507),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_650),
.B(n_349),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_658),
.B(n_481),
.Y(n_824)
);

NAND3xp33_ASAP7_75t_L g825 ( 
.A(n_650),
.B(n_256),
.C(n_241),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_658),
.B(n_482),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_667),
.B(n_664),
.Y(n_827)
);

OR2x6_ASAP7_75t_L g828 ( 
.A(n_646),
.B(n_467),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_639),
.Y(n_829)
);

NOR2xp67_ASAP7_75t_L g830 ( 
.A(n_639),
.B(n_640),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_664),
.B(n_665),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_665),
.B(n_482),
.Y(n_832)
);

O2A1O1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_646),
.A2(n_468),
.B(n_471),
.C(n_473),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_668),
.B(n_483),
.Y(n_834)
);

O2A1O1Ixp5_ASAP7_75t_L g835 ( 
.A1(n_569),
.A2(n_451),
.B(n_431),
.C(n_523),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_569),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_582),
.B(n_366),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_637),
.A2(n_300),
.B1(n_341),
.B2(n_351),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_582),
.B(n_367),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_582),
.B(n_308),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_637),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_668),
.B(n_483),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_572),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_575),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_582),
.B(n_370),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_673),
.B(n_485),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_582),
.B(n_370),
.Y(n_847)
);

BUFx6f_ASAP7_75t_SL g848 ( 
.A(n_682),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_673),
.B(n_485),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_674),
.B(n_488),
.Y(n_850)
);

AND2x4_ASAP7_75t_L g851 ( 
.A(n_648),
.B(n_471),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_572),
.A2(n_473),
.B(n_474),
.C(n_475),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_488),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_574),
.A2(n_362),
.B1(n_252),
.B2(n_260),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_582),
.B(n_300),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_675),
.A2(n_549),
.B(n_538),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_679),
.B(n_242),
.Y(n_857)
);

OAI22x1_ASAP7_75t_SL g858 ( 
.A1(n_679),
.A2(n_307),
.B1(n_313),
.B2(n_298),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_574),
.A2(n_300),
.B1(n_341),
.B2(n_351),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_685),
.B(n_496),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_685),
.B(n_512),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_701),
.B(n_300),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_701),
.B(n_341),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_576),
.A2(n_341),
.B1(n_351),
.B2(n_476),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_705),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_838),
.A2(n_578),
.B1(n_585),
.B2(n_592),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_709),
.B(n_706),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_764),
.B(n_687),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_766),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_713),
.B(n_701),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_767),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_774),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_706),
.B(n_687),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_R g874 ( 
.A(n_718),
.B(n_277),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_769),
.B(n_702),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_789),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_755),
.B(n_474),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_769),
.B(n_702),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_763),
.B(n_648),
.Y(n_879)
);

OR2x6_ASAP7_75t_L g880 ( 
.A(n_792),
.B(n_444),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_838),
.A2(n_578),
.B1(n_585),
.B2(n_592),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_812),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_812),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_722),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_851),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_715),
.B(n_294),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_711),
.B(n_649),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_744),
.A2(n_597),
.B(n_576),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_790),
.A2(n_691),
.B1(n_653),
.B2(n_649),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_711),
.B(n_653),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_851),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_762),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_780),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_830),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_789),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_789),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_761),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_759),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_794),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_728),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_746),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_790),
.B(n_596),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_798),
.B(n_670),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_816),
.B(n_596),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_798),
.B(n_701),
.Y(n_905)
);

O2A1O1Ixp5_ASAP7_75t_L g906 ( 
.A1(n_827),
.A2(n_600),
.B(n_575),
.C(n_577),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_828),
.A2(n_670),
.B1(n_690),
.B2(n_691),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_816),
.B(n_596),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_708),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_727),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_743),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_725),
.B(n_444),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_733),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_725),
.B(n_445),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_735),
.A2(n_597),
.B1(n_341),
.B2(n_351),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_717),
.B(n_692),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_789),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_819),
.A2(n_730),
.B1(n_731),
.B2(n_723),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_SL g919 ( 
.A(n_793),
.B(n_701),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_819),
.A2(n_692),
.B1(n_596),
.B2(n_644),
.Y(n_920)
);

BUFx4f_ASAP7_75t_L g921 ( 
.A(n_792),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_754),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_757),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_799),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_843),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_717),
.B(n_609),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_792),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_707),
.Y(n_928)
);

INVx6_ASAP7_75t_L g929 ( 
.A(n_797),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_793),
.B(n_712),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_829),
.B(n_609),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_797),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_745),
.B(n_609),
.Y(n_933)
);

AND2x6_ASAP7_75t_L g934 ( 
.A(n_736),
.B(n_604),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_714),
.B(n_609),
.Y(n_935)
);

INVx1_ASAP7_75t_SL g936 ( 
.A(n_821),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_802),
.B(n_701),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_777),
.A2(n_606),
.B(n_631),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_738),
.Y(n_939)
);

AND3x2_ASAP7_75t_SL g940 ( 
.A(n_735),
.B(n_1),
.C(n_3),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_804),
.Y(n_941)
);

BUFx4f_ASAP7_75t_L g942 ( 
.A(n_797),
.Y(n_942)
);

BUFx2_ASAP7_75t_L g943 ( 
.A(n_829),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_823),
.B(n_619),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_828),
.A2(n_703),
.B1(n_699),
.B2(n_604),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_808),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_740),
.B(n_619),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_800),
.Y(n_948)
);

INVx5_ASAP7_75t_L g949 ( 
.A(n_828),
.Y(n_949)
);

INVx4_ASAP7_75t_L g950 ( 
.A(n_808),
.Y(n_950)
);

NOR3xp33_ASAP7_75t_SL g951 ( 
.A(n_825),
.B(n_317),
.C(n_316),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_750),
.B(n_604),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_801),
.B(n_605),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_732),
.B(n_445),
.Y(n_954)
);

NOR3xp33_ASAP7_75t_SL g955 ( 
.A(n_719),
.B(n_323),
.C(n_325),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_726),
.B(n_446),
.Y(n_956)
);

A2O1A1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_787),
.A2(n_726),
.B(n_747),
.C(n_739),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_841),
.A2(n_351),
.B1(n_341),
.B2(n_601),
.Y(n_958)
);

INVx3_ASAP7_75t_L g959 ( 
.A(n_799),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_772),
.B(n_619),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_857),
.B(n_619),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_739),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_857),
.B(n_636),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_858),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_827),
.B(n_636),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_737),
.B(n_636),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_747),
.A2(n_636),
.B1(n_644),
.B2(n_684),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_817),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_758),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_748),
.B(n_605),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_770),
.B(n_446),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_741),
.B(n_644),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_859),
.A2(n_351),
.B1(n_341),
.B2(n_601),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_R g974 ( 
.A(n_742),
.B(n_331),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_820),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_806),
.B(n_613),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_770),
.A2(n_684),
.B1(n_699),
.B2(n_613),
.Y(n_977)
);

NAND3xp33_ASAP7_75t_SL g978 ( 
.A(n_787),
.B(n_338),
.C(n_333),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_SL g979 ( 
.A1(n_721),
.A2(n_340),
.B1(n_346),
.B2(n_378),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_795),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_724),
.B(n_684),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_751),
.A2(n_684),
.B1(n_699),
.B2(n_676),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_786),
.B(n_613),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_752),
.B(n_621),
.Y(n_984)
);

OR2x2_ASAP7_75t_L g985 ( 
.A(n_779),
.B(n_348),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_809),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_781),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_716),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_756),
.B(n_621),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_824),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_826),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_721),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_832),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_729),
.B(n_621),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_834),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_808),
.B(n_623),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_803),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_808),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_859),
.A2(n_351),
.B1(n_583),
.B2(n_581),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_776),
.B(n_703),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_734),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_753),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_803),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_749),
.B(n_447),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_805),
.B(n_703),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_810),
.A2(n_623),
.B(n_696),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_814),
.Y(n_1007)
);

OR2x6_ASAP7_75t_L g1008 ( 
.A(n_771),
.B(n_852),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_831),
.B(n_626),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_842),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_846),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_809),
.Y(n_1012)
);

INVx5_ASAP7_75t_L g1013 ( 
.A(n_753),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_710),
.B(n_447),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_778),
.B(n_626),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_720),
.A2(n_583),
.B1(n_577),
.B2(n_579),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_836),
.Y(n_1017)
);

INVx2_ASAP7_75t_SL g1018 ( 
.A(n_844),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_811),
.B(n_448),
.Y(n_1019)
);

NAND3xp33_ASAP7_75t_SL g1020 ( 
.A(n_833),
.B(n_361),
.C(n_352),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_753),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_854),
.B(n_657),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_854),
.B(n_626),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_849),
.B(n_627),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_788),
.B(n_657),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_782),
.B(n_627),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_848),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_850),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_753),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_853),
.B(n_627),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_860),
.B(n_671),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_861),
.B(n_671),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_784),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_785),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_815),
.B(n_671),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_760),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_SL g1037 ( 
.A1(n_753),
.A2(n_371),
.B1(n_363),
.B2(n_682),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_822),
.B(n_448),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_768),
.B(n_676),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_773),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_783),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_775),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_835),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_856),
.Y(n_1044)
);

INVxp67_ASAP7_75t_L g1045 ( 
.A(n_840),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_867),
.A2(n_791),
.B(n_835),
.C(n_845),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_867),
.A2(n_847),
.B1(n_839),
.B2(n_837),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_938),
.A2(n_765),
.B(n_680),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_910),
.Y(n_1049)
);

AOI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_1003),
.A2(n_848),
.B1(n_796),
.B2(n_661),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_1035),
.A2(n_765),
.B(n_680),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_969),
.B(n_579),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_1005),
.A2(n_680),
.B(n_631),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_901),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_873),
.B(n_581),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_899),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_SL g1057 ( 
.A1(n_979),
.A2(n_864),
.B1(n_450),
.B2(n_452),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_957),
.A2(n_864),
.B1(n_807),
.B2(n_813),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_902),
.A2(n_818),
.B(n_681),
.C(n_683),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_965),
.A2(n_602),
.B(n_606),
.Y(n_1060)
);

NAND2x2_ASAP7_75t_L g1061 ( 
.A(n_997),
.B(n_321),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_946),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_946),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_933),
.A2(n_602),
.B(n_606),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_913),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_962),
.A2(n_863),
.B(n_862),
.C(n_855),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1003),
.A2(n_681),
.B(n_696),
.C(n_676),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1028),
.B(n_584),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_962),
.B(n_681),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_961),
.A2(n_602),
.B(n_631),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1028),
.B(n_912),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_914),
.B(n_584),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_979),
.A2(n_586),
.B1(n_590),
.B2(n_599),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_874),
.B(n_686),
.C(n_454),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_897),
.B(n_697),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_873),
.B(n_586),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_992),
.A2(n_682),
.B1(n_696),
.B2(n_683),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_963),
.A2(n_631),
.B(n_680),
.Y(n_1078)
);

OR2x6_ASAP7_75t_SL g1079 ( 
.A(n_927),
.B(n_683),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_923),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_892),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_876),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_956),
.B(n_589),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_971),
.B(n_589),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_936),
.B(n_450),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_909),
.B(n_980),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_943),
.B(n_661),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_898),
.B(n_657),
.Y(n_1088)
);

INVxp33_ASAP7_75t_SL g1089 ( 
.A(n_932),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_930),
.B(n_697),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_904),
.A2(n_600),
.B(n_599),
.C(n_590),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_978),
.B(n_454),
.C(n_452),
.Y(n_1092)
);

BUFx4f_ASAP7_75t_L g1093 ( 
.A(n_929),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_876),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_990),
.B(n_697),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_904),
.A2(n_431),
.B(n_451),
.C(n_549),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_894),
.B(n_697),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1001),
.A2(n_682),
.B1(n_516),
.B2(n_538),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_894),
.A2(n_512),
.B(n_516),
.C(n_523),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_925),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_879),
.A2(n_697),
.B(n_682),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_892),
.Y(n_1102)
);

OA21x2_ASAP7_75t_L g1103 ( 
.A1(n_888),
.A2(n_492),
.B(n_476),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_960),
.A2(n_1),
.B(n_6),
.C(n_10),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_869),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_949),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1025),
.A2(n_492),
.B(n_476),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_886),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_887),
.A2(n_492),
.B(n_476),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_908),
.A2(n_14),
.B(n_22),
.C(n_25),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_L g1111 ( 
.A(n_949),
.B(n_492),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_876),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_929),
.B(n_85),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_SL g1114 ( 
.A(n_874),
.B(n_25),
.C(n_28),
.Y(n_1114)
);

BUFx2_ASAP7_75t_L g1115 ( 
.A(n_884),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_908),
.A2(n_29),
.B(n_32),
.C(n_33),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_987),
.B(n_101),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_890),
.A2(n_492),
.B(n_476),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_981),
.A2(n_492),
.B(n_98),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_SL g1120 ( 
.A1(n_988),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_872),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_926),
.A2(n_492),
.B(n_105),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_922),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1007),
.B(n_36),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_948),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_882),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_877),
.B(n_37),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_954),
.B(n_40),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_868),
.A2(n_115),
.B(n_177),
.Y(n_1129)
);

OAI21xp33_ASAP7_75t_L g1130 ( 
.A1(n_974),
.A2(n_40),
.B(n_41),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1000),
.A2(n_97),
.B(n_175),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_883),
.Y(n_1132)
);

INVxp67_ASAP7_75t_SL g1133 ( 
.A(n_876),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_SL g1134 ( 
.A1(n_974),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_SL g1135 ( 
.A1(n_964),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_991),
.B(n_124),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_949),
.A2(n_49),
.B1(n_50),
.B2(n_54),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_916),
.A2(n_129),
.B(n_174),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_960),
.B(n_55),
.Y(n_1139)
);

INVx3_ASAP7_75t_L g1140 ( 
.A(n_950),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_931),
.A2(n_55),
.B(n_56),
.C(n_58),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_949),
.A2(n_881),
.B1(n_866),
.B2(n_1010),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_968),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_921),
.Y(n_1144)
);

AND2x2_ASAP7_75t_SL g1145 ( 
.A(n_921),
.B(n_58),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_928),
.B(n_941),
.Y(n_1146)
);

AND2x4_ASAP7_75t_SL g1147 ( 
.A(n_880),
.B(n_142),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1006),
.A2(n_131),
.B(n_173),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_895),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1004),
.B(n_61),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_880),
.B(n_61),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_L g1153 ( 
.A(n_985),
.B(n_63),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_935),
.A2(n_151),
.B(n_75),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_895),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_885),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_902),
.A2(n_154),
.B(n_77),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_866),
.A2(n_65),
.B1(n_80),
.B2(n_121),
.Y(n_1158)
);

XOR2xp5_ASAP7_75t_L g1159 ( 
.A(n_1027),
.B(n_125),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_895),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_993),
.B(n_995),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_929),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_1045),
.A2(n_156),
.B1(n_160),
.B2(n_166),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1009),
.A2(n_168),
.B(n_190),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_891),
.Y(n_1165)
);

O2A1O1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_931),
.A2(n_875),
.B(n_878),
.C(n_903),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_880),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_1045),
.B(n_1020),
.C(n_1011),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_955),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_953),
.B(n_976),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_939),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1031),
.A2(n_1032),
.B(n_919),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_953),
.Y(n_1173)
);

OAI22xp33_ASAP7_75t_SL g1174 ( 
.A1(n_940),
.A2(n_1008),
.B1(n_1022),
.B2(n_1041),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1008),
.A2(n_983),
.B1(n_994),
.B2(n_900),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_976),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1013),
.A2(n_1019),
.B(n_1038),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1013),
.A2(n_1030),
.B(n_1024),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1013),
.A2(n_1030),
.B(n_1024),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_900),
.B(n_911),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_865),
.B(n_871),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_911),
.B(n_1036),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1040),
.B(n_1042),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_893),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_970),
.A2(n_984),
.B(n_989),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1017),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_L g1188 ( 
.A1(n_966),
.A2(n_972),
.B(n_944),
.C(n_1023),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1018),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_895),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_942),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_865),
.B(n_918),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_896),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1039),
.B(n_1015),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_951),
.A2(n_1008),
.B(n_955),
.C(n_952),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1039),
.B(n_1015),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_942),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_947),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_924),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_896),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1188),
.A2(n_944),
.B(n_966),
.C(n_972),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1162),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1071),
.B(n_905),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1056),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1178),
.A2(n_1013),
.B(n_907),
.Y(n_1205)
);

AOI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1153),
.A2(n_983),
.B(n_994),
.Y(n_1206)
);

INVx4_ASAP7_75t_L g1207 ( 
.A(n_1093),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_SL g1208 ( 
.A1(n_1106),
.A2(n_952),
.B(n_1026),
.C(n_984),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1067),
.A2(n_945),
.A3(n_1043),
.B(n_1044),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1054),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1161),
.B(n_881),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1127),
.B(n_1014),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_SL g1213 ( 
.A1(n_1124),
.A2(n_1134),
.B(n_1130),
.Y(n_1213)
);

OAI22x1_ASAP7_75t_L g1214 ( 
.A1(n_1169),
.A2(n_940),
.B1(n_905),
.B2(n_977),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1123),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1086),
.B(n_1146),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1128),
.B(n_1014),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1172),
.A2(n_1179),
.B(n_1059),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1051),
.A2(n_906),
.B(n_970),
.Y(n_1220)
);

AOI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1177),
.A2(n_1055),
.B(n_1192),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1161),
.B(n_1180),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1182),
.B(n_958),
.Y(n_1223)
);

NAND2x1p5_ASAP7_75t_L g1224 ( 
.A(n_1150),
.B(n_950),
.Y(n_1224)
);

AO21x2_ASAP7_75t_L g1225 ( 
.A1(n_1046),
.A2(n_1148),
.B(n_1055),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1115),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1142),
.A2(n_1026),
.B(n_996),
.Y(n_1227)
);

AO32x2_ASAP7_75t_L g1228 ( 
.A1(n_1142),
.A2(n_1158),
.A3(n_1058),
.B1(n_1073),
.B2(n_1057),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1076),
.A2(n_1196),
.B(n_1194),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1089),
.B(n_1029),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_1174),
.A2(n_996),
.B(n_967),
.Y(n_1231)
);

CKINVDCx9p33_ASAP7_75t_R g1232 ( 
.A(n_1087),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1070),
.A2(n_1078),
.B(n_1060),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1194),
.A2(n_920),
.B(n_889),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1100),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1064),
.A2(n_982),
.B(n_1016),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1146),
.B(n_1197),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1183),
.B(n_958),
.Y(n_1238)
);

OAI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1175),
.A2(n_1037),
.B1(n_1021),
.B2(n_1002),
.Y(n_1239)
);

OA21x2_ASAP7_75t_L g1240 ( 
.A1(n_1091),
.A2(n_973),
.B(n_915),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_1058),
.A2(n_870),
.B(n_937),
.C(n_986),
.Y(n_1241)
);

OR2x2_ASAP7_75t_L g1242 ( 
.A(n_1085),
.B(n_1012),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1186),
.B(n_1151),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1166),
.A2(n_1037),
.B(n_915),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1196),
.A2(n_896),
.B(n_917),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1081),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1105),
.Y(n_1247)
);

INVx5_ASAP7_75t_L g1248 ( 
.A(n_1200),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1168),
.A2(n_1012),
.B1(n_924),
.B2(n_959),
.Y(n_1249)
);

AOI221xp5_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_973),
.B1(n_1016),
.B2(n_999),
.C(n_1021),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1047),
.A2(n_999),
.B(n_934),
.Y(n_1251)
);

NOR2xp67_ASAP7_75t_L g1252 ( 
.A(n_1108),
.B(n_986),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1053),
.A2(n_959),
.B(n_934),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1107),
.A2(n_934),
.B(n_1002),
.Y(n_1254)
);

O2A1O1Ixp5_ASAP7_75t_SL g1255 ( 
.A1(n_1106),
.A2(n_1014),
.B(n_934),
.C(n_917),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1176),
.B(n_1002),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1186),
.B(n_1173),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1170),
.A2(n_1021),
.B1(n_917),
.B2(n_998),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1072),
.B(n_1021),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1083),
.A2(n_998),
.B(n_1084),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1121),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1101),
.A2(n_998),
.B(n_1073),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1102),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_1093),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1184),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1068),
.B(n_998),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1096),
.A2(n_1090),
.A3(n_1158),
.B(n_1110),
.Y(n_1267)
);

INVx5_ASAP7_75t_L g1268 ( 
.A(n_1094),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1170),
.B(n_1139),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1136),
.A2(n_1052),
.B(n_1095),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1198),
.B(n_1171),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1109),
.A2(n_1118),
.B(n_1052),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1136),
.A2(n_1095),
.B(n_1097),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1103),
.A2(n_1181),
.B(n_1131),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1122),
.A2(n_1119),
.B(n_1138),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1195),
.A2(n_1157),
.B(n_1129),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1103),
.A2(n_1164),
.B(n_1154),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1102),
.B(n_1132),
.Y(n_1279)
);

OAI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1066),
.A2(n_1069),
.B(n_1050),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1111),
.A2(n_1150),
.B(n_1190),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1150),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1150),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1187),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1049),
.A2(n_1125),
.B(n_1143),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_L g1286 ( 
.A1(n_1156),
.A2(n_1165),
.B(n_1104),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1065),
.Y(n_1287)
);

NOR2x1_ASAP7_75t_L g1288 ( 
.A(n_1082),
.B(n_1140),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1152),
.B(n_1145),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1190),
.A2(n_1075),
.B(n_1077),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1088),
.B(n_1117),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1116),
.A2(n_1141),
.B(n_1137),
.C(n_1092),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1117),
.B(n_1189),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1190),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1080),
.B(n_1149),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1191),
.A2(n_1144),
.B1(n_1167),
.B2(n_1113),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1199),
.B(n_1074),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1190),
.A2(n_1098),
.B1(n_1133),
.B2(n_1063),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1137),
.A2(n_1082),
.A3(n_1099),
.B(n_1114),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1062),
.A2(n_1140),
.B(n_1063),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1094),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1079),
.B(n_1062),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1113),
.A2(n_1061),
.B(n_1163),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1094),
.Y(n_1304)
);

AOI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1113),
.A2(n_1159),
.B(n_1112),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1147),
.B(n_1112),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1112),
.A2(n_1155),
.B(n_1160),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1155),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1135),
.B(n_1160),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1160),
.A2(n_1193),
.B(n_1200),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1193),
.Y(n_1311)
);

OR2x6_ASAP7_75t_L g1312 ( 
.A(n_1193),
.B(n_1162),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1127),
.B(n_867),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1102),
.Y(n_1315)
);

O2A1O1Ixp5_ASAP7_75t_L g1316 ( 
.A1(n_1188),
.A2(n_957),
.B(n_1179),
.C(n_1178),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1071),
.B(n_867),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1188),
.A2(n_867),
.B(n_957),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1130),
.A2(n_867),
.B1(n_838),
.B2(n_979),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1071),
.B(n_867),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1056),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1071),
.B(n_867),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1056),
.Y(n_1325)
);

NAND2xp33_ASAP7_75t_L g1326 ( 
.A(n_1142),
.B(n_949),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1056),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1062),
.Y(n_1328)
);

AO21x2_ASAP7_75t_L g1329 ( 
.A1(n_1178),
.A2(n_1179),
.B(n_957),
.Y(n_1329)
);

BUFx4_ASAP7_75t_SL g1330 ( 
.A(n_1144),
.Y(n_1330)
);

INVxp67_ASAP7_75t_SL g1331 ( 
.A(n_1142),
.Y(n_1331)
);

OAI22x1_ASAP7_75t_L g1332 ( 
.A1(n_1153),
.A2(n_867),
.B1(n_558),
.B2(n_709),
.Y(n_1332)
);

AOI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1178),
.A2(n_1179),
.B(n_1172),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1123),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1067),
.A2(n_1046),
.A3(n_957),
.B(n_1058),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1336)
);

O2A1O1Ixp5_ASAP7_75t_L g1337 ( 
.A1(n_1188),
.A2(n_957),
.B(n_1179),
.C(n_1178),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1056),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1056),
.Y(n_1340)
);

A2O1A1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1153),
.A2(n_867),
.B(n_709),
.C(n_957),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1056),
.Y(n_1343)
);

AOI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1153),
.A2(n_867),
.B1(n_709),
.B2(n_790),
.Y(n_1344)
);

INVx5_ASAP7_75t_SL g1345 ( 
.A(n_1113),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1071),
.B(n_867),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1071),
.B(n_867),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1178),
.A2(n_1179),
.B(n_1177),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1056),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1188),
.A2(n_867),
.B(n_957),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1048),
.A2(n_1185),
.B(n_906),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1127),
.B(n_867),
.Y(n_1353)
);

BUFx6f_ASAP7_75t_L g1354 ( 
.A(n_1150),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1071),
.B(n_616),
.Y(n_1355)
);

CKINVDCx11_ASAP7_75t_R g1356 ( 
.A(n_1079),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1071),
.B(n_867),
.Y(n_1357)
);

NAND2x1p5_ASAP7_75t_L g1358 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1358)
);

INVxp67_ASAP7_75t_SL g1359 ( 
.A(n_1279),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1344),
.A2(n_1341),
.B(n_1244),
.C(n_1250),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1204),
.Y(n_1361)
);

NAND2x1p5_ASAP7_75t_L g1362 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1362)
);

INVx8_ASAP7_75t_L g1363 ( 
.A(n_1248),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1305),
.B(n_1292),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1205),
.A2(n_1221),
.B(n_1274),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1264),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1253),
.A2(n_1273),
.B(n_1233),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1314),
.B(n_1353),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1332),
.A2(n_1341),
.B1(n_1319),
.B2(n_1213),
.C(n_1292),
.Y(n_1369)
);

OAI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1319),
.A2(n_1222),
.B1(n_1357),
.B2(n_1320),
.Y(n_1370)
);

OR2x6_ASAP7_75t_L g1371 ( 
.A(n_1251),
.B(n_1303),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1316),
.A2(n_1337),
.B(n_1323),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1247),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1317),
.B(n_1324),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1327),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1215),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1215),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1349),
.A2(n_1274),
.A3(n_1205),
.B(n_1227),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_SL g1379 ( 
.A1(n_1250),
.A2(n_1206),
.B(n_1211),
.C(n_1286),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1340),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1349),
.A2(n_1326),
.B(n_1271),
.Y(n_1381)
);

AO21x1_ASAP7_75t_L g1382 ( 
.A1(n_1326),
.A2(n_1280),
.B(n_1203),
.Y(n_1382)
);

OA21x2_ASAP7_75t_L g1383 ( 
.A1(n_1316),
.A2(n_1338),
.B(n_1352),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1347),
.A2(n_1348),
.B1(n_1331),
.B2(n_1203),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1315),
.Y(n_1385)
);

OAI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1291),
.A2(n_1345),
.B1(n_1355),
.B2(n_1243),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1322),
.A2(n_1346),
.B(n_1342),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1235),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1210),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1257),
.B(n_1272),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_1210),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1261),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1336),
.A2(n_1201),
.B(n_1220),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1265),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1321),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1263),
.B(n_1270),
.Y(n_1396)
);

A2O1A1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1331),
.A2(n_1229),
.B(n_1201),
.C(n_1227),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1226),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1283),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1271),
.A2(n_1236),
.B(n_1278),
.Y(n_1400)
);

AOI22x1_ASAP7_75t_L g1401 ( 
.A1(n_1214),
.A2(n_1277),
.B1(n_1275),
.B2(n_1290),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_1334),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1234),
.A2(n_1241),
.B(n_1260),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1256),
.B(n_1306),
.Y(n_1404)
);

AO21x2_ASAP7_75t_L g1405 ( 
.A1(n_1333),
.A2(n_1275),
.B(n_1225),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1217),
.B(n_1223),
.Y(n_1406)
);

NOR2xp67_ASAP7_75t_L g1407 ( 
.A(n_1207),
.B(n_1293),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1345),
.A2(n_1296),
.B1(n_1252),
.B2(n_1242),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1245),
.A2(n_1254),
.B(n_1260),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1289),
.B(n_1246),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1325),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1218),
.B(n_1212),
.C(n_1309),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1226),
.Y(n_1413)
);

AOI22x1_ASAP7_75t_L g1414 ( 
.A1(n_1290),
.A2(n_1350),
.B1(n_1343),
.B2(n_1339),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1241),
.A2(n_1234),
.B(n_1208),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1217),
.B(n_1237),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1309),
.A2(n_1356),
.B1(n_1238),
.B2(n_1225),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1356),
.A2(n_1269),
.B1(n_1284),
.B2(n_1287),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1259),
.A2(n_1266),
.B(n_1285),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1295),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1202),
.Y(n_1421)
);

AOI22x1_ASAP7_75t_L g1422 ( 
.A1(n_1207),
.A2(n_1281),
.B1(n_1328),
.B2(n_1294),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1219),
.A2(n_1255),
.B(n_1276),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1209),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1330),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_SL g1426 ( 
.A1(n_1281),
.A2(n_1239),
.B(n_1307),
.Y(n_1426)
);

INVx8_ASAP7_75t_L g1427 ( 
.A(n_1248),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1301),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1230),
.B(n_1302),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1297),
.A2(n_1249),
.B(n_1298),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1330),
.Y(n_1431)
);

BUFx3_ASAP7_75t_L g1432 ( 
.A(n_1311),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1302),
.A2(n_1329),
.B1(n_1228),
.B2(n_1258),
.C(n_1308),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1304),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1312),
.Y(n_1435)
);

CKINVDCx20_ASAP7_75t_R g1436 ( 
.A(n_1232),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1209),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_1312),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_SL g1439 ( 
.A(n_1283),
.B(n_1354),
.Y(n_1439)
);

AO21x2_ASAP7_75t_L g1440 ( 
.A1(n_1329),
.A2(n_1307),
.B(n_1300),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1312),
.A2(n_1328),
.B1(n_1294),
.B2(n_1268),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1248),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1219),
.A2(n_1276),
.B(n_1240),
.Y(n_1443)
);

OAI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1228),
.A2(n_1240),
.B1(n_1354),
.B2(n_1268),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1219),
.A2(n_1276),
.B(n_1240),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1228),
.A2(n_1335),
.B(n_1267),
.C(n_1288),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1224),
.A2(n_1310),
.B(n_1335),
.Y(n_1447)
);

AO31x2_ASAP7_75t_L g1448 ( 
.A1(n_1228),
.A2(n_1267),
.A3(n_1209),
.B(n_1299),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1268),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1224),
.A2(n_1209),
.B(n_1267),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_L g1451 ( 
.A1(n_1267),
.A2(n_1232),
.B(n_1299),
.Y(n_1451)
);

NAND3xp33_ASAP7_75t_SL g1452 ( 
.A(n_1299),
.B(n_1344),
.C(n_867),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1299),
.A2(n_867),
.B(n_1341),
.C(n_957),
.Y(n_1453)
);

INVx3_ASAP7_75t_SL g1454 ( 
.A(n_1354),
.Y(n_1454)
);

AOI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1205),
.A2(n_1179),
.B(n_1178),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1282),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1314),
.B(n_1353),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_SL g1458 ( 
.A(n_1344),
.B(n_1341),
.Y(n_1458)
);

O2A1O1Ixp33_ASAP7_75t_L g1459 ( 
.A1(n_1341),
.A2(n_867),
.B(n_957),
.C(n_709),
.Y(n_1459)
);

NOR2xp67_ASAP7_75t_R g1460 ( 
.A(n_1207),
.B(n_1162),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1204),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1317),
.B(n_867),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1344),
.A2(n_867),
.B1(n_1319),
.B2(n_1341),
.Y(n_1464)
);

INVx5_ASAP7_75t_L g1465 ( 
.A(n_1282),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1332),
.A2(n_867),
.B1(n_1344),
.B2(n_1319),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1204),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1282),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1204),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1204),
.Y(n_1474)
);

NAND2x1p5_ASAP7_75t_L g1475 ( 
.A(n_1282),
.B(n_1283),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1207),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1349),
.A2(n_1351),
.B(n_1318),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1344),
.B(n_867),
.C(n_790),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1215),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1344),
.A2(n_867),
.B(n_957),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1349),
.A2(n_1351),
.B(n_1318),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1317),
.B(n_867),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1226),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1205),
.A2(n_1179),
.B(n_1178),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1215),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1244),
.A2(n_1179),
.B(n_1178),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1355),
.B(n_1317),
.Y(n_1487)
);

AOI211xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1344),
.A2(n_867),
.B(n_1341),
.C(n_1174),
.Y(n_1488)
);

BUFx8_ASAP7_75t_SL g1489 ( 
.A(n_1215),
.Y(n_1489)
);

NAND3xp33_ASAP7_75t_SL g1490 ( 
.A(n_1344),
.B(n_867),
.C(n_709),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1204),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1332),
.A2(n_867),
.B1(n_1344),
.B2(n_1319),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1256),
.B(n_1170),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1244),
.A2(n_1179),
.B(n_1178),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1262),
.A2(n_1313),
.B(n_1216),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1349),
.A2(n_1351),
.B(n_1318),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_SL g1498 ( 
.A1(n_1303),
.A2(n_1231),
.B(n_1292),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1332),
.A2(n_867),
.B1(n_1344),
.B2(n_1319),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1204),
.Y(n_1500)
);

BUFx3_ASAP7_75t_L g1501 ( 
.A(n_1366),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1359),
.B(n_1374),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1360),
.A2(n_1467),
.B1(n_1499),
.B2(n_1493),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1368),
.B(n_1457),
.Y(n_1504)
);

AND2x4_ASAP7_75t_SL g1505 ( 
.A(n_1376),
.B(n_1479),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_SL g1506 ( 
.A(n_1364),
.B(n_1371),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_1489),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1396),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1384),
.B(n_1370),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1366),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1360),
.A2(n_1499),
.B1(n_1493),
.B2(n_1467),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1406),
.B(n_1410),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1404),
.B(n_1410),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1478),
.A2(n_1464),
.B1(n_1480),
.B2(n_1482),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_1490),
.A2(n_1459),
.B(n_1458),
.C(n_1452),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1463),
.B(n_1390),
.Y(n_1516)
);

O2A1O1Ixp33_ASAP7_75t_L g1517 ( 
.A1(n_1458),
.A2(n_1453),
.B(n_1379),
.C(n_1488),
.Y(n_1517)
);

CKINVDCx16_ASAP7_75t_R g1518 ( 
.A(n_1376),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1434),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1384),
.A2(n_1369),
.B1(n_1444),
.B2(n_1436),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1442),
.A2(n_1386),
.B(n_1397),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1494),
.B(n_1416),
.Y(n_1522)
);

O2A1O1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1379),
.A2(n_1397),
.B(n_1498),
.C(n_1408),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1442),
.A2(n_1364),
.B(n_1381),
.Y(n_1524)
);

OA22x2_ASAP7_75t_L g1525 ( 
.A1(n_1364),
.A2(n_1371),
.B1(n_1430),
.B2(n_1394),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1486),
.A2(n_1495),
.B(n_1497),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1420),
.B(n_1385),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1417),
.B(n_1433),
.Y(n_1528)
);

INVx3_ASAP7_75t_SL g1529 ( 
.A(n_1402),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1412),
.B(n_1417),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1429),
.A2(n_1403),
.B(n_1407),
.C(n_1418),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1429),
.B(n_1436),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1446),
.A2(n_1432),
.B(n_1441),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1388),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1415),
.A2(n_1423),
.B(n_1443),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_1489),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1444),
.A2(n_1446),
.B1(n_1395),
.B2(n_1411),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1392),
.A2(n_1413),
.B1(n_1361),
.B2(n_1491),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1371),
.A2(n_1426),
.B(n_1439),
.C(n_1373),
.Y(n_1539)
);

O2A1O1Ixp33_ASAP7_75t_L g1540 ( 
.A1(n_1439),
.A2(n_1500),
.B(n_1380),
.C(n_1461),
.Y(n_1540)
);

BUFx6f_ASAP7_75t_L g1541 ( 
.A(n_1363),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1398),
.B(n_1483),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1476),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1358),
.A2(n_1475),
.B(n_1362),
.Y(n_1544)
);

AOI221xp5_ASAP7_75t_L g1545 ( 
.A1(n_1477),
.A2(n_1481),
.B1(n_1375),
.B2(n_1469),
.C(n_1474),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1473),
.A2(n_1425),
.B(n_1428),
.C(n_1431),
.Y(n_1546)
);

BUFx12f_ASAP7_75t_L g1547 ( 
.A(n_1377),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1358),
.A2(n_1362),
.B(n_1475),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_SL g1549 ( 
.A1(n_1449),
.A2(n_1419),
.B(n_1402),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1419),
.B(n_1448),
.Y(n_1550)
);

O2A1O1Ixp5_ASAP7_75t_L g1551 ( 
.A1(n_1365),
.A2(n_1484),
.B(n_1455),
.C(n_1437),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1413),
.A2(n_1479),
.B1(n_1389),
.B2(n_1465),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1419),
.A2(n_1427),
.B(n_1363),
.Y(n_1553)
);

AOI21x1_ASAP7_75t_SL g1554 ( 
.A1(n_1460),
.A2(n_1401),
.B(n_1422),
.Y(n_1554)
);

O2A1O1Ixp33_ASAP7_75t_L g1555 ( 
.A1(n_1454),
.A2(n_1456),
.B(n_1472),
.C(n_1399),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1415),
.A2(n_1423),
.B(n_1443),
.Y(n_1556)
);

O2A1O1Ixp5_ASAP7_75t_L g1557 ( 
.A1(n_1424),
.A2(n_1437),
.B(n_1414),
.C(n_1451),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1389),
.A2(n_1465),
.B1(n_1391),
.B2(n_1421),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1405),
.A2(n_1400),
.B(n_1447),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1424),
.A2(n_1421),
.B(n_1440),
.C(n_1405),
.Y(n_1560)
);

AOI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1400),
.A2(n_1447),
.B(n_1440),
.Y(n_1561)
);

O2A1O1Ixp5_ASAP7_75t_L g1562 ( 
.A1(n_1451),
.A2(n_1378),
.B(n_1450),
.C(n_1409),
.Y(n_1562)
);

AOI21x1_ASAP7_75t_SL g1563 ( 
.A1(n_1427),
.A2(n_1465),
.B(n_1476),
.Y(n_1563)
);

AOI221x1_ASAP7_75t_SL g1564 ( 
.A1(n_1448),
.A2(n_1485),
.B1(n_1377),
.B2(n_1378),
.C(n_1476),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1372),
.A2(n_1400),
.B1(n_1393),
.B2(n_1383),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1372),
.B(n_1383),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1383),
.B(n_1445),
.Y(n_1567)
);

INVx5_ASAP7_75t_L g1568 ( 
.A(n_1387),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1445),
.B(n_1393),
.Y(n_1569)
);

A2O1A1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1367),
.A2(n_1468),
.B(n_1492),
.C(n_1462),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1393),
.A2(n_1470),
.B1(n_1462),
.B2(n_1466),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1468),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1470),
.B(n_1471),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1471),
.A2(n_1492),
.B(n_1496),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1496),
.Y(n_1575)
);

AND2x4_ASAP7_75t_L g1576 ( 
.A(n_1435),
.B(n_1438),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1364),
.B(n_1371),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1478),
.A2(n_867),
.B(n_1344),
.C(n_1341),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1487),
.B(n_1396),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1384),
.B(n_1370),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1459),
.A2(n_1341),
.B(n_867),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1487),
.B(n_1396),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1363),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1459),
.A2(n_1341),
.B(n_867),
.Y(n_1584)
);

AOI21x1_ASAP7_75t_SL g1585 ( 
.A1(n_1463),
.A2(n_1482),
.B(n_1320),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1459),
.A2(n_1341),
.B(n_867),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1384),
.B(n_1370),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1368),
.B(n_1457),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1381),
.A2(n_957),
.B(n_1480),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1381),
.A2(n_957),
.B(n_1480),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1384),
.B(n_1370),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1489),
.Y(n_1592)
);

AOI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1381),
.A2(n_957),
.B(n_1480),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1360),
.A2(n_867),
.B1(n_1344),
.B2(n_1319),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1490),
.A2(n_867),
.B(n_1341),
.C(n_957),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1384),
.B(n_1370),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1487),
.B(n_1396),
.Y(n_1597)
);

O2A1O1Ixp5_ASAP7_75t_L g1598 ( 
.A1(n_1488),
.A2(n_957),
.B(n_1458),
.C(n_1382),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1381),
.A2(n_957),
.B(n_1480),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1368),
.B(n_1457),
.Y(n_1600)
);

INVx1_ASAP7_75t_SL g1601 ( 
.A(n_1396),
.Y(n_1601)
);

CKINVDCx20_ASAP7_75t_R g1602 ( 
.A(n_1489),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1569),
.Y(n_1603)
);

NOR2x1_ASAP7_75t_SL g1604 ( 
.A(n_1577),
.B(n_1537),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1594),
.B(n_1514),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_SL g1606 ( 
.A1(n_1594),
.A2(n_1578),
.B(n_1595),
.Y(n_1606)
);

OR2x6_ASAP7_75t_L g1607 ( 
.A(n_1524),
.B(n_1589),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1550),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1502),
.B(n_1509),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1566),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1550),
.B(n_1567),
.Y(n_1611)
);

AO21x2_ASAP7_75t_L g1612 ( 
.A1(n_1526),
.A2(n_1559),
.B(n_1561),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1535),
.Y(n_1613)
);

NAND2xp33_ASAP7_75t_R g1614 ( 
.A(n_1530),
.B(n_1577),
.Y(n_1614)
);

AO21x2_ASAP7_75t_L g1615 ( 
.A1(n_1590),
.A2(n_1599),
.B(n_1593),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1519),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1537),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1556),
.B(n_1525),
.Y(n_1618)
);

AOI221xp5_ASAP7_75t_L g1619 ( 
.A1(n_1503),
.A2(n_1511),
.B1(n_1514),
.B2(n_1517),
.C(n_1598),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1572),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1575),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1515),
.A2(n_1581),
.B(n_1586),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1568),
.Y(n_1623)
);

AOI222xp33_ASAP7_75t_L g1624 ( 
.A1(n_1503),
.A2(n_1511),
.B1(n_1520),
.B2(n_1596),
.C1(n_1580),
.C2(n_1587),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1562),
.B(n_1506),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1545),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1568),
.B(n_1570),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1573),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1565),
.B(n_1551),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1601),
.B(n_1528),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1571),
.A2(n_1574),
.B(n_1554),
.Y(n_1632)
);

AO21x2_ASAP7_75t_L g1633 ( 
.A1(n_1528),
.A2(n_1591),
.B(n_1580),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1539),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1591),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1540),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1560),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1564),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1564),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1521),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1538),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1549),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1523),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1538),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1553),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1508),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1579),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1584),
.B(n_1513),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1582),
.B(n_1597),
.Y(n_1649)
);

AO21x2_ASAP7_75t_L g1650 ( 
.A1(n_1531),
.A2(n_1520),
.B(n_1533),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1516),
.A2(n_1558),
.B1(n_1532),
.B2(n_1552),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1546),
.A2(n_1555),
.B(n_1527),
.Y(n_1652)
);

BUFx4f_ASAP7_75t_SL g1653 ( 
.A(n_1507),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1637),
.B(n_1558),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1620),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1633),
.B(n_1512),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1633),
.B(n_1635),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1611),
.B(n_1588),
.Y(n_1658)
);

INVxp67_ASAP7_75t_SL g1659 ( 
.A(n_1608),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1611),
.B(n_1504),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1621),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1600),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1610),
.B(n_1542),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1613),
.Y(n_1664)
);

NOR4xp25_ASAP7_75t_SL g1665 ( 
.A(n_1614),
.B(n_1592),
.C(n_1563),
.D(n_1585),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1607),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1633),
.B(n_1576),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1603),
.B(n_1518),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1613),
.Y(n_1669)
);

OAI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1619),
.A2(n_1605),
.B1(n_1622),
.B2(n_1617),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1629),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1619),
.A2(n_1547),
.B1(n_1505),
.B2(n_1522),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1623),
.B(n_1627),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1633),
.B(n_1501),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_L g1675 ( 
.A(n_1622),
.B(n_1510),
.C(n_1548),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1623),
.B(n_1583),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1605),
.A2(n_1602),
.B1(n_1536),
.B2(n_1529),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1618),
.B(n_1628),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1670),
.A2(n_1606),
.B1(n_1651),
.B2(n_1617),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1664),
.Y(n_1680)
);

OAI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1670),
.A2(n_1607),
.B1(n_1640),
.B2(n_1641),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1675),
.A2(n_1650),
.B1(n_1640),
.B2(n_1604),
.Y(n_1682)
);

OAI211xp5_ASAP7_75t_L g1683 ( 
.A1(n_1654),
.A2(n_1624),
.B(n_1626),
.C(n_1652),
.Y(n_1683)
);

OR2x2_ASAP7_75t_L g1684 ( 
.A(n_1678),
.B(n_1646),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1668),
.Y(n_1687)
);

NAND3xp33_ASAP7_75t_L g1688 ( 
.A(n_1654),
.B(n_1624),
.C(n_1626),
.Y(n_1688)
);

OAI21xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1659),
.A2(n_1640),
.B(n_1607),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1655),
.Y(n_1690)
);

AOI222xp33_ASAP7_75t_L g1691 ( 
.A1(n_1677),
.A2(n_1641),
.B1(n_1643),
.B2(n_1639),
.C1(n_1638),
.C2(n_1644),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1666),
.B(n_1607),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1673),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1678),
.B(n_1618),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1672),
.A2(n_1651),
.B1(n_1607),
.B2(n_1609),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1668),
.Y(n_1696)
);

INVxp67_ASAP7_75t_L g1697 ( 
.A(n_1668),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1675),
.A2(n_1652),
.B1(n_1607),
.B2(n_1642),
.C(n_1631),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1673),
.B(n_1627),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1666),
.A2(n_1650),
.B1(n_1615),
.B2(n_1633),
.Y(n_1700)
);

OAI31xp33_ASAP7_75t_L g1701 ( 
.A1(n_1677),
.A2(n_1634),
.A3(n_1636),
.B(n_1650),
.Y(n_1701)
);

AOI21xp33_ASAP7_75t_L g1702 ( 
.A1(n_1674),
.A2(n_1650),
.B(n_1615),
.Y(n_1702)
);

OAI211xp5_ASAP7_75t_L g1703 ( 
.A1(n_1674),
.A2(n_1634),
.B(n_1631),
.C(n_1616),
.Y(n_1703)
);

OA21x2_ASAP7_75t_L g1704 ( 
.A1(n_1657),
.A2(n_1632),
.B(n_1630),
.Y(n_1704)
);

NAND3xp33_ASAP7_75t_L g1705 ( 
.A(n_1656),
.B(n_1636),
.C(n_1630),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1608),
.Y(n_1706)
);

AO21x2_ASAP7_75t_L g1707 ( 
.A1(n_1669),
.A2(n_1612),
.B(n_1625),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1666),
.Y(n_1708)
);

INVx1_ASAP7_75t_SL g1709 ( 
.A(n_1663),
.Y(n_1709)
);

NOR2xp33_ASAP7_75t_R g1710 ( 
.A(n_1663),
.B(n_1653),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1676),
.Y(n_1711)
);

NAND4xp25_ASAP7_75t_SL g1712 ( 
.A(n_1667),
.B(n_1642),
.C(n_1645),
.D(n_1648),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1665),
.A2(n_1635),
.B1(n_1647),
.B2(n_1649),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1685),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1688),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1685),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1692),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1692),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1686),
.Y(n_1719)
);

INVx3_ASAP7_75t_L g1720 ( 
.A(n_1699),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1680),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1690),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1687),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1709),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1683),
.B(n_1649),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1692),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_SL g1727 ( 
.A(n_1688),
.B(n_1665),
.C(n_1650),
.Y(n_1727)
);

INVx4_ASAP7_75t_SL g1728 ( 
.A(n_1692),
.Y(n_1728)
);

NOR2x1p5_ASAP7_75t_L g1729 ( 
.A(n_1687),
.B(n_1666),
.Y(n_1729)
);

OR2x6_ASAP7_75t_L g1730 ( 
.A(n_1692),
.B(n_1666),
.Y(n_1730)
);

INVx5_ASAP7_75t_L g1731 ( 
.A(n_1708),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1705),
.B(n_1706),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1707),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1706),
.B(n_1659),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1705),
.B(n_1671),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1701),
.B(n_1666),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1707),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1707),
.Y(n_1738)
);

OA21x2_ASAP7_75t_L g1739 ( 
.A1(n_1702),
.A2(n_1628),
.B(n_1661),
.Y(n_1739)
);

INVx3_ASAP7_75t_R g1740 ( 
.A(n_1735),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1714),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1714),
.Y(n_1742)
);

NAND4xp75_ASAP7_75t_L g1743 ( 
.A(n_1736),
.B(n_1701),
.C(n_1689),
.D(n_1704),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1724),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1729),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1732),
.B(n_1684),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1715),
.A2(n_1679),
.B(n_1682),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1723),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1699),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1728),
.B(n_1699),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1725),
.B(n_1696),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1728),
.B(n_1699),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1731),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1714),
.Y(n_1754)
);

INVx1_ASAP7_75t_SL g1755 ( 
.A(n_1723),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1725),
.B(n_1697),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1716),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1715),
.B(n_1658),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1717),
.Y(n_1759)
);

OR2x2_ASAP7_75t_L g1760 ( 
.A(n_1732),
.B(n_1684),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1728),
.B(n_1693),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1728),
.B(n_1693),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1728),
.B(n_1693),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1724),
.B(n_1658),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1736),
.B(n_1658),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1716),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1716),
.Y(n_1767)
);

NOR2xp33_ASAP7_75t_L g1768 ( 
.A(n_1718),
.B(n_1653),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1717),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1719),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1728),
.B(n_1708),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1727),
.A2(n_1700),
.B1(n_1698),
.B2(n_1689),
.C(n_1695),
.Y(n_1772)
);

NAND4xp25_ASAP7_75t_L g1773 ( 
.A(n_1727),
.B(n_1691),
.C(n_1717),
.D(n_1726),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1734),
.B(n_1660),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1720),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1734),
.B(n_1703),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1731),
.B(n_1710),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1719),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1721),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1734),
.B(n_1660),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1720),
.B(n_1711),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1721),
.Y(n_1782)
);

INVx3_ASAP7_75t_L g1783 ( 
.A(n_1718),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1719),
.Y(n_1784)
);

AOI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1718),
.A2(n_1615),
.B(n_1681),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1755),
.B(n_1660),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1748),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1741),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1759),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1747),
.B(n_1758),
.Y(n_1790)
);

INVxp33_ASAP7_75t_L g1791 ( 
.A(n_1777),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1750),
.B(n_1717),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1741),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1771),
.Y(n_1794)
);

OAI21xp33_ASAP7_75t_L g1795 ( 
.A1(n_1773),
.A2(n_1726),
.B(n_1712),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1742),
.Y(n_1796)
);

OAI211xp5_ASAP7_75t_L g1797 ( 
.A1(n_1772),
.A2(n_1718),
.B(n_1739),
.C(n_1726),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1779),
.Y(n_1798)
);

INVxp67_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1751),
.B(n_1663),
.Y(n_1800)
);

OR2x6_ASAP7_75t_L g1801 ( 
.A(n_1753),
.B(n_1743),
.Y(n_1801)
);

INVx1_ASAP7_75t_SL g1802 ( 
.A(n_1769),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1742),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1746),
.B(n_1735),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1754),
.Y(n_1805)
);

INVx4_ASAP7_75t_L g1806 ( 
.A(n_1783),
.Y(n_1806)
);

INVxp67_ASAP7_75t_SL g1807 ( 
.A(n_1776),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1750),
.B(n_1726),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1746),
.B(n_1735),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1754),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1756),
.B(n_1662),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1744),
.B(n_1662),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1765),
.B(n_1662),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1752),
.B(n_1720),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1779),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1776),
.B(n_1694),
.Y(n_1816)
);

AND2x2_ASAP7_75t_SL g1817 ( 
.A(n_1768),
.B(n_1718),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1760),
.B(n_1694),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1757),
.Y(n_1819)
);

OAI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1743),
.A2(n_1731),
.B(n_1713),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1757),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1785),
.B(n_1783),
.C(n_1731),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1788),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1789),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1793),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1796),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1803),
.Y(n_1827)
);

AND2x2_ASAP7_75t_SL g1828 ( 
.A(n_1817),
.B(n_1771),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1805),
.Y(n_1829)
);

CKINVDCx16_ASAP7_75t_R g1830 ( 
.A(n_1801),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1799),
.B(n_1783),
.Y(n_1831)
);

NAND4xp75_ASAP7_75t_L g1832 ( 
.A(n_1820),
.B(n_1740),
.C(n_1753),
.D(n_1775),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1810),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1792),
.B(n_1749),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1819),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1821),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1792),
.B(n_1749),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1787),
.Y(n_1838)
);

BUFx3_ASAP7_75t_L g1839 ( 
.A(n_1794),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1806),
.Y(n_1840)
);

INVx1_ASAP7_75t_SL g1841 ( 
.A(n_1802),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1808),
.B(n_1752),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1806),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1798),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_L g1845 ( 
.A1(n_1801),
.A2(n_1615),
.B1(n_1771),
.B2(n_1730),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1806),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1798),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1807),
.B(n_1760),
.Y(n_1848)
);

OR2x2_ASAP7_75t_L g1849 ( 
.A(n_1804),
.B(n_1774),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1832),
.A2(n_1797),
.B1(n_1801),
.B2(n_1795),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1830),
.A2(n_1790),
.B1(n_1801),
.B2(n_1791),
.Y(n_1851)
);

OAI211xp5_ASAP7_75t_L g1852 ( 
.A1(n_1845),
.A2(n_1822),
.B(n_1794),
.C(n_1808),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1828),
.B(n_1817),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1839),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1839),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1839),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1824),
.B(n_1791),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1844),
.Y(n_1858)
);

OAI32xp33_ASAP7_75t_L g1859 ( 
.A1(n_1830),
.A2(n_1809),
.A3(n_1804),
.B1(n_1740),
.B2(n_1816),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1841),
.B(n_1811),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1844),
.Y(n_1861)
);

CKINVDCx16_ASAP7_75t_R g1862 ( 
.A(n_1831),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1842),
.B(n_1814),
.Y(n_1863)
);

AOI322xp5_ASAP7_75t_L g1864 ( 
.A1(n_1838),
.A2(n_1818),
.A3(n_1786),
.B1(n_1813),
.B2(n_1812),
.C1(n_1764),
.C2(n_1780),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1847),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1828),
.B(n_1800),
.Y(n_1866)
);

AOI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1832),
.A2(n_1775),
.B1(n_1763),
.B2(n_1762),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1828),
.B(n_1809),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1847),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1838),
.B(n_1814),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1855),
.B(n_1848),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1854),
.B(n_1834),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1855),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1857),
.B(n_1849),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1863),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1856),
.B(n_1834),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1860),
.B(n_1849),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1868),
.B(n_1837),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1862),
.B(n_1842),
.Y(n_1879)
);

OA21x2_ASAP7_75t_L g1880 ( 
.A1(n_1851),
.A2(n_1843),
.B(n_1840),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1851),
.B(n_1837),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1866),
.B(n_1840),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1870),
.B(n_1843),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1879),
.B(n_1853),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_1880),
.B(n_1850),
.C(n_1852),
.Y(n_1885)
);

NAND4xp25_ASAP7_75t_L g1886 ( 
.A(n_1881),
.B(n_1859),
.C(n_1867),
.D(n_1865),
.Y(n_1886)
);

OAI221xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1878),
.A2(n_1864),
.B1(n_1846),
.B2(n_1869),
.C(n_1858),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1875),
.A2(n_1846),
.B1(n_1615),
.B2(n_1861),
.Y(n_1888)
);

AOI21xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1880),
.A2(n_1874),
.B(n_1871),
.Y(n_1889)
);

NOR2x1_ASAP7_75t_L g1890 ( 
.A(n_1871),
.B(n_1823),
.Y(n_1890)
);

AND2x2_ASAP7_75t_SL g1891 ( 
.A(n_1882),
.B(n_1823),
.Y(n_1891)
);

NAND3xp33_ASAP7_75t_L g1892 ( 
.A(n_1873),
.B(n_1826),
.C(n_1825),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1872),
.A2(n_1836),
.B1(n_1835),
.B2(n_1833),
.C(n_1829),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1876),
.B(n_1825),
.Y(n_1894)
);

INVxp67_ASAP7_75t_L g1895 ( 
.A(n_1890),
.Y(n_1895)
);

AOI221x1_ASAP7_75t_L g1896 ( 
.A1(n_1889),
.A2(n_1883),
.B1(n_1835),
.B2(n_1826),
.C(n_1836),
.Y(n_1896)
);

AND4x1_ASAP7_75t_L g1897 ( 
.A(n_1884),
.B(n_1827),
.C(n_1833),
.D(n_1829),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1891),
.Y(n_1898)
);

XOR2x2_ASAP7_75t_L g1899 ( 
.A(n_1885),
.B(n_1877),
.Y(n_1899)
);

OAI311xp33_ASAP7_75t_L g1900 ( 
.A1(n_1886),
.A2(n_1827),
.A3(n_1761),
.B1(n_1762),
.C1(n_1763),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1895),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1898),
.B(n_1887),
.C(n_1892),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1895),
.Y(n_1903)
);

CKINVDCx20_ASAP7_75t_R g1904 ( 
.A(n_1899),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1897),
.B(n_1894),
.Y(n_1905)
);

OAI32xp33_ASAP7_75t_L g1906 ( 
.A1(n_1900),
.A2(n_1888),
.A3(n_1815),
.B1(n_1761),
.B2(n_1893),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1904),
.A2(n_1731),
.B1(n_1815),
.B2(n_1720),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_SL g1908 ( 
.A1(n_1905),
.A2(n_1896),
.B1(n_1781),
.B2(n_1739),
.Y(n_1908)
);

AO221x1_ASAP7_75t_L g1909 ( 
.A1(n_1901),
.A2(n_1720),
.B1(n_1766),
.B2(n_1778),
.C(n_1770),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1903),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1902),
.B(n_1781),
.Y(n_1911)
);

XOR2x1_ASAP7_75t_L g1912 ( 
.A(n_1911),
.B(n_1906),
.Y(n_1912)
);

OAI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1907),
.A2(n_1731),
.B(n_1782),
.Y(n_1913)
);

NOR3x1_ASAP7_75t_L g1914 ( 
.A(n_1910),
.B(n_1909),
.C(n_1908),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1912),
.B(n_1766),
.Y(n_1915)
);

AOI322xp5_ASAP7_75t_L g1916 ( 
.A1(n_1915),
.A2(n_1914),
.A3(n_1913),
.B1(n_1737),
.B2(n_1733),
.C1(n_1738),
.C2(n_1731),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1916),
.A2(n_1731),
.B1(n_1782),
.B2(n_1784),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1916),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1918),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1917),
.Y(n_1920)
);

OAI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1919),
.A2(n_1784),
.B1(n_1767),
.B2(n_1778),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1920),
.Y(n_1922)
);

OAI22xp5_ASAP7_75t_SL g1923 ( 
.A1(n_1922),
.A2(n_1731),
.B1(n_1543),
.B2(n_1767),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1923),
.B(n_1921),
.Y(n_1924)
);

AOI22xp33_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1770),
.B1(n_1737),
.B2(n_1738),
.Y(n_1925)
);

OA22x2_ASAP7_75t_L g1926 ( 
.A1(n_1925),
.A2(n_1738),
.B1(n_1737),
.B2(n_1733),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1926),
.A2(n_1733),
.B1(n_1737),
.B2(n_1738),
.C(n_1722),
.Y(n_1927)
);

AOI211xp5_ASAP7_75t_L g1928 ( 
.A1(n_1927),
.A2(n_1541),
.B(n_1733),
.C(n_1544),
.Y(n_1928)
);


endmodule