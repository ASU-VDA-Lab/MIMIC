module real_aes_882_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_478;
wire n_356;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_500;
wire n_307;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_0), .B(n_210), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_1), .A2(n_205), .B(n_269), .Y(n_268) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_2), .A2(n_54), .B1(n_92), .B2(n_96), .Y(n_95) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_3), .A2(n_81), .B1(n_160), .B2(n_161), .Y(n_80) );
INVx1_ASAP7_75t_L g160 ( .A(n_3), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_4), .B(n_221), .Y(n_249) );
INVx1_ASAP7_75t_L g189 ( .A(n_5), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_6), .B(n_221), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_7), .A2(n_81), .B1(n_161), .B2(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g510 ( .A(n_7), .Y(n_510) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_8), .A2(n_23), .B1(n_92), .B2(n_93), .Y(n_91) );
NAND2xp33_ASAP7_75t_L g321 ( .A(n_9), .B(n_219), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g146 ( .A1(n_10), .A2(n_57), .B1(n_147), .B2(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g202 ( .A(n_11), .Y(n_202) );
AOI221x1_ASAP7_75t_L g204 ( .A1(n_12), .A2(n_20), .B1(n_205), .B2(n_210), .C(n_217), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g317 ( .A(n_13), .B(n_210), .Y(n_317) );
AO21x2_ASAP7_75t_L g314 ( .A1(n_14), .A2(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_15), .B(n_200), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_16), .B(n_221), .Y(n_303) );
AO21x1_ASAP7_75t_L g243 ( .A1(n_17), .A2(n_210), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g172 ( .A(n_18), .Y(n_172) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_19), .A2(n_171), .B1(n_172), .B2(n_173), .Y(n_170) );
INVx1_ASAP7_75t_L g173 ( .A(n_19), .Y(n_173) );
NAND2x1_ASAP7_75t_L g231 ( .A(n_21), .B(n_221), .Y(n_231) );
NAND2x1_ASAP7_75t_L g277 ( .A(n_22), .B(n_219), .Y(n_277) );
AOI22xp33_ASAP7_75t_SL g501 ( .A1(n_22), .A2(n_81), .B1(n_161), .B2(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_22), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g181 ( .A1(n_23), .A2(n_54), .B1(n_59), .B2(n_182), .C(n_184), .Y(n_181) );
OR2x2_ASAP7_75t_L g203 ( .A(n_24), .B(n_68), .Y(n_203) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_24), .A2(n_68), .B(n_202), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_25), .B(n_219), .Y(n_271) );
INVx3_ASAP7_75t_L g92 ( .A(n_26), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_27), .B(n_221), .Y(n_320) );
OAI22xp5_ASAP7_75t_SL g175 ( .A1(n_28), .A2(n_63), .B1(n_176), .B2(n_177), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_28), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g139 ( .A1(n_29), .A2(n_39), .B1(n_140), .B2(n_142), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_30), .B(n_219), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_31), .A2(n_205), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_SL g101 ( .A(n_32), .Y(n_101) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_33), .A2(n_50), .B1(n_129), .B2(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g191 ( .A(n_34), .Y(n_191) );
AND2x2_ASAP7_75t_L g206 ( .A(n_34), .B(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g216 ( .A(n_34), .B(n_189), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_35), .B(n_210), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g307 ( .A(n_36), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g119 ( .A1(n_37), .A2(n_42), .B1(n_120), .B2(n_124), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_38), .B(n_219), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_40), .A2(n_205), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g522 ( .A(n_40), .Y(n_522) );
AO22x2_ASAP7_75t_L g104 ( .A1(n_41), .A2(n_59), .B1(n_92), .B2(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g166 ( .A1(n_43), .A2(n_69), .B1(n_167), .B2(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_43), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_43), .B(n_219), .Y(n_232) );
INVx1_ASAP7_75t_L g209 ( .A(n_44), .Y(n_209) );
INVx1_ASAP7_75t_L g213 ( .A(n_44), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g85 ( .A1(n_45), .A2(n_64), .B1(n_86), .B2(n_106), .Y(n_85) );
INVx1_ASAP7_75t_L g102 ( .A(n_46), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g109 ( .A1(n_47), .A2(n_60), .B1(n_110), .B2(n_114), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_48), .B(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_49), .A2(n_205), .B(n_230), .Y(n_229) );
AO21x1_ASAP7_75t_L g246 ( .A1(n_51), .A2(n_205), .B(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_52), .B(n_210), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_53), .B(n_210), .Y(n_279) );
INVxp33_ASAP7_75t_L g186 ( .A(n_54), .Y(n_186) );
AND2x2_ASAP7_75t_L g260 ( .A(n_55), .B(n_201), .Y(n_260) );
INVx1_ASAP7_75t_L g207 ( .A(n_56), .Y(n_207) );
INVx1_ASAP7_75t_L g215 ( .A(n_56), .Y(n_215) );
AND2x2_ASAP7_75t_L g281 ( .A(n_58), .B(n_235), .Y(n_281) );
INVxp67_ASAP7_75t_L g185 ( .A(n_59), .Y(n_185) );
AND2x2_ASAP7_75t_L g265 ( .A(n_61), .B(n_235), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_62), .B(n_210), .Y(n_305) );
INVx1_ASAP7_75t_L g177 ( .A(n_63), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_65), .B(n_135), .Y(n_134) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_66), .A2(n_75), .B1(n_154), .B2(n_156), .Y(n_153) );
AND2x2_ASAP7_75t_L g244 ( .A(n_67), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g168 ( .A(n_69), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_69), .B(n_219), .Y(n_304) );
AND2x2_ASAP7_75t_L g238 ( .A(n_70), .B(n_235), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_71), .B(n_221), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_72), .B(n_219), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g301 ( .A1(n_73), .A2(n_205), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_74), .B(n_221), .Y(n_270) );
BUFx2_ASAP7_75t_SL g183 ( .A(n_76), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_77), .A2(n_205), .B(n_319), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_178), .B1(n_192), .B2(n_499), .C(n_500), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_162), .Y(n_79) );
INVxp67_ASAP7_75t_SL g161 ( .A(n_81), .Y(n_161) );
INVxp33_ASAP7_75t_SL g81 ( .A(n_82), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_83), .Y(n_82) );
NOR2x1_ASAP7_75t_L g83 ( .A(n_84), .B(n_133), .Y(n_83) );
NAND4xp25_ASAP7_75t_L g84 ( .A(n_85), .B(n_109), .C(n_119), .D(n_128), .Y(n_84) );
INVx2_ASAP7_75t_SL g86 ( .A(n_87), .Y(n_86) );
INVx8_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x4_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x2_ASAP7_75t_L g112 ( .A(n_89), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g122 ( .A(n_89), .B(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g137 ( .A(n_89), .B(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g89 ( .A(n_90), .B(n_94), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x4_ASAP7_75t_L g108 ( .A(n_91), .B(n_94), .Y(n_108) );
INVx1_ASAP7_75t_L g118 ( .A(n_91), .Y(n_118) );
AND2x2_ASAP7_75t_L g127 ( .A(n_91), .B(n_95), .Y(n_127) );
INVx2_ASAP7_75t_L g93 ( .A(n_92), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
OAI22x1_ASAP7_75t_L g99 ( .A1(n_92), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_92), .Y(n_100) );
INVx1_ASAP7_75t_L g105 ( .A(n_92), .Y(n_105) );
INVxp67_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x2_ASAP7_75t_L g117 ( .A(n_95), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g107 ( .A(n_97), .B(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g116 ( .A(n_97), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g126 ( .A(n_97), .B(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g97 ( .A(n_98), .B(n_103), .Y(n_97) );
AND2x2_ASAP7_75t_L g113 ( .A(n_98), .B(n_104), .Y(n_113) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g123 ( .A(n_99), .B(n_103), .Y(n_123) );
AND2x2_ASAP7_75t_L g138 ( .A(n_99), .B(n_104), .Y(n_138) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_99), .Y(n_152) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x4_ASAP7_75t_L g141 ( .A(n_108), .B(n_113), .Y(n_141) );
AND2x2_ASAP7_75t_L g148 ( .A(n_108), .B(n_123), .Y(n_148) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g130 ( .A(n_113), .B(n_117), .Y(n_130) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx8_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g155 ( .A(n_117), .B(n_123), .Y(n_155) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx6_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g131 ( .A(n_127), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g151 ( .A(n_127), .B(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND4xp25_ASAP7_75t_SL g133 ( .A(n_134), .B(n_139), .C(n_146), .D(n_153), .Y(n_133) );
INVx4_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
INVx6_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g144 ( .A(n_138), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g157 ( .A(n_138), .B(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx6_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx5_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx4f_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_SL g162 ( .A1(n_163), .A2(n_164), .B1(n_174), .B2(n_175), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_164), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B1(n_169), .B2(n_170), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g178 ( .A(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
AND3x1_ASAP7_75t_SL g180 ( .A(n_181), .B(n_187), .C(n_190), .Y(n_180) );
INVxp67_ASAP7_75t_L g508 ( .A(n_181), .Y(n_508) );
CKINVDCx8_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g184 ( .A(n_185), .B(n_186), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_187), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_187), .A2(n_516), .B(n_519), .Y(n_515) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_SL g513 ( .A(n_188), .B(n_190), .Y(n_513) );
AND2x2_ASAP7_75t_L g520 ( .A(n_188), .B(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g208 ( .A(n_189), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_190), .B(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND4xp75_ASAP7_75t_L g193 ( .A(n_194), .B(n_409), .C(n_449), .D(n_478), .Y(n_193) );
NOR2x1_ASAP7_75t_L g194 ( .A(n_195), .B(n_371), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_196), .B(n_328), .Y(n_195) );
AOI21xp5_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_261), .B(n_282), .Y(n_196) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_198), .B(n_224), .Y(n_197) );
AND2x4_ASAP7_75t_L g327 ( .A(n_198), .B(n_287), .Y(n_327) );
INVx1_ASAP7_75t_SL g380 ( .A(n_198), .Y(n_380) );
AOI21xp33_ASAP7_75t_L g415 ( .A1(n_198), .A2(n_416), .B(n_419), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_SL g419 ( .A1(n_198), .A2(n_420), .B(n_421), .C(n_422), .Y(n_419) );
NAND2x1_ASAP7_75t_L g460 ( .A(n_198), .B(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_198), .B(n_421), .Y(n_482) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g285 ( .A(n_199), .Y(n_285) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_199), .Y(n_359) );
OA21x2_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_204), .B(n_223), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_200), .A2(n_267), .B(n_268), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_200), .Y(n_280) );
OA21x2_ASAP7_75t_L g369 ( .A1(n_200), .A2(n_204), .B(n_223), .Y(n_369) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AND2x4_ASAP7_75t_L g245 ( .A(n_202), .B(n_203), .Y(n_245) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_205), .Y(n_499) );
AND2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
BUFx3_ASAP7_75t_L g518 ( .A(n_206), .Y(n_518) );
AND2x6_ASAP7_75t_L g219 ( .A(n_207), .B(n_212), .Y(n_219) );
AND2x4_ASAP7_75t_L g221 ( .A(n_209), .B(n_214), .Y(n_221) );
INVx2_ASAP7_75t_L g521 ( .A(n_209), .Y(n_521) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_216), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_214), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx5_ASAP7_75t_L g222 ( .A(n_216), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_220), .B(n_222), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_222), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_248), .B(n_249), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_257), .B(n_258), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_222), .A2(n_270), .B(n_271), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_222), .A2(n_277), .B(n_278), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_222), .A2(n_303), .B(n_304), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_222), .A2(n_320), .B(n_321), .Y(n_319) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_239), .Y(n_224) );
AND2x2_ASAP7_75t_L g351 ( .A(n_225), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g432 ( .A(n_225), .B(n_287), .Y(n_432) );
INVx1_ASAP7_75t_L g492 ( .A(n_225), .Y(n_492) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g336 ( .A(n_226), .B(n_252), .Y(n_336) );
AND2x2_ASAP7_75t_L g461 ( .A(n_226), .B(n_253), .Y(n_461) );
AND2x2_ASAP7_75t_L g466 ( .A(n_226), .B(n_426), .Y(n_466) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVxp67_ASAP7_75t_L g342 ( .A(n_227), .Y(n_342) );
BUFx3_ASAP7_75t_L g375 ( .A(n_227), .Y(n_375) );
AND2x2_ASAP7_75t_L g421 ( .A(n_227), .B(n_253), .Y(n_421) );
AO21x2_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_234), .B(n_238), .Y(n_227) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_228), .A2(n_234), .B(n_238), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_234), .A2(n_254), .B(n_260), .Y(n_253) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_234), .A2(n_254), .B(n_260), .Y(n_288) );
INVx3_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
BUFx4f_ASAP7_75t_L g315 ( .A(n_237), .Y(n_315) );
AND2x2_ASAP7_75t_L g406 ( .A(n_239), .B(n_284), .Y(n_406) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_252), .Y(n_239) );
AND2x4_ASAP7_75t_L g287 ( .A(n_240), .B(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g398 ( .A(n_240), .B(n_382), .Y(n_398) );
AND2x2_ASAP7_75t_SL g441 ( .A(n_240), .B(n_369), .Y(n_441) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
BUFx2_ASAP7_75t_L g377 ( .A(n_241), .Y(n_377) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g338 ( .A(n_242), .Y(n_338) );
OAI21x1_ASAP7_75t_SL g242 ( .A1(n_243), .A2(n_246), .B(n_250), .Y(n_242) );
INVx1_ASAP7_75t_L g251 ( .A(n_244), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_245), .B(n_251), .Y(n_250) );
INVx1_ASAP7_75t_SL g299 ( .A(n_245), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_245), .A2(n_317), .B(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_252), .B(n_338), .Y(n_341) );
AND2x2_ASAP7_75t_L g426 ( .A(n_252), .B(n_369), .Y(n_426) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g423 ( .A(n_253), .B(n_285), .Y(n_423) );
AND2x2_ASAP7_75t_L g443 ( .A(n_253), .B(n_369), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_255), .B(n_259), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_261), .B(n_332), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_261), .A2(n_455), .B1(n_456), .B2(n_457), .C(n_459), .Y(n_454) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OAI332xp33_ASAP7_75t_L g488 ( .A1(n_262), .A2(n_348), .A3(n_355), .B1(n_414), .B2(n_489), .B3(n_490), .C1(n_491), .C2(n_493), .Y(n_488) );
NAND2x1p5_ASAP7_75t_L g262 ( .A(n_263), .B(n_272), .Y(n_262) );
AND2x2_ASAP7_75t_L g293 ( .A(n_263), .B(n_273), .Y(n_293) );
AND2x2_ASAP7_75t_L g310 ( .A(n_263), .B(n_311), .Y(n_310) );
INVx4_ASAP7_75t_L g323 ( .A(n_263), .Y(n_323) );
AND2x2_ASAP7_75t_SL g383 ( .A(n_263), .B(n_324), .Y(n_383) );
INVx5_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2x1_ASAP7_75t_SL g345 ( .A(n_264), .B(n_311), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_264), .B(n_272), .Y(n_349) );
AND2x2_ASAP7_75t_L g356 ( .A(n_264), .B(n_273), .Y(n_356) );
BUFx2_ASAP7_75t_L g391 ( .A(n_264), .Y(n_391) );
AND2x2_ASAP7_75t_L g446 ( .A(n_264), .B(n_314), .Y(n_446) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
OR2x2_ASAP7_75t_L g313 ( .A(n_272), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g324 ( .A(n_272), .B(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g364 ( .A(n_272), .Y(n_364) );
AND2x2_ASAP7_75t_L g434 ( .A(n_272), .B(n_333), .Y(n_434) );
AND2x2_ASAP7_75t_L g447 ( .A(n_272), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_272), .B(n_448), .Y(n_465) );
INVx4_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_273), .Y(n_331) );
AO21x2_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_280), .B(n_281), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_279), .Y(n_274) );
OAI32xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_289), .A3(n_294), .B1(n_308), .B2(n_326), .Y(n_282) );
INVx2_ASAP7_75t_L g392 ( .A(n_283), .Y(n_392) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g403 ( .A(n_284), .Y(n_403) );
BUFx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g337 ( .A(n_285), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g470 ( .A(n_285), .B(n_375), .Y(n_470) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g382 ( .A(n_288), .Y(n_382) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx2_ASAP7_75t_L g370 ( .A(n_291), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_291), .B(n_413), .Y(n_412) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x4_ASAP7_75t_SL g381 ( .A(n_292), .B(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g458 ( .A(n_292), .Y(n_458) );
AND2x2_ASAP7_75t_L g476 ( .A(n_292), .B(n_338), .Y(n_476) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NOR2xp67_ASAP7_75t_SL g420 ( .A(n_295), .B(n_349), .Y(n_420) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_296), .B(n_331), .Y(n_418) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g494 ( .A(n_297), .B(n_364), .Y(n_494) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g325 ( .A(n_298), .Y(n_325) );
INVx2_ASAP7_75t_L g366 ( .A(n_298), .Y(n_366) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_306), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_299), .B(n_307), .Y(n_306) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_299), .A2(n_300), .B(n_306), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_305), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_309), .B(n_322), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_309), .B(n_368), .Y(n_453) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
AND3x2_ASAP7_75t_L g408 ( .A(n_310), .B(n_355), .C(n_364), .Y(n_408) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_311), .B(n_314), .Y(n_389) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g343 ( .A(n_313), .B(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g333 ( .A(n_314), .Y(n_333) );
INVx1_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
BUFx3_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_314), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x4_ASAP7_75t_L g374 ( .A(n_323), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_323), .B(n_333), .Y(n_417) );
AND2x2_ASAP7_75t_L g373 ( .A(n_324), .B(n_348), .Y(n_373) );
INVx2_ASAP7_75t_L g400 ( .A(n_324), .Y(n_400) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_334), .B(n_339), .C(n_360), .Y(n_328) );
OAI21xp5_ASAP7_75t_L g480 ( .A1(n_329), .A2(n_456), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_332), .B(n_391), .Y(n_390) );
AOI211xp5_ASAP7_75t_SL g410 ( .A1(n_332), .A2(n_411), .B(n_415), .C(n_424), .Y(n_410) );
AND2x2_ASAP7_75t_L g396 ( .A(n_333), .B(n_356), .Y(n_396) );
OR2x2_ASAP7_75t_L g399 ( .A(n_333), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_336), .B(n_441), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_337), .B(n_382), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_337), .A2(n_363), .B1(n_443), .B2(n_446), .C(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g368 ( .A(n_338), .B(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g414 ( .A(n_338), .B(n_369), .Y(n_414) );
OAI221xp5_ASAP7_75t_SL g339 ( .A1(n_340), .A2(n_343), .B1(n_346), .B2(n_350), .C(n_353), .Y(n_339) );
AND2x2_ASAP7_75t_L g485 ( .A(n_340), .B(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g352 ( .A(n_341), .Y(n_352) );
INVx1_ASAP7_75t_L g438 ( .A(n_342), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_343), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g357 ( .A(n_345), .B(n_348), .Y(n_357) );
AND2x2_ASAP7_75t_L g433 ( .A(n_345), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g358 ( .A(n_352), .B(n_359), .Y(n_358) );
OAI21xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_357), .B(n_358), .Y(n_353) );
INVx1_ASAP7_75t_L g477 ( .A(n_354), .Y(n_477) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
AND2x2_ASAP7_75t_L g456 ( .A(n_355), .B(n_383), .Y(n_456) );
AND2x2_ASAP7_75t_SL g429 ( .A(n_356), .B(n_365), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_362), .B(n_367), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g397 ( .A1(n_361), .A2(n_395), .B1(n_398), .B2(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g467 ( .A(n_361), .Y(n_467) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g387 ( .A(n_364), .Y(n_387) );
INVx1_ASAP7_75t_L g448 ( .A(n_366), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g367 ( .A(n_368), .B(n_370), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_368), .B(n_438), .Y(n_489) );
AND2x2_ASAP7_75t_L g457 ( .A(n_369), .B(n_458), .Y(n_457) );
OAI211xp5_ASAP7_75t_L g450 ( .A1(n_370), .A2(n_451), .B(n_454), .C(n_462), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_393), .Y(n_371) );
AOI322xp5_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .A3(n_376), .B1(n_378), .B2(n_383), .C1(n_384), .C2(n_392), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_374), .Y(n_490) );
AND2x2_ASAP7_75t_L g440 ( .A(n_375), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g474 ( .A(n_375), .Y(n_474) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g425 ( .A(n_377), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_SL g431 ( .A(n_377), .B(n_423), .Y(n_431) );
AND2x2_ASAP7_75t_L g455 ( .A(n_377), .B(n_421), .Y(n_455) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx1_ASAP7_75t_L g427 ( .A(n_381), .Y(n_427) );
NAND2xp33_ASAP7_75t_SL g384 ( .A(n_385), .B(n_390), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_SL g430 ( .A1(n_386), .A2(n_431), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_430) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g497 ( .A(n_389), .Y(n_497) );
AOI211xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B(n_397), .C(n_401), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g472 ( .A(n_396), .Y(n_472) );
INVx1_ASAP7_75t_L g404 ( .A(n_398), .Y(n_404) );
OR2x2_ASAP7_75t_L g491 ( .A(n_398), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_SL g487 ( .A(n_399), .Y(n_487) );
AOI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_405), .B(n_407), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_403), .B(n_421), .Y(n_498) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_430), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_413), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g464 ( .A(n_417), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_SL g424 ( .A1(n_425), .A2(n_427), .B(n_428), .Y(n_424) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
AOI31xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .A3(n_442), .B(n_444), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_441), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_466), .B1(n_467), .B2(n_468), .C(n_471), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_475), .B2(n_477), .Y(n_471) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .C(n_495), .Y(n_478) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_480), .B(n_483), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_SL g493 ( .A(n_494), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
OAI222xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_503), .B1(n_509), .B2(n_511), .C1(n_514), .C2(n_522), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_504), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
CKINVDCx16_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
INVxp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
endmodule