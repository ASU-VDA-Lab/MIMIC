module fake_jpeg_1592_n_152 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_12),
.B(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_9),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_35),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_10),
.Y(n_35)
);

BUFx12f_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_17),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_14),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_47),
.B(n_16),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_0),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_25),
.B1(n_30),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_59),
.B1(n_60),
.B2(n_18),
.Y(n_75)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_19),
.A3(n_16),
.B1(n_47),
.B2(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_71),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_58),
.B(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_17),
.B1(n_22),
.B2(n_18),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_62),
.B(n_1),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_34),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_48),
.C(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_83),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_65),
.A2(n_15),
.B(n_19),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_78),
.B(n_93),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_40),
.B(n_44),
.C(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_40),
.B1(n_26),
.B2(n_4),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_58),
.B1(n_73),
.B2(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_58),
.B(n_3),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_67),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_92),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_5),
.B(n_26),
.C(n_57),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_5),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_5),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_96),
.B(n_101),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_100),
.B1(n_108),
.B2(n_89),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_73),
.B(n_53),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_84),
.B(n_91),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_105),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_64),
.B1(n_68),
.B2(n_51),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_85),
.B1(n_90),
.B2(n_56),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_51),
.B1(n_56),
.B2(n_76),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_81),
.C(n_80),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_118),
.B(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_94),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_98),
.C(n_99),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_105),
.C(n_110),
.Y(n_128)
);

INVx2_ASAP7_75t_R g122 ( 
.A(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_97),
.B1(n_95),
.B2(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_109),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_125),
.A2(n_115),
.B1(n_124),
.B2(n_131),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_111),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_126),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_113),
.C(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_119),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_132),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_121),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.C(n_138),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_117),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_138),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_122),
.B(n_123),
.C(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_139),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_135),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_128),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_139),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_146),
.B(n_147),
.C(n_141),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_129),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_149),
.B(n_141),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_134),
.B(n_140),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_137),
.Y(n_151)
);

XNOR2x2_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_130),
.Y(n_152)
);


endmodule