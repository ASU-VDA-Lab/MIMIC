module fake_jpeg_26100_n_273 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_273);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_273;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_3),
.B(n_11),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_20),
.B1(n_23),
.B2(n_18),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

AO22x2_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_32),
.B1(n_30),
.B2(n_35),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_53),
.A2(n_35),
.B1(n_32),
.B2(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_41),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_61),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_20),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_36),
.A2(n_18),
.B1(n_14),
.B2(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_35),
.B1(n_32),
.B2(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_78),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_53),
.B1(n_66),
.B2(n_61),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_76),
.Y(n_88)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_53),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_42),
.A3(n_28),
.B1(n_34),
.B2(n_48),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_80),
.A2(n_31),
.B(n_57),
.C(n_48),
.Y(n_102)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_62),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_91),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_97),
.A2(n_96),
.B1(n_78),
.B2(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_83),
.B(n_21),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx24_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_71),
.B(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_30),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_71),
.B1(n_80),
.B2(n_76),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_102),
.B1(n_104),
.B2(n_93),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_29),
.B(n_77),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_69),
.B1(n_100),
.B2(n_31),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_85),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_118),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_95),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_75),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_86),
.B(n_16),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_16),
.CI(n_25),
.CON(n_146),
.SN(n_146)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_105),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_73),
.B1(n_32),
.B2(n_84),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_104),
.B1(n_93),
.B2(n_84),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_88),
.B1(n_97),
.B2(n_102),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_121),
.B1(n_110),
.B2(n_52),
.Y(n_161)
);

NOR3xp33_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_98),
.C(n_91),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_132),
.Y(n_165)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_129),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_86),
.B1(n_101),
.B2(n_104),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_131),
.A2(n_136),
.B1(n_121),
.B2(n_110),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_14),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_15),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_139),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_143),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_93),
.B1(n_77),
.B2(n_51),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_123),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_142),
.Y(n_167)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_115),
.B(n_17),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_144),
.B(n_19),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_147),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_16),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_58),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_131),
.A2(n_124),
.B(n_116),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_129),
.B(n_134),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_119),
.C(n_106),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_162),
.C(n_140),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_161),
.B1(n_139),
.B2(n_134),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_172),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_130),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_30),
.C(n_27),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_16),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_123),
.Y(n_174)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_145),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_29),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_151),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_150),
.C(n_163),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_186),
.C(n_188),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g178 ( 
.A(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_187),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_172),
.B1(n_157),
.B2(n_160),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_169),
.B(n_167),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_129),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_129),
.C(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_26),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_154),
.B(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_192),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_193),
.A2(n_190),
.B1(n_180),
.B2(n_94),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_185),
.A2(n_160),
.B1(n_152),
.B2(n_167),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_201),
.B1(n_208),
.B2(n_52),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_19),
.B(n_39),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_177),
.A2(n_153),
.B1(n_142),
.B2(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_202),
.B(n_204),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_207),
.B(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_42),
.B1(n_50),
.B2(n_44),
.Y(n_224)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_173),
.A2(n_100),
.B1(n_99),
.B2(n_94),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_183),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_198),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_212),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_175),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_214),
.A2(n_220),
.B1(n_44),
.B2(n_54),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_190),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_225),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_225),
.B1(n_199),
.B2(n_22),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_54),
.C(n_27),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_212),
.C(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_195),
.A2(n_42),
.B1(n_46),
.B2(n_22),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_203),
.A2(n_50),
.B(n_12),
.Y(n_221)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_200),
.A2(n_12),
.B(n_11),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_194),
.A2(n_11),
.B(n_12),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_226)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_54),
.C(n_27),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_10),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_9),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_215),
.C(n_41),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_248),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_8),
.B(n_9),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_246),
.B1(n_239),
.B2(n_248),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_233),
.B(n_27),
.C(n_30),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_230),
.B(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_250),
.B(n_251),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_243),
.A2(n_237),
.B1(n_234),
.B2(n_227),
.Y(n_251)
);

NOR2x1_ASAP7_75t_SL g252 ( 
.A(n_245),
.B(n_237),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_252),
.A2(n_253),
.A3(n_5),
.B1(n_4),
.B2(n_3),
.C1(n_2),
.C2(n_1),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_7),
.B1(n_8),
.B2(n_6),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_256),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_5),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_5),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_261),
.B(n_3),
.C(n_4),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_26),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_262),
.C(n_30),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_26),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_254),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_259),
.C(n_263),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_25),
.C(n_4),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_267),
.C(n_25),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_22),
.B(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_0),
.C(n_29),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_SL g273 ( 
.A1(n_272),
.A2(n_0),
.B(n_234),
.C(n_241),
.Y(n_273)
);


endmodule