module fake_jpeg_30509_n_51 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_51);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_51;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_21),
.Y(n_23)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_25),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_20),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_22),
.B1(n_9),
.B2(n_10),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_3),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_20),
.B(n_18),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_18),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_28),
.B(n_5),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_31),
.C(n_34),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_22),
.B1(n_5),
.B2(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_43),
.B(n_44),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_45),
.A2(n_35),
.B(n_40),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_45),
.B(n_14),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_47),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_48),
.Y(n_51)
);


endmodule