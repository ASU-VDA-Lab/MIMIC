module fake_ariane_1661_n_1138 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1138);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1138;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_349;
wire n_391;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_194;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_202;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_1134;
wire n_485;
wire n_401;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_600;
wire n_481;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_928;
wire n_839;
wire n_1099;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_920;
wire n_1080;
wire n_576;
wire n_843;
wire n_899;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_617;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_217;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_212;
wire n_851;
wire n_278;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_234;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_998;
wire n_999;
wire n_967;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_204;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_1051;
wire n_608;
wire n_959;
wire n_494;
wire n_892;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_934;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_111),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_166),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_83),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_70),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_60),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_193),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_167),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_107),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_39),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_190),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_169),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_5),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_148),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_58),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_51),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_13),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_24),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_8),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_52),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_75),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_170),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_67),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_116),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_72),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_172),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_42),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_112),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_115),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_119),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_174),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_171),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_160),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_79),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_95),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_165),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_11),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_92),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_122),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_162),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_100),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_3),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_44),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_13),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_155),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_82),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_35),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_31),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_118),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_98),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_46),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_163),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_136),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_18),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_219),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_219),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g273 ( 
.A(n_254),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_257),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_223),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_211),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_254),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_207),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_207),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_246),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_210),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_210),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_246),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_195),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_197),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g291 ( 
.A(n_208),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_232),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_250),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_214),
.Y(n_296)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_222),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_224),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_199),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_200),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_247),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_202),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_204),
.Y(n_303)
);

INVxp33_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_260),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_221),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_266),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g308 ( 
.A(n_215),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_220),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_238),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_194),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_256),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_255),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_206),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_267),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_267),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_278),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_268),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_271),
.A2(n_259),
.B1(n_263),
.B2(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_268),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_270),
.A2(n_240),
.B(n_227),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_296),
.Y(n_326)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

AND2x4_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_264),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_275),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_306),
.B(n_236),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_308),
.B(n_245),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_277),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_269),
.B(n_248),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_277),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_226),
.Y(n_342)
);

AOI22x1_ASAP7_75t_SL g343 ( 
.A1(n_274),
.A2(n_265),
.B1(n_262),
.B2(n_244),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_292),
.B(n_196),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_273),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_315),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_282),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_307),
.Y(n_351)
);

AND2x4_ASAP7_75t_L g352 ( 
.A(n_310),
.B(n_226),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_287),
.B(n_198),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_283),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_293),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_284),
.A2(n_228),
.B1(n_242),
.B2(n_241),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_201),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_295),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_279),
.Y(n_363)
);

INVx4_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_285),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_285),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_286),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_288),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_298),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_286),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_226),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_281),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

OAI22xp33_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_280),
.B1(n_301),
.B2(n_313),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_328),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_363),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_359),
.B(n_280),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_340),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_320),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_337),
.B(n_297),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_337),
.B(n_284),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_317),
.B(n_314),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_348),
.B(n_301),
.Y(n_387)
);

NOR2x1p5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_313),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_326),
.B(n_369),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_333),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_320),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_333),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_326),
.B(n_289),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVx2_ASAP7_75t_SL g399 ( 
.A(n_317),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_335),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_335),
.Y(n_401)
);

AND2x6_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_226),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_339),
.B(n_316),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_338),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_339),
.B(n_316),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_335),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_338),
.Y(n_408)
);

OR2x6_ASAP7_75t_L g409 ( 
.A(n_323),
.B(n_290),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_319),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_324),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

AND3x2_ASAP7_75t_L g414 ( 
.A(n_369),
.B(n_281),
.C(n_299),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_349),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_349),
.Y(n_416)
);

INVx5_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_363),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_R g421 ( 
.A(n_343),
.B(n_302),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_355),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_350),
.B(n_303),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_334),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_341),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_321),
.B(n_309),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_341),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_321),
.B(n_318),
.Y(n_432)
);

INVx5_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_361),
.Y(n_435)
);

BUFx6f_ASAP7_75t_SL g436 ( 
.A(n_318),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_372),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_327),
.B(n_346),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_372),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_354),
.B(n_311),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_361),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_365),
.Y(n_443)
);

INVxp33_ASAP7_75t_SL g444 ( 
.A(n_344),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_365),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_L g446 ( 
.A(n_353),
.B(n_203),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_383),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_377),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_351),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_379),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_399),
.B(n_332),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_427),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_376),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_404),
.B(n_406),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_376),
.B(n_368),
.Y(n_462)
);

INVxp33_ASAP7_75t_L g463 ( 
.A(n_386),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_404),
.B(n_318),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_347),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_394),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_444),
.B(n_364),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_327),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_420),
.B(n_329),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_398),
.B(n_329),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_386),
.B(n_329),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_327),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_406),
.B(n_371),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_408),
.B(n_345),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_389),
.B(n_384),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_443),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_388),
.B(n_343),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_408),
.A2(n_325),
.B(n_360),
.Y(n_484)
);

OR2x2_ASAP7_75t_L g485 ( 
.A(n_396),
.B(n_356),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_429),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_385),
.B(n_356),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_388),
.B(n_342),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_R g490 ( 
.A(n_414),
.B(n_325),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_431),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_387),
.B(n_364),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_378),
.B(n_342),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_435),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_447),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_381),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_409),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_409),
.B(n_364),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_381),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_409),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_374),
.B(n_342),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_423),
.B(n_352),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_436),
.B(n_357),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_411),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_441),
.B(n_357),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_357),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_411),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_412),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_430),
.B(n_352),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_412),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_373),
.B(n_352),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_423),
.B(n_350),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_375),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_375),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_380),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_409),
.B(n_325),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_409),
.B(n_350),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_380),
.B(n_358),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_382),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_421),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_446),
.B(n_362),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_382),
.B(n_312),
.Y(n_531)
);

NOR2x1p5_ASAP7_75t_L g532 ( 
.A(n_419),
.B(n_366),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_424),
.Y(n_533)
);

INVx4_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_366),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_469),
.B(n_395),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_463),
.B(n_419),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_461),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_367),
.C(n_419),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_458),
.B(n_419),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_484),
.A2(n_391),
.B(n_390),
.Y(n_541)
);

AND2x6_ASAP7_75t_SL g542 ( 
.A(n_480),
.B(n_367),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_464),
.B(n_440),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_448),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_468),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_459),
.B(n_440),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_450),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_468),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_459),
.B(n_395),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_522),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_455),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_463),
.B(n_440),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_460),
.Y(n_554)
);

NOR3xp33_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_440),
.C(n_403),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_449),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_467),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_484),
.A2(n_479),
.B(n_533),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_460),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_474),
.B(n_370),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_478),
.B(n_473),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_504),
.A2(n_403),
.B1(n_407),
.B2(n_395),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_478),
.B(n_395),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_472),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_476),
.B(n_403),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_502),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_478),
.B(n_403),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g569 ( 
.A1(n_503),
.A2(n_402),
.B1(n_325),
.B2(n_251),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_477),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_462),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_478),
.B(n_407),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_489),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_452),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_530),
.B(n_407),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_454),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_511),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_478),
.A2(n_402),
.B1(n_416),
.B2(n_415),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_501),
.B(n_439),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_502),
.B(n_407),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_525),
.A2(n_424),
.B1(n_391),
.B2(n_393),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_502),
.B(n_390),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_473),
.B(n_415),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_501),
.B(n_416),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_526),
.B(n_418),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_520),
.B(n_418),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_511),
.B(n_507),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_509),
.B(n_422),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_513),
.Y(n_590)
);

NOR3xp33_ASAP7_75t_L g591 ( 
.A(n_492),
.B(n_397),
.C(n_393),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_516),
.B(n_422),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_510),
.B(n_425),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_517),
.B(n_425),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_487),
.B(n_426),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_519),
.B(n_426),
.Y(n_596)
);

AND2x6_ASAP7_75t_SL g597 ( 
.A(n_483),
.B(n_0),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_485),
.B(n_493),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_525),
.A2(n_397),
.B1(n_400),
.B2(n_401),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_531),
.B(n_428),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_518),
.B(n_428),
.Y(n_601)
);

OAI221xp5_ASAP7_75t_L g602 ( 
.A1(n_514),
.A2(n_439),
.B1(n_434),
.B2(n_400),
.C(n_413),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_514),
.B(n_401),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_532),
.B(n_413),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_505),
.Y(n_605)
);

A2O1A1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_530),
.A2(n_434),
.B(n_437),
.C(n_433),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_545),
.Y(n_607)
);

NOR3xp33_ASAP7_75t_SL g608 ( 
.A(n_566),
.B(n_479),
.C(n_521),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_590),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_605),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_605),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_605),
.Y(n_612)
);

INVxp33_ASAP7_75t_L g613 ( 
.A(n_598),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_554),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_538),
.B(n_512),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_548),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_605),
.B(n_505),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_551),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_538),
.B(n_535),
.Y(n_619)
);

AND3x2_ASAP7_75t_SL g620 ( 
.A(n_542),
.B(n_508),
.C(n_503),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_557),
.Y(n_621)
);

AO22x1_ASAP7_75t_L g622 ( 
.A1(n_598),
.A2(n_512),
.B1(n_475),
.B2(n_529),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_574),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_571),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_560),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_562),
.B(n_486),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_567),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_577),
.B(n_508),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_555),
.B(n_488),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_587),
.B(n_470),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_561),
.B(n_475),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_586),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_544),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_547),
.Y(n_636)
);

OR2x6_ASAP7_75t_L g637 ( 
.A(n_573),
.B(n_505),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_593),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_534),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_549),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_SL g641 ( 
.A(n_566),
.B(n_553),
.C(n_537),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_579),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_579),
.B(n_491),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_SL g644 ( 
.A(n_537),
.B(n_490),
.C(n_495),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_567),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_553),
.B(n_470),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_552),
.B(n_556),
.Y(n_647)
);

OAI21xp33_ASAP7_75t_SL g648 ( 
.A1(n_558),
.A2(n_515),
.B(n_497),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_588),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_SL g650 ( 
.A(n_559),
.B(n_490),
.C(n_496),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_565),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_579),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_570),
.B(n_515),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_604),
.B(n_529),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_589),
.Y(n_655)
);

INVx1_ASAP7_75t_SL g656 ( 
.A(n_585),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_540),
.B(n_499),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_539),
.A2(n_528),
.B1(n_506),
.B2(n_524),
.Y(n_658)
);

A2O1A1Ixp33_ASAP7_75t_L g659 ( 
.A1(n_555),
.A2(n_523),
.B(n_527),
.C(n_500),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_539),
.B(n_457),
.Y(n_660)
);

BUFx4f_ASAP7_75t_L g661 ( 
.A(n_584),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_534),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_588),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_595),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_584),
.B(n_465),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_536),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_592),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_594),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_596),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_600),
.B(n_481),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_619),
.B(n_546),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_618),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_625),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_632),
.A2(n_646),
.B(n_648),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_653),
.A2(n_606),
.B(n_541),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_646),
.A2(n_657),
.B(n_659),
.Y(n_676)
);

AOI21xp33_ASAP7_75t_L g677 ( 
.A1(n_613),
.A2(n_568),
.B(n_564),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_662),
.Y(n_678)
);

NAND2x1p5_ASAP7_75t_L g679 ( 
.A(n_661),
.B(n_642),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_657),
.A2(n_603),
.B(n_575),
.Y(n_680)
);

AOI21x1_ASAP7_75t_L g681 ( 
.A1(n_631),
.A2(n_582),
.B(n_601),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_632),
.A2(n_603),
.B(n_591),
.C(n_572),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_659),
.A2(n_580),
.B(n_602),
.Y(n_683)
);

A2O1A1Ixp33_ASAP7_75t_L g684 ( 
.A1(n_650),
.A2(n_591),
.B(n_543),
.C(n_569),
.Y(n_684)
);

AO21x2_ASAP7_75t_L g685 ( 
.A1(n_650),
.A2(n_582),
.B(n_581),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_L g686 ( 
.A1(n_608),
.A2(n_563),
.B(n_550),
.Y(n_686)
);

AOI21xp5_ASAP7_75t_L g687 ( 
.A1(n_631),
.A2(n_580),
.B(n_583),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_642),
.B(n_578),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_668),
.A2(n_498),
.A3(n_494),
.B(n_482),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_656),
.B(n_597),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_614),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_609),
.Y(n_692)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_660),
.A2(n_578),
.B(n_569),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_661),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_610),
.Y(n_695)
);

NAND2x1p5_ASAP7_75t_L g696 ( 
.A(n_611),
.B(n_599),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_647),
.A2(n_433),
.B(n_417),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_626),
.A2(n_433),
.B(n_417),
.Y(n_698)
);

INVx4_ASAP7_75t_L g699 ( 
.A(n_662),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_638),
.B(n_402),
.Y(n_700)
);

AOI21xp5_ASAP7_75t_SL g701 ( 
.A1(n_633),
.A2(n_615),
.B(n_655),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_607),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_626),
.A2(n_433),
.B(n_417),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_643),
.B(n_417),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_664),
.B(n_402),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_658),
.A2(n_433),
.B(n_417),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_611),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_664),
.B(n_402),
.Y(n_708)
);

AOI21x1_ASAP7_75t_L g709 ( 
.A1(n_622),
.A2(n_433),
.B(n_417),
.Y(n_709)
);

CKINVDCx8_ASAP7_75t_R g710 ( 
.A(n_624),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_667),
.A2(n_437),
.B(n_251),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_643),
.A2(n_402),
.B1(n_437),
.B2(n_230),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_637),
.B(n_437),
.Y(n_713)
);

OAI21xp5_ASAP7_75t_L g714 ( 
.A1(n_641),
.A2(n_437),
.B(n_402),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_628),
.B(n_0),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_635),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_669),
.Y(n_717)
);

OAI21x1_ASAP7_75t_L g718 ( 
.A1(n_617),
.A2(n_437),
.B(n_37),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_630),
.B(n_1),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_630),
.B(n_1),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_634),
.B(n_2),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_613),
.B(n_2),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_616),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_636),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_640),
.A2(n_251),
.B(n_234),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_654),
.B(n_641),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_628),
.B(n_3),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_651),
.B(n_4),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_670),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_617),
.A2(n_251),
.B(n_234),
.Y(n_730)
);

AOI21xp5_ASAP7_75t_SL g731 ( 
.A1(n_682),
.A2(n_666),
.B(n_637),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_692),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_676),
.A2(n_639),
.B(n_662),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_674),
.A2(n_639),
.B(n_662),
.Y(n_734)
);

AO31x2_ASAP7_75t_L g735 ( 
.A1(n_684),
.A2(n_629),
.A3(n_621),
.B(n_623),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_716),
.Y(n_736)
);

O2A1O1Ixp5_ASAP7_75t_L g737 ( 
.A1(n_726),
.A2(n_610),
.B(n_612),
.C(n_665),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_675),
.A2(n_706),
.B(n_680),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_683),
.A2(n_645),
.B(n_627),
.Y(n_739)
);

AO31x2_ASAP7_75t_L g740 ( 
.A1(n_693),
.A2(n_652),
.A3(n_612),
.B(n_644),
.Y(n_740)
);

BUFx6f_ASAP7_75t_L g741 ( 
.A(n_673),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_701),
.A2(n_711),
.B(n_687),
.Y(n_742)
);

A2O1A1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_686),
.A2(n_644),
.B(n_608),
.C(n_665),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_710),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_715),
.B(n_637),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_717),
.Y(n_746)
);

AO32x2_ASAP7_75t_L g747 ( 
.A1(n_678),
.A2(n_620),
.A3(n_654),
.B1(n_649),
.B2(n_645),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_714),
.A2(n_671),
.B(n_703),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_694),
.B(n_627),
.Y(n_749)
);

OAI21xp5_ASAP7_75t_L g750 ( 
.A1(n_722),
.A2(n_649),
.B(n_212),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_672),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_717),
.Y(n_752)
);

AO31x2_ASAP7_75t_L g753 ( 
.A1(n_725),
.A2(n_620),
.A3(n_663),
.B(n_234),
.Y(n_753)
);

O2A1O1Ixp5_ASAP7_75t_SL g754 ( 
.A1(n_724),
.A2(n_663),
.B(n_234),
.C(n_237),
.Y(n_754)
);

OAI21x1_ASAP7_75t_L g755 ( 
.A1(n_698),
.A2(n_663),
.B(n_38),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_694),
.B(n_663),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_697),
.A2(n_213),
.B(n_205),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_702),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_721),
.B(n_4),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_681),
.A2(n_40),
.B(n_36),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_723),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_719),
.B(n_217),
.C(n_216),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_688),
.A2(n_239),
.B1(n_235),
.B2(n_233),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_729),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_718),
.A2(n_43),
.B(n_41),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_685),
.A2(n_225),
.B(n_218),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_691),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_685),
.A2(n_229),
.B(n_5),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_720),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_769)
);

AO31x2_ASAP7_75t_L g770 ( 
.A1(n_729),
.A2(n_124),
.A3(n_189),
.B(n_188),
.Y(n_770)
);

OAI21x1_ASAP7_75t_L g771 ( 
.A1(n_709),
.A2(n_47),
.B(n_45),
.Y(n_771)
);

AO31x2_ASAP7_75t_L g772 ( 
.A1(n_730),
.A2(n_125),
.A3(n_187),
.B(n_185),
.Y(n_772)
);

BUFx8_ASAP7_75t_L g773 ( 
.A(n_707),
.Y(n_773)
);

AO31x2_ASAP7_75t_L g774 ( 
.A1(n_705),
.A2(n_121),
.A3(n_184),
.B(n_183),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_688),
.A2(n_6),
.B(n_9),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_690),
.A2(n_677),
.B1(n_727),
.B2(n_700),
.Y(n_776)
);

AOI221xp5_ASAP7_75t_SL g777 ( 
.A1(n_728),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_14),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_712),
.A2(n_10),
.B(n_12),
.C(n_14),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_708),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_696),
.A2(n_49),
.B(n_48),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_695),
.A2(n_15),
.B(n_16),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_707),
.B(n_17),
.Y(n_782)
);

NOR4xp25_ASAP7_75t_L g783 ( 
.A(n_695),
.B(n_18),
.C(n_19),
.D(n_20),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_689),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_678),
.A2(n_19),
.B(n_20),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_699),
.A2(n_21),
.B(n_22),
.Y(n_786)
);

AO31x2_ASAP7_75t_L g787 ( 
.A1(n_689),
.A2(n_132),
.A3(n_182),
.B(n_181),
.Y(n_787)
);

NOR2x1_ASAP7_75t_SL g788 ( 
.A(n_699),
.B(n_21),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_694),
.B(n_22),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_689),
.A2(n_131),
.A3(n_180),
.B(n_179),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_707),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_713),
.Y(n_792)
);

CKINVDCx20_ASAP7_75t_R g793 ( 
.A(n_679),
.Y(n_793)
);

AO31x2_ASAP7_75t_L g794 ( 
.A1(n_713),
.A2(n_129),
.A3(n_178),
.B(n_177),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_704),
.Y(n_795)
);

NAND3xp33_ASAP7_75t_L g796 ( 
.A(n_704),
.B(n_23),
.C(n_24),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_676),
.A2(n_23),
.B(n_25),
.Y(n_797)
);

AO31x2_ASAP7_75t_L g798 ( 
.A1(n_684),
.A2(n_128),
.A3(n_176),
.B(n_175),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_729),
.B(n_25),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_672),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_732),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_796),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_751),
.Y(n_803)
);

INVx6_ASAP7_75t_L g804 ( 
.A(n_773),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_791),
.Y(n_805)
);

BUFx4f_ASAP7_75t_SL g806 ( 
.A(n_741),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_736),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_746),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_776),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_809)
);

OAI21xp33_ASAP7_75t_L g810 ( 
.A1(n_783),
.A2(n_29),
.B(n_30),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_758),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_741),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_SL g813 ( 
.A1(n_768),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_752),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_738),
.A2(n_32),
.B(n_33),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_744),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_782),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_SL g818 ( 
.A1(n_775),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_764),
.B(n_50),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_769),
.A2(n_34),
.B1(n_54),
.B2(n_56),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_761),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_800),
.A2(n_57),
.B1(n_59),
.B2(n_62),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_767),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_759),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_SL g825 ( 
.A1(n_750),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_825)
);

CKINVDCx6p67_ASAP7_75t_R g826 ( 
.A(n_793),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_784),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_745),
.B(n_73),
.Y(n_828)
);

INVx5_ASAP7_75t_L g829 ( 
.A(n_756),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_777),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_756),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_763),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_747),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_795),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_SL g835 ( 
.A1(n_788),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_SL g836 ( 
.A1(n_797),
.A2(n_766),
.B1(n_742),
.B2(n_789),
.Y(n_836)
);

CKINVDCx11_ASAP7_75t_R g837 ( 
.A(n_795),
.Y(n_837)
);

BUFx4f_ASAP7_75t_SL g838 ( 
.A(n_749),
.Y(n_838)
);

BUFx2_ASAP7_75t_R g839 ( 
.A(n_792),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_731),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_762),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_799),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_735),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_735),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_740),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_740),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_778),
.A2(n_743),
.B1(n_779),
.B2(n_785),
.Y(n_847)
);

INVx6_ASAP7_75t_L g848 ( 
.A(n_737),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_787),
.Y(n_849)
);

OAI22xp33_ASAP7_75t_L g850 ( 
.A1(n_786),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_734),
.Y(n_851)
);

CKINVDCx6p67_ASAP7_75t_R g852 ( 
.A(n_747),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_753),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_770),
.Y(n_854)
);

NAND2x1p5_ASAP7_75t_L g855 ( 
.A(n_739),
.B(n_96),
.Y(n_855)
);

OAI22xp33_ASAP7_75t_L g856 ( 
.A1(n_781),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_733),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_770),
.Y(n_858)
);

INVx4_ASAP7_75t_L g859 ( 
.A(n_798),
.Y(n_859)
);

BUFx2_ASAP7_75t_L g860 ( 
.A(n_753),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_757),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_787),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_748),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_863)
);

OAI21x1_ASAP7_75t_L g864 ( 
.A1(n_854),
.A2(n_771),
.B(n_760),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_801),
.B(n_798),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_858),
.A2(n_755),
.B(n_754),
.Y(n_866)
);

OR2x2_ASAP7_75t_L g867 ( 
.A(n_833),
.B(n_807),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_827),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_843),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_808),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_844),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_814),
.B(n_774),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_845),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_848),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_846),
.B(n_794),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_852),
.B(n_790),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_853),
.B(n_780),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_805),
.B(n_794),
.Y(n_878)
);

BUFx3_ASAP7_75t_L g879 ( 
.A(n_848),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_855),
.Y(n_880)
);

INVx2_ASAP7_75t_SL g881 ( 
.A(n_805),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_842),
.B(n_790),
.Y(n_882)
);

OAI21x1_ASAP7_75t_L g883 ( 
.A1(n_862),
.A2(n_765),
.B(n_774),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_821),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_816),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_859),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_823),
.B(n_772),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_857),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_851),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_803),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_815),
.B(n_772),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_859),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_860),
.B(n_117),
.Y(n_893)
);

AO21x2_ASAP7_75t_L g894 ( 
.A1(n_849),
.A2(n_815),
.B(n_830),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_811),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_819),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_855),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_819),
.B(n_120),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_831),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_831),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_810),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_829),
.Y(n_902)
);

BUFx2_ASAP7_75t_SL g903 ( 
.A(n_829),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_810),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_830),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_847),
.A2(n_123),
.B(n_126),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_828),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_829),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_868),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_865),
.B(n_836),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_868),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_905),
.A2(n_904),
.B1(n_901),
.B2(n_847),
.Y(n_912)
);

AO21x2_ASAP7_75t_L g913 ( 
.A1(n_891),
.A2(n_820),
.B(n_802),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_869),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_869),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_868),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_870),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_869),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_871),
.Y(n_919)
);

OA21x2_ASAP7_75t_L g920 ( 
.A1(n_891),
.A2(n_863),
.B(n_840),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_870),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_872),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_871),
.Y(n_923)
);

OA21x2_ASAP7_75t_L g924 ( 
.A1(n_883),
.A2(n_820),
.B(n_809),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_871),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_886),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_873),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_865),
.B(n_812),
.Y(n_928)
);

OA21x2_ASAP7_75t_L g929 ( 
.A1(n_883),
.A2(n_824),
.B(n_802),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_867),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_867),
.Y(n_931)
);

AO21x1_ASAP7_75t_SL g932 ( 
.A1(n_905),
.A2(n_904),
.B(n_901),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_873),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_886),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_881),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_884),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_887),
.B(n_872),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_887),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_906),
.A2(n_813),
.B(n_818),
.Y(n_939)
);

BUFx2_ASAP7_75t_SL g940 ( 
.A(n_910),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_927),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_914),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_927),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_927),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_913),
.Y(n_945)
);

INVxp67_ASAP7_75t_SL g946 ( 
.A(n_937),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_933),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_933),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_938),
.B(n_889),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_930),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_938),
.B(n_888),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_930),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_926),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_932),
.B(n_888),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_933),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_914),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_932),
.B(n_888),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_928),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_909),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_909),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_912),
.A2(n_906),
.B(n_876),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_935),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_959),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_941),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_940),
.Y(n_965)
);

OAI33xp33_ASAP7_75t_L g966 ( 
.A1(n_959),
.A2(n_937),
.A3(n_931),
.B1(n_936),
.B2(n_917),
.B3(n_921),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_942),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_941),
.Y(n_968)
);

OAI211xp5_ASAP7_75t_SL g969 ( 
.A1(n_961),
.A2(n_912),
.B(n_939),
.C(n_917),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_940),
.B(n_931),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_954),
.Y(n_971)
);

NOR2x1p5_ASAP7_75t_L g972 ( 
.A(n_954),
.B(n_826),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_946),
.B(n_910),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_957),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_957),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_950),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_951),
.B(n_910),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_943),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_943),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_977),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_977),
.B(n_945),
.Y(n_981)
);

INVx1_ASAP7_75t_SL g982 ( 
.A(n_973),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_975),
.B(n_951),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_976),
.B(n_952),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_975),
.B(n_949),
.Y(n_985)
);

INVx1_ASAP7_75t_SL g986 ( 
.A(n_971),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_972),
.B(n_949),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_963),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_974),
.B(n_958),
.Y(n_989)
);

OR2x2_ASAP7_75t_L g990 ( 
.A(n_970),
.B(n_945),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_963),
.Y(n_991)
);

OR2x2_ASAP7_75t_L g992 ( 
.A(n_965),
.B(n_945),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_965),
.B(n_945),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_983),
.B(n_985),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_982),
.B(n_964),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_983),
.B(n_962),
.Y(n_996)
);

NAND2x1_ASAP7_75t_L g997 ( 
.A(n_981),
.B(n_953),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_988),
.Y(n_998)
);

NOR2x1_ASAP7_75t_SL g999 ( 
.A(n_980),
.B(n_932),
.Y(n_999)
);

AND2x2_ASAP7_75t_SL g1000 ( 
.A(n_980),
.B(n_929),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_984),
.B(n_968),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_991),
.B(n_978),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_994),
.B(n_986),
.Y(n_1003)
);

OAI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_995),
.A2(n_961),
.B1(n_969),
.B2(n_874),
.Y(n_1004)
);

OAI22xp33_ASAP7_75t_L g1005 ( 
.A1(n_1001),
.A2(n_969),
.B1(n_874),
.B2(n_879),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_996),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_998),
.B(n_989),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_1000),
.B(n_1002),
.Y(n_1008)
);

OAI22xp33_ASAP7_75t_L g1009 ( 
.A1(n_1002),
.A2(n_874),
.B1(n_879),
.B2(n_920),
.Y(n_1009)
);

OR2x2_ASAP7_75t_L g1010 ( 
.A(n_1007),
.B(n_985),
.Y(n_1010)
);

NOR2xp67_ASAP7_75t_L g1011 ( 
.A(n_1006),
.B(n_981),
.Y(n_1011)
);

AOI22xp33_ASAP7_75t_L g1012 ( 
.A1(n_1004),
.A2(n_1000),
.B1(n_1008),
.B2(n_1005),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1003),
.B(n_981),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1009),
.Y(n_1014)
);

INVxp33_ASAP7_75t_L g1015 ( 
.A(n_1003),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_1006),
.B(n_987),
.Y(n_1016)
);

INVxp67_ASAP7_75t_L g1017 ( 
.A(n_1003),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1003),
.B(n_999),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1006),
.B(n_992),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_1015),
.A2(n_993),
.B(n_997),
.Y(n_1020)
);

AND3x2_ASAP7_75t_L g1021 ( 
.A(n_1017),
.B(n_898),
.C(n_806),
.Y(n_1021)
);

NAND2x1_ASAP7_75t_L g1022 ( 
.A(n_1011),
.B(n_990),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1017),
.B(n_885),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1014),
.A2(n_913),
.B1(n_920),
.B2(n_966),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1010),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1019),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1016),
.B(n_993),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_L g1028 ( 
.A(n_1012),
.B(n_939),
.C(n_835),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_1028),
.A2(n_1018),
.B(n_1013),
.C(n_879),
.Y(n_1029)
);

OAI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_1024),
.A2(n_929),
.B1(n_924),
.B2(n_920),
.Y(n_1030)
);

OA21x2_ASAP7_75t_L g1031 ( 
.A1(n_1023),
.A2(n_967),
.B(n_979),
.Y(n_1031)
);

AOI31xp33_ASAP7_75t_L g1032 ( 
.A1(n_1026),
.A2(n_804),
.A3(n_966),
.B(n_898),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_1025),
.B(n_962),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_1021),
.B(n_962),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_1022),
.B(n_953),
.Y(n_1035)
);

AOI211xp5_ASAP7_75t_L g1036 ( 
.A1(n_1020),
.A2(n_850),
.B(n_856),
.C(n_804),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_1027),
.B(n_921),
.Y(n_1037)
);

OAI211xp5_ASAP7_75t_L g1038 ( 
.A1(n_1034),
.A2(n_953),
.B(n_825),
.C(n_935),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_1029),
.A2(n_913),
.B(n_929),
.C(n_893),
.Y(n_1039)
);

OAI32xp33_ASAP7_75t_L g1040 ( 
.A1(n_1035),
.A2(n_893),
.A3(n_953),
.B1(n_967),
.B2(n_876),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1030),
.A2(n_913),
.B1(n_920),
.B2(n_929),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1037),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_1032),
.A2(n_1036),
.B(n_1033),
.C(n_1031),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_1031),
.A2(n_913),
.B(n_929),
.C(n_924),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1037),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1042),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_1045),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1043),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1039),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1044),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_1041),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_1038),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_1040),
.B(n_837),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1042),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1042),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1042),
.B(n_935),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1047),
.Y(n_1057)
);

NOR2x1_ASAP7_75t_L g1058 ( 
.A(n_1046),
.B(n_926),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_1047),
.B(n_832),
.C(n_841),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_L g1060 ( 
.A(n_1048),
.B(n_861),
.C(n_822),
.Y(n_1060)
);

NAND5xp2_ASAP7_75t_L g1061 ( 
.A(n_1053),
.B(n_896),
.C(n_928),
.D(n_907),
.E(n_882),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1054),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_1055),
.B(n_924),
.C(n_920),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1052),
.B(n_817),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1049),
.A2(n_924),
.B1(n_894),
.B2(n_960),
.Y(n_1065)
);

OAI32xp33_ASAP7_75t_L g1066 ( 
.A1(n_1050),
.A2(n_960),
.A3(n_934),
.B1(n_926),
.B2(n_948),
.Y(n_1066)
);

NAND4xp25_ASAP7_75t_L g1067 ( 
.A(n_1056),
.B(n_926),
.C(n_934),
.D(n_896),
.Y(n_1067)
);

AOI21xp33_ASAP7_75t_SL g1068 ( 
.A1(n_1062),
.A2(n_1051),
.B(n_924),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1064),
.A2(n_894),
.B1(n_882),
.B2(n_922),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_1060),
.A2(n_955),
.B(n_948),
.C(n_947),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_L g1071 ( 
.A(n_1057),
.B(n_922),
.C(n_907),
.Y(n_1071)
);

NOR4xp25_ASAP7_75t_L g1072 ( 
.A(n_1067),
.B(n_955),
.C(n_947),
.D(n_944),
.Y(n_1072)
);

NAND3xp33_ASAP7_75t_L g1073 ( 
.A(n_1058),
.B(n_944),
.C(n_936),
.Y(n_1073)
);

NOR2x1_ASAP7_75t_L g1074 ( 
.A(n_1059),
.B(n_926),
.Y(n_1074)
);

AOI211xp5_ASAP7_75t_L g1075 ( 
.A1(n_1072),
.A2(n_1066),
.B(n_1061),
.C(n_1063),
.Y(n_1075)
);

NOR4xp25_ASAP7_75t_L g1076 ( 
.A(n_1070),
.B(n_1073),
.C(n_1074),
.D(n_1068),
.Y(n_1076)
);

AOI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1071),
.A2(n_1065),
.B(n_880),
.C(n_928),
.Y(n_1077)
);

NAND4xp25_ASAP7_75t_L g1078 ( 
.A(n_1069),
.B(n_934),
.C(n_834),
.D(n_900),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1074),
.B(n_942),
.Y(n_1079)
);

NOR3xp33_ASAP7_75t_SL g1080 ( 
.A(n_1070),
.B(n_900),
.C(n_838),
.Y(n_1080)
);

AOI211xp5_ASAP7_75t_L g1081 ( 
.A1(n_1072),
.A2(n_880),
.B(n_878),
.C(n_897),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1074),
.B(n_942),
.Y(n_1082)
);

NOR4xp75_ASAP7_75t_L g1083 ( 
.A(n_1074),
.B(n_934),
.C(n_881),
.D(n_886),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_1076),
.B(n_956),
.Y(n_1084)
);

NOR2x1_ASAP7_75t_L g1085 ( 
.A(n_1078),
.B(n_934),
.Y(n_1085)
);

OA22x2_ASAP7_75t_L g1086 ( 
.A1(n_1079),
.A2(n_956),
.B1(n_903),
.B2(n_892),
.Y(n_1086)
);

NOR3xp33_ASAP7_75t_L g1087 ( 
.A(n_1075),
.B(n_897),
.C(n_866),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1080),
.A2(n_956),
.B(n_866),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_1082),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_1077),
.B(n_897),
.C(n_839),
.Y(n_1090)
);

AND4x1_ASAP7_75t_L g1091 ( 
.A(n_1081),
.B(n_839),
.C(n_903),
.D(n_135),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_1083),
.B(n_880),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_1079),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1092),
.A2(n_1084),
.B1(n_1085),
.B2(n_1086),
.Y(n_1094)
);

NAND4xp75_ASAP7_75t_L g1095 ( 
.A(n_1089),
.B(n_916),
.C(n_911),
.D(n_908),
.Y(n_1095)
);

INVx3_ASAP7_75t_SL g1096 ( 
.A(n_1093),
.Y(n_1096)
);

NOR3x2_ASAP7_75t_L g1097 ( 
.A(n_1087),
.B(n_127),
.C(n_133),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_L g1098 ( 
.A(n_1090),
.B(n_1088),
.C(n_1091),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1084),
.B(n_894),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1084),
.B(n_894),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1092),
.B(n_911),
.Y(n_1101)
);

NAND4xp75_ASAP7_75t_L g1102 ( 
.A(n_1089),
.B(n_916),
.C(n_908),
.D(n_902),
.Y(n_1102)
);

AND2x4_ASAP7_75t_L g1103 ( 
.A(n_1089),
.B(n_880),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1084),
.B(n_892),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1084),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_L g1106 ( 
.A(n_1089),
.B(n_866),
.C(n_138),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1096),
.A2(n_880),
.B1(n_878),
.B2(n_877),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1105),
.B(n_880),
.C(n_878),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_1094),
.A2(n_878),
.B(n_886),
.C(n_902),
.Y(n_1109)
);

NAND4xp25_ASAP7_75t_SL g1110 ( 
.A(n_1098),
.B(n_908),
.C(n_902),
.D(n_899),
.Y(n_1110)
);

XNOR2xp5_ASAP7_75t_L g1111 ( 
.A(n_1097),
.B(n_137),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1106),
.A2(n_875),
.B1(n_877),
.B2(n_884),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_1100),
.B(n_139),
.C(n_140),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_SL g1114 ( 
.A1(n_1103),
.A2(n_875),
.B1(n_883),
.B2(n_864),
.Y(n_1114)
);

NOR2x1_ASAP7_75t_L g1115 ( 
.A(n_1104),
.B(n_141),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1115),
.A2(n_1101),
.B1(n_1099),
.B2(n_1102),
.Y(n_1116)
);

AO22x2_ASAP7_75t_L g1117 ( 
.A1(n_1111),
.A2(n_1095),
.B1(n_899),
.B2(n_875),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1112),
.A2(n_875),
.B1(n_877),
.B2(n_890),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1108),
.A2(n_1114),
.B1(n_1109),
.B2(n_1113),
.Y(n_1119)
);

OAI22x1_ASAP7_75t_L g1120 ( 
.A1(n_1110),
.A2(n_899),
.B1(n_923),
.B2(n_919),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_1107),
.A2(n_925),
.B1(n_923),
.B2(n_919),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1112),
.A2(n_877),
.B1(n_890),
.B2(n_895),
.Y(n_1122)
);

OAI22x1_ASAP7_75t_L g1123 ( 
.A1(n_1118),
.A2(n_142),
.B1(n_143),
.B2(n_146),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1117),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1116),
.B(n_877),
.Y(n_1125)
);

AOI221x1_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_1119),
.B1(n_1117),
.B2(n_1121),
.C(n_1120),
.Y(n_1126)
);

NOR4xp25_ASAP7_75t_L g1127 ( 
.A(n_1126),
.B(n_1125),
.C(n_1123),
.D(n_1122),
.Y(n_1127)
);

OAI21x1_ASAP7_75t_SL g1128 ( 
.A1(n_1127),
.A2(n_147),
.B(n_149),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1128),
.A2(n_864),
.B1(n_923),
.B2(n_919),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1128),
.A2(n_925),
.B1(n_918),
.B2(n_915),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_1128),
.A2(n_925),
.B1(n_918),
.B2(n_915),
.Y(n_1131)
);

AOI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1129),
.A2(n_150),
.B(n_151),
.Y(n_1132)
);

XNOR2xp5_ASAP7_75t_L g1133 ( 
.A(n_1130),
.B(n_152),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_1131),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1134),
.B(n_153),
.Y(n_1135)
);

OA21x2_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_1132),
.B(n_156),
.Y(n_1136)
);

AOI221xp5_ASAP7_75t_L g1137 ( 
.A1(n_1136),
.A2(n_154),
.B1(n_157),
.B2(n_158),
.C(n_159),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_1135),
.B(n_161),
.C(n_164),
.Y(n_1138)
);


endmodule