module fake_netlist_6_3519_n_2823 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_92, n_599, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2823);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_599;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2823;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_1575;
wire n_798;
wire n_2324;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_612;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1796;
wire n_1757;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_811;
wire n_683;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_1837;
wire n_964;
wire n_831;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_2801;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_2439;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_1405;
wire n_972;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1848;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_1362;
wire n_1156;
wire n_829;
wire n_2600;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_88),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_427),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_366),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_558),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_189),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_460),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_476),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_237),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_553),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_200),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_71),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_293),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_306),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_276),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_146),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_588),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_217),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_357),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_557),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_428),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_493),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_452),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_391),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_601),
.Y(n_634)
);

INVx1_ASAP7_75t_SL g635 ( 
.A(n_156),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_444),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_46),
.Y(n_637)
);

CKINVDCx14_ASAP7_75t_R g638 ( 
.A(n_82),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_469),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_74),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_492),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_41),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_305),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_370),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_235),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_561),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_31),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_539),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_260),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_96),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_544),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_500),
.Y(n_652)
);

CKINVDCx14_ASAP7_75t_R g653 ( 
.A(n_484),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_308),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_571),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_234),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_402),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_313),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_126),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_312),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_337),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_475),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_444),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_512),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_455),
.Y(n_665)
);

CKINVDCx16_ASAP7_75t_R g666 ( 
.A(n_338),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_126),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_440),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_180),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_479),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_174),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_432),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_219),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_147),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_455),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_467),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_607),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_477),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_434),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_110),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_176),
.Y(n_681)
);

INVxp67_ASAP7_75t_SL g682 ( 
.A(n_379),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_381),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_472),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_308),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_206),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_592),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_198),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_73),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_132),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_37),
.Y(n_691)
);

BUFx10_ASAP7_75t_L g692 ( 
.A(n_597),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_424),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_478),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_189),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_378),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_291),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_132),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_559),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_157),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_146),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_286),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_610),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_31),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_288),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_388),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_496),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_417),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_407),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_123),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_228),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_115),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_75),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_274),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_260),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_124),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_282),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_397),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_564),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_84),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_453),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_556),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_303),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_173),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_490),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_573),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_356),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_253),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_114),
.Y(n_729)
);

BUFx10_ASAP7_75t_L g730 ( 
.A(n_123),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_53),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_413),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_354),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_71),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_52),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_33),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_50),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_168),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_474),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_519),
.Y(n_740)
);

CKINVDCx20_ASAP7_75t_R g741 ( 
.A(n_167),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_550),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_271),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_266),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_525),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_375),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_13),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_223),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_325),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_324),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_470),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_51),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_139),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_328),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_482),
.Y(n_755)
);

CKINVDCx20_ASAP7_75t_R g756 ( 
.A(n_274),
.Y(n_756)
);

BUFx10_ASAP7_75t_L g757 ( 
.A(n_578),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_397),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_468),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_319),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_224),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_532),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_50),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_84),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_369),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_114),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_587),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_183),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_554),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_480),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_364),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_364),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_187),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_226),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_434),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_133),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_41),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_76),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_590),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_395),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_186),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_341),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_509),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_401),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_268),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_405),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_449),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_85),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_335),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_527),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_471),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_169),
.Y(n_792)
);

CKINVDCx16_ASAP7_75t_R g793 ( 
.A(n_270),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_76),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_224),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_10),
.Y(n_796)
);

BUFx2_ASAP7_75t_L g797 ( 
.A(n_456),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_61),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_104),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_23),
.Y(n_800)
);

BUFx2_ASAP7_75t_SL g801 ( 
.A(n_426),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_494),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_314),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_47),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_428),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_358),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_387),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_64),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_105),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_429),
.Y(n_810)
);

BUFx8_ASAP7_75t_SL g811 ( 
.A(n_211),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_111),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_486),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_180),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_88),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_473),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_78),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_450),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_276),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_221),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_359),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_432),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_345),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_201),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_255),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_489),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_446),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_515),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_291),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_221),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_86),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_545),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_292),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_54),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_421),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_128),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_373),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_232),
.Y(n_838)
);

BUFx5_ASAP7_75t_L g839 ( 
.A(n_476),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_426),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_313),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_593),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_316),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_108),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_289),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_446),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_595),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_240),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_332),
.Y(n_849)
);

BUFx2_ASAP7_75t_L g850 ( 
.A(n_457),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_511),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_61),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_526),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_29),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_336),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_112),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_504),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_380),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_367),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_21),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_839),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_839),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_839),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_839),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_839),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_839),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_839),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_811),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_670),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_619),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_728),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_728),
.Y(n_872)
);

INVxp33_ASAP7_75t_L g873 ( 
.A(n_843),
.Y(n_873)
);

INVxp67_ASAP7_75t_SL g874 ( 
.A(n_783),
.Y(n_874)
);

INVxp33_ASAP7_75t_L g875 ( 
.A(n_671),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_738),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_728),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_728),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_774),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_774),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_824),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_774),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_774),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_761),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_824),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_855),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_855),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_824),
.Y(n_888)
);

INVxp33_ASAP7_75t_L g889 ( 
.A(n_797),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_811),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_855),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_619),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_855),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_628),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_628),
.Y(n_895)
);

CKINVDCx14_ASAP7_75t_R g896 ( 
.A(n_638),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_692),
.Y(n_897)
);

NOR2xp67_ASAP7_75t_L g898 ( 
.A(n_633),
.B(n_0),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_637),
.Y(n_899)
);

INVxp67_ASAP7_75t_SL g900 ( 
.A(n_620),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_620),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_692),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_725),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_804),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_799),
.Y(n_905)
);

CKINVDCx16_ASAP7_75t_R g906 ( 
.A(n_640),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_804),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_859),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_859),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_666),
.Y(n_910)
);

INVxp33_ASAP7_75t_L g911 ( 
.A(n_850),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_612),
.Y(n_912)
);

INVxp33_ASAP7_75t_SL g913 ( 
.A(n_630),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_613),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_725),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_621),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_725),
.Y(n_917)
);

INVxp33_ASAP7_75t_L g918 ( 
.A(n_622),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_627),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_636),
.Y(n_920)
);

INVxp33_ASAP7_75t_L g921 ( 
.A(n_639),
.Y(n_921)
);

INVx1_ASAP7_75t_SL g922 ( 
.A(n_775),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_650),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_793),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_634),
.B(n_0),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_725),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_654),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_654),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_680),
.Y(n_929)
);

NOR2xp67_ASAP7_75t_L g930 ( 
.A(n_709),
.B(n_1),
.Y(n_930)
);

INVxp67_ASAP7_75t_SL g931 ( 
.A(n_629),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_680),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_611),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_661),
.Y(n_934)
);

INVxp33_ASAP7_75t_SL g935 ( 
.A(n_630),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_730),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_616),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_662),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_632),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_663),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_675),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_725),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_678),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_641),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_641),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_681),
.Y(n_946)
);

INVx1_ASAP7_75t_SL g947 ( 
.A(n_730),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_696),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_634),
.B(n_1),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_696),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_692),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_712),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_725),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_725),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_712),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_753),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_753),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_809),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_809),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_858),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_858),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_617),
.Y(n_962)
);

CKINVDCx14_ASAP7_75t_R g963 ( 
.A(n_653),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_683),
.Y(n_964)
);

INVx4_ASAP7_75t_L g965 ( 
.A(n_903),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_871),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_881),
.B(n_655),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_888),
.B(n_655),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_871),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_963),
.B(n_664),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_872),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_861),
.B(n_652),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_903),
.Y(n_973)
);

BUFx8_ASAP7_75t_SL g974 ( 
.A(n_868),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_881),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_885),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_900),
.B(n_664),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_861),
.Y(n_978)
);

BUFx8_ASAP7_75t_SL g979 ( 
.A(n_868),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_885),
.Y(n_980)
);

INVx3_ASAP7_75t_L g981 ( 
.A(n_862),
.Y(n_981)
);

BUFx8_ASAP7_75t_SL g982 ( 
.A(n_890),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_872),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_877),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_877),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_901),
.B(n_709),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_878),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_878),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_904),
.B(n_721),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_879),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_910),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_879),
.Y(n_992)
);

AND2x4_ASAP7_75t_L g993 ( 
.A(n_931),
.B(n_707),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_922),
.B(n_947),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_906),
.B(n_757),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_896),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_880),
.B(n_707),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_874),
.B(n_769),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_915),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_880),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_915),
.Y(n_1001)
);

INVx5_ASAP7_75t_L g1002 ( 
.A(n_917),
.Y(n_1002)
);

INVx5_ASAP7_75t_L g1003 ( 
.A(n_917),
.Y(n_1003)
);

INVx6_ASAP7_75t_L g1004 ( 
.A(n_897),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_890),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_882),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_897),
.B(n_902),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_882),
.B(n_769),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_883),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_883),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_902),
.B(n_699),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_886),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_886),
.Y(n_1013)
);

INVx5_ASAP7_75t_L g1014 ( 
.A(n_926),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_907),
.B(n_908),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_887),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_887),
.Y(n_1017)
);

INVx5_ASAP7_75t_L g1018 ( 
.A(n_926),
.Y(n_1018)
);

INVx4_ASAP7_75t_L g1019 ( 
.A(n_942),
.Y(n_1019)
);

INVx5_ASAP7_75t_L g1020 ( 
.A(n_942),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_891),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_891),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_893),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_893),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_910),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_862),
.B(n_703),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_909),
.B(n_721),
.Y(n_1027)
);

HB1xp67_ASAP7_75t_L g1028 ( 
.A(n_899),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_960),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_863),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_951),
.B(n_842),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1030),
.Y(n_1033)
);

OA21x2_ASAP7_75t_L g1034 ( 
.A1(n_1026),
.A2(n_866),
.B(n_864),
.Y(n_1034)
);

BUFx6f_ASAP7_75t_L g1035 ( 
.A(n_1010),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_970),
.B(n_913),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1030),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_1029),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_981),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_1028),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_981),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_993),
.B(n_865),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_993),
.B(n_865),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_994),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_981),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_981),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_1010),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_1026),
.A2(n_949),
.B(n_925),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_1010),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_1031),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_978),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_1029),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1026),
.B(n_960),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_978),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_1022),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1026),
.B(n_912),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_993),
.B(n_978),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1022),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1022),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_965),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_965),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_1004),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_1007),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_1015),
.B(n_914),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1015),
.B(n_916),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_SL g1066 ( 
.A(n_996),
.B(n_905),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_965),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_993),
.B(n_986),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1029),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1029),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1029),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_971),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_996),
.B(n_933),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_999),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_991),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_986),
.B(n_894),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_965),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_SL g1078 ( 
.A(n_1005),
.B(n_913),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1025),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_968),
.A2(n_867),
.B(n_953),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_973),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_973),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_967),
.B(n_919),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_973),
.B(n_867),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_973),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_966),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1019),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1019),
.B(n_933),
.Y(n_1088)
);

INVx6_ASAP7_75t_L g1089 ( 
.A(n_1019),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_975),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_967),
.B(n_920),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1019),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_966),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_967),
.B(n_923),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_967),
.B(n_1027),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_975),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_969),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_971),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_969),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_1004),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_989),
.B(n_894),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_983),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_987),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_977),
.B(n_937),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_983),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_998),
.B(n_937),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_987),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_985),
.B(n_962),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_989),
.B(n_895),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1006),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_984),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_984),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_975),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1006),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1023),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1011),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_975),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_975),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1027),
.B(n_934),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_999),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1086),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1086),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1051),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1093),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1093),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1040),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_L g1127 ( 
.A(n_1048),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1097),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1097),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1051),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1061),
.B(n_976),
.Y(n_1131)
);

INVx2_ASAP7_75t_SL g1132 ( 
.A(n_1068),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1053),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1050),
.B(n_924),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1061),
.B(n_976),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1061),
.B(n_976),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1099),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1099),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1103),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1103),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1107),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1107),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_SL g1143 ( 
.A(n_1119),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_1063),
.B(n_935),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_1100),
.B(n_997),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1081),
.B(n_976),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1060),
.A2(n_935),
.B1(n_1008),
.B2(n_997),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1081),
.B(n_976),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_1079),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1110),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1110),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1053),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_1035),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_SL g1154 ( 
.A(n_1116),
.B(n_962),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1060),
.A2(n_997),
.B1(n_1008),
.B2(n_801),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_1053),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1081),
.B(n_1116),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1114),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1058),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1098),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1068),
.B(n_1004),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1076),
.B(n_1101),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1067),
.B(n_980),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1058),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1106),
.B(n_995),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1034),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1076),
.B(n_1004),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1054),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1036),
.B(n_631),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1098),
.Y(n_1170)
);

INVxp33_ASAP7_75t_SL g1171 ( 
.A(n_1066),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1102),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1104),
.B(n_875),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1054),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1059),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1035),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1059),
.Y(n_1177)
);

OR2x2_ASAP7_75t_L g1178 ( 
.A(n_1044),
.B(n_939),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1095),
.B(n_631),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1101),
.B(n_889),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1102),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1034),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1032),
.Y(n_1183)
);

OR2x6_ASAP7_75t_L g1184 ( 
.A(n_1108),
.B(n_787),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1088),
.B(n_876),
.C(n_869),
.Y(n_1185)
);

INVx8_ASAP7_75t_L g1186 ( 
.A(n_1095),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1100),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1105),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1119),
.B(n_847),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1119),
.B(n_851),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1105),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1034),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1075),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1034),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1064),
.B(n_851),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1073),
.B(n_911),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1064),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_L g1198 ( 
.A(n_1039),
.B(n_1041),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1111),
.Y(n_1199)
);

NAND2xp33_ASAP7_75t_L g1200 ( 
.A(n_1039),
.B(n_652),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1078),
.A2(n_884),
.B1(n_936),
.B2(n_951),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1111),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1112),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1067),
.B(n_980),
.Y(n_1204)
);

OR2x2_ASAP7_75t_L g1205 ( 
.A(n_1064),
.B(n_1005),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1112),
.Y(n_1206)
);

CKINVDCx14_ASAP7_75t_R g1207 ( 
.A(n_1065),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1115),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1115),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1077),
.B(n_980),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1056),
.B(n_870),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1065),
.B(n_857),
.Y(n_1212)
);

CKINVDCx11_ASAP7_75t_R g1213 ( 
.A(n_1065),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_1056),
.B(n_892),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1041),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1045),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1109),
.B(n_873),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1032),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1062),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1045),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1109),
.B(n_997),
.Y(n_1221)
);

INVx3_ASAP7_75t_L g1222 ( 
.A(n_1089),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1077),
.B(n_980),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1046),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1046),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1056),
.B(n_944),
.Y(n_1226)
);

OR2x2_ASAP7_75t_L g1227 ( 
.A(n_1083),
.B(n_624),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1033),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1082),
.B(n_980),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1089),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_SL g1231 ( 
.A(n_1062),
.B(n_974),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1083),
.B(n_635),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1082),
.B(n_1008),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1083),
.A2(n_945),
.B1(n_615),
.B2(n_642),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1033),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1091),
.B(n_857),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1037),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1037),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1085),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1042),
.A2(n_1043),
.B(n_1057),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1085),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1091),
.B(n_1094),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1091),
.B(n_614),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_SL g1244 ( 
.A(n_1094),
.Y(n_1244)
);

INVx3_ASAP7_75t_L g1245 ( 
.A(n_1089),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1094),
.B(n_626),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1087),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1035),
.B(n_648),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1087),
.B(n_1008),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1092),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_1072),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1092),
.B(n_985),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1084),
.Y(n_1253)
);

HB1xp67_ASAP7_75t_L g1254 ( 
.A(n_1048),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1089),
.B(n_918),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1080),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1220),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1255),
.B(n_1048),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1217),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1157),
.A2(n_1048),
.B(n_1080),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1186),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1144),
.B(n_1035),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1220),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1225),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1225),
.Y(n_1265)
);

INVxp67_ASAP7_75t_SL g1266 ( 
.A(n_1153),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1123),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1132),
.B(n_1035),
.Y(n_1268)
);

INVxp33_ASAP7_75t_SL g1269 ( 
.A(n_1231),
.Y(n_1269)
);

XOR2xp5_ASAP7_75t_L g1270 ( 
.A(n_1207),
.B(n_615),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1123),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1130),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1132),
.B(n_1253),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1130),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1253),
.B(n_1047),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1221),
.B(n_1047),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1168),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1168),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1174),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1153),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1174),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1175),
.Y(n_1282)
);

NAND2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1244),
.B(n_625),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1171),
.B(n_979),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1217),
.B(n_1180),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1175),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1177),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1177),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1215),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1215),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1221),
.B(n_1047),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1188),
.B(n_1047),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1216),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1216),
.Y(n_1294)
);

XOR2xp5_ASAP7_75t_L g1295 ( 
.A(n_1171),
.B(n_625),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1224),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1224),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_L g1298 ( 
.A(n_1173),
.B(n_1047),
.Y(n_1298)
);

AND2x6_ASAP7_75t_L g1299 ( 
.A(n_1166),
.B(n_1038),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1160),
.Y(n_1300)
);

CKINVDCx16_ASAP7_75t_R g1301 ( 
.A(n_1143),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1180),
.B(n_921),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1160),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1178),
.B(n_1049),
.Y(n_1304)
);

XOR2xp5_ASAP7_75t_L g1305 ( 
.A(n_1234),
.B(n_642),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1170),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1170),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1172),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1162),
.Y(n_1309)
);

INVxp67_ASAP7_75t_SL g1310 ( 
.A(n_1153),
.Y(n_1310)
);

INVx2_ASAP7_75t_SL g1311 ( 
.A(n_1149),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1172),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1181),
.Y(n_1313)
);

INVxp67_ASAP7_75t_L g1314 ( 
.A(n_1162),
.Y(n_1314)
);

AND2x2_ASAP7_75t_SL g1315 ( 
.A(n_1127),
.B(n_652),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_SL g1316 ( 
.A(n_1126),
.B(n_982),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1181),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1191),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1191),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1178),
.B(n_1049),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1199),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1134),
.B(n_643),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1197),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1199),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1197),
.Y(n_1325)
);

AND2x2_ASAP7_75t_SL g1326 ( 
.A(n_1127),
.B(n_1254),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1188),
.B(n_1049),
.Y(n_1327)
);

XNOR2x2_ASAP7_75t_L g1328 ( 
.A(n_1196),
.B(n_711),
.Y(n_1328)
);

AND2x2_ASAP7_75t_SL g1329 ( 
.A(n_1127),
.B(n_652),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1202),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1202),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1203),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1203),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1206),
.Y(n_1334)
);

AND2x2_ASAP7_75t_L g1335 ( 
.A(n_1134),
.B(n_898),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1242),
.B(n_1049),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1193),
.B(n_730),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1206),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1208),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1208),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1209),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1154),
.B(n_1049),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1209),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1227),
.B(n_744),
.Y(n_1344)
);

XOR2xp5_ASAP7_75t_L g1345 ( 
.A(n_1205),
.B(n_1185),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1228),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1228),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1235),
.Y(n_1348)
);

NAND2xp33_ASAP7_75t_R g1349 ( 
.A(n_1251),
.B(n_632),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1235),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1241),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1133),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1241),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1133),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1133),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1227),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1233),
.A2(n_1118),
.B(n_1052),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1152),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1152),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1247),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1152),
.Y(n_1361)
);

CKINVDCx20_ASAP7_75t_R g1362 ( 
.A(n_1213),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1156),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1165),
.B(n_1055),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1156),
.Y(n_1365)
);

NOR2xp67_ASAP7_75t_L g1366 ( 
.A(n_1205),
.B(n_1211),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1156),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1167),
.B(n_1055),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1251),
.Y(n_1369)
);

XOR2xp5_ASAP7_75t_L g1370 ( 
.A(n_1242),
.B(n_658),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1247),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1240),
.A2(n_1052),
.B(n_1038),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1159),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1164),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1183),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1218),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1232),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1237),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1213),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1238),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1239),
.Y(n_1381)
);

AND2x2_ASAP7_75t_SL g1382 ( 
.A(n_1239),
.B(n_740),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1121),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1232),
.B(n_744),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_1167),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1121),
.Y(n_1386)
);

INVxp33_ASAP7_75t_L g1387 ( 
.A(n_1214),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1143),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1122),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_1242),
.B(n_1055),
.Y(n_1390)
);

XNOR2xp5_ASAP7_75t_L g1391 ( 
.A(n_1201),
.B(n_658),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1169),
.B(n_744),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1226),
.B(n_729),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1122),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1124),
.Y(n_1395)
);

XOR2xp5_ASAP7_75t_L g1396 ( 
.A(n_1179),
.B(n_665),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1250),
.B(n_1055),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1124),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1125),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1125),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1128),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1184),
.B(n_736),
.Y(n_1402)
);

NAND2xp33_ASAP7_75t_SL g1403 ( 
.A(n_1244),
.B(n_676),
.Y(n_1403)
);

BUFx3_ASAP7_75t_L g1404 ( 
.A(n_1187),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1184),
.B(n_764),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1184),
.B(n_938),
.Y(n_1406)
);

XOR2xp5_ASAP7_75t_L g1407 ( 
.A(n_1243),
.B(n_676),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1184),
.B(n_940),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1128),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1195),
.B(n_1055),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_1189),
.Y(n_1411)
);

CKINVDCx14_ASAP7_75t_R g1412 ( 
.A(n_1161),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1129),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1143),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1129),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1137),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1190),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1250),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1137),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1212),
.B(n_731),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1236),
.B(n_731),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1138),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1219),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1138),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1139),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1139),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1161),
.B(n_941),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1219),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1244),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1140),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1141),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1141),
.Y(n_1432)
);

INVxp33_ASAP7_75t_L g1433 ( 
.A(n_1246),
.Y(n_1433)
);

AND2x2_ASAP7_75t_SL g1434 ( 
.A(n_1198),
.B(n_767),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1187),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1161),
.B(n_943),
.Y(n_1436)
);

AND2x2_ASAP7_75t_SL g1437 ( 
.A(n_1198),
.B(n_779),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1142),
.Y(n_1438)
);

INVx1_ASAP7_75t_SL g1439 ( 
.A(n_1161),
.Y(n_1439)
);

CKINVDCx11_ASAP7_75t_R g1440 ( 
.A(n_1186),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1240),
.B(n_741),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1145),
.B(n_1118),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1249),
.B(n_741),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1142),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1145),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1145),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1150),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1150),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1147),
.B(n_946),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1151),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1222),
.B(n_964),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1166),
.B(n_756),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1155),
.B(n_964),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1158),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1285),
.A2(n_1186),
.B1(n_1248),
.B2(n_1230),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1366),
.A2(n_1186),
.B1(n_1230),
.B2(n_1222),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1297),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1315),
.A2(n_756),
.B1(n_765),
.B2(n_758),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1314),
.B(n_1166),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1441),
.A2(n_1230),
.B1(n_1245),
.B2(n_1222),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1314),
.B(n_1182),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1258),
.A2(n_1245),
.B(n_1135),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1387),
.B(n_1182),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1309),
.B(n_1182),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1311),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1351),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1309),
.B(n_1192),
.Y(n_1467)
);

AO221x1_ASAP7_75t_L g1468 ( 
.A1(n_1356),
.A2(n_1176),
.B1(n_1153),
.B2(n_686),
.C(n_694),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1353),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1441),
.A2(n_1158),
.B1(n_1194),
.B2(n_1192),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1273),
.B(n_1192),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1257),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1360),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1381),
.B(n_1194),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1371),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1259),
.B(n_1153),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1302),
.B(n_682),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1263),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1259),
.B(n_1176),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1418),
.Y(n_1480)
);

BUFx6f_ASAP7_75t_L g1481 ( 
.A(n_1440),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_1435),
.Y(n_1482)
);

INVx4_ASAP7_75t_L g1483 ( 
.A(n_1261),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1440),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1385),
.B(n_1194),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1262),
.B(n_1298),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1317),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1369),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1298),
.B(n_1163),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1443),
.A2(n_1204),
.B1(n_1223),
.B2(n_1210),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1264),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1443),
.B(n_930),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1304),
.B(n_1229),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1265),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1420),
.A2(n_645),
.B1(n_747),
.B2(n_644),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1320),
.B(n_1252),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1452),
.B(n_1176),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_SL g1498 ( 
.A(n_1382),
.B(n_1176),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1382),
.A2(n_1420),
.B1(n_1421),
.B2(n_1434),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1412),
.A2(n_651),
.B1(n_687),
.B2(n_677),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1266),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1267),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1373),
.B(n_1131),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1322),
.B(n_1256),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1374),
.B(n_1136),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1412),
.A2(n_719),
.B1(n_726),
.B2(n_722),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1375),
.B(n_1146),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1271),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1421),
.A2(n_813),
.B1(n_853),
.B2(n_832),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1376),
.B(n_1148),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1377),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1321),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1378),
.B(n_1256),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1434),
.A2(n_646),
.B1(n_757),
.B2(n_1069),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1380),
.B(n_1070),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1324),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1282),
.B(n_1070),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1272),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1426),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1404),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1450),
.Y(n_1521)
);

NOR2xp67_ASAP7_75t_L g1522 ( 
.A(n_1356),
.B(n_742),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1336),
.Y(n_1523)
);

INVxp33_ASAP7_75t_L g1524 ( 
.A(n_1370),
.Y(n_1524)
);

INVx8_ASAP7_75t_L g1525 ( 
.A(n_1261),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1274),
.B(n_1071),
.Y(n_1526)
);

INVxp67_ASAP7_75t_L g1527 ( 
.A(n_1335),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1337),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1286),
.B(n_1071),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1387),
.B(n_758),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1261),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1423),
.B(n_745),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1428),
.B(n_762),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1277),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1287),
.B(n_1023),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1261),
.Y(n_1536)
);

BUFx12f_ASAP7_75t_L g1537 ( 
.A(n_1388),
.Y(n_1537)
);

BUFx8_ASAP7_75t_L g1538 ( 
.A(n_1406),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1289),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1278),
.B(n_1090),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1279),
.B(n_1090),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_SL g1542 ( 
.A(n_1439),
.B(n_790),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_SL g1543 ( 
.A(n_1404),
.Y(n_1543)
);

BUFx6f_ASAP7_75t_SL g1544 ( 
.A(n_1336),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1408),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1437),
.A2(n_757),
.B1(n_772),
.B2(n_765),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1427),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1393),
.B(n_772),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1288),
.B(n_1090),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_SL g1550 ( 
.A1(n_1305),
.A2(n_810),
.B1(n_817),
.B2(n_815),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1437),
.A2(n_815),
.B1(n_817),
.B2(n_810),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1281),
.B(n_1090),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1436),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1344),
.B(n_823),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1346),
.B(n_1090),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1347),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1348),
.B(n_1096),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1384),
.B(n_823),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1350),
.B(n_1096),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1290),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1300),
.B(n_1096),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1446),
.A2(n_802),
.B1(n_828),
.B2(n_826),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1315),
.A2(n_787),
.B1(n_693),
.B2(n_698),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1449),
.B(n_1096),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1402),
.B(n_895),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1446),
.B(n_1113),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_L g1567 ( 
.A(n_1445),
.B(n_1113),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1295),
.B(n_618),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1451),
.B(n_927),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1303),
.B(n_1113),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1293),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1405),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1306),
.B(n_1113),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1392),
.B(n_927),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1396),
.B(n_623),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1433),
.B(n_1113),
.Y(n_1576)
);

BUFx8_ASAP7_75t_L g1577 ( 
.A(n_1451),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1414),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1442),
.Y(n_1579)
);

O2A1O1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1342),
.A2(n_1433),
.B(n_1275),
.C(n_1308),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1453),
.B(n_1117),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1307),
.B(n_1117),
.Y(n_1582)
);

BUFx3_ASAP7_75t_L g1583 ( 
.A(n_1429),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1329),
.A2(n_705),
.B1(n_708),
.B2(n_691),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1312),
.B(n_1117),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1329),
.B(n_1117),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1313),
.B(n_1117),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1368),
.A2(n_1291),
.B(n_1276),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1349),
.A2(n_645),
.B1(n_747),
.B2(n_644),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1318),
.B(n_647),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1294),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1326),
.B(n_649),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1296),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1319),
.Y(n_1594)
);

O2A1O1Ixp5_ASAP7_75t_L g1595 ( 
.A1(n_1364),
.A2(n_717),
.B(n_718),
.C(n_714),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1411),
.A2(n_1200),
.B1(n_972),
.B2(n_657),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1407),
.B(n_656),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1345),
.B(n_1270),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1301),
.B(n_928),
.Y(n_1599)
);

INVx4_ASAP7_75t_L g1600 ( 
.A(n_1442),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1330),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1331),
.B(n_659),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1411),
.B(n_928),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_SL g1604 ( 
.A(n_1326),
.B(n_660),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1269),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1417),
.B(n_667),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1332),
.B(n_668),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1364),
.B(n_669),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1333),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1266),
.A2(n_1310),
.B1(n_1280),
.B2(n_1334),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_SL g1611 ( 
.A(n_1410),
.B(n_672),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1338),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1328),
.A2(n_1200),
.B1(n_733),
.B2(n_734),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1339),
.B(n_673),
.Y(n_1614)
);

BUFx3_ASAP7_75t_L g1615 ( 
.A(n_1325),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1340),
.B(n_674),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1280),
.A2(n_1310),
.B1(n_1343),
.B2(n_1341),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1352),
.B(n_953),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1383),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1354),
.B(n_954),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1386),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1355),
.B(n_954),
.Y(n_1622)
);

INVx8_ASAP7_75t_L g1623 ( 
.A(n_1299),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1417),
.B(n_1391),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1284),
.B(n_679),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1410),
.A2(n_972),
.B1(n_685),
.B2(n_688),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1358),
.B(n_972),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1389),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1283),
.B(n_684),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1394),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1359),
.B(n_689),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_SL g1632 ( 
.A(n_1361),
.B(n_690),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1395),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1363),
.B(n_972),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1365),
.B(n_972),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1283),
.A2(n_972),
.B1(n_697),
.B2(n_700),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1349),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1403),
.A2(n_972),
.B1(n_701),
.B2(n_702),
.Y(n_1638)
);

INVx4_ASAP7_75t_L g1639 ( 
.A(n_1299),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1367),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1398),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1399),
.B(n_985),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1454),
.B(n_985),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1400),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_SL g1645 ( 
.A(n_1403),
.B(n_695),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1379),
.B(n_704),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1401),
.B(n_985),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1409),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1325),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1413),
.B(n_988),
.Y(n_1650)
);

NOR3xp33_ASAP7_75t_L g1651 ( 
.A(n_1323),
.B(n_710),
.C(n_706),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1268),
.B(n_713),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1415),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1416),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_SL g1655 ( 
.A(n_1292),
.B(n_715),
.Y(n_1655)
);

INVxp33_ASAP7_75t_SL g1656 ( 
.A(n_1316),
.Y(n_1656)
);

A2O1A1Ixp33_ASAP7_75t_L g1657 ( 
.A1(n_1260),
.A2(n_746),
.B(n_752),
.C(n_723),
.Y(n_1657)
);

NAND2xp33_ASAP7_75t_SL g1658 ( 
.A(n_1362),
.B(n_837),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_R g1659 ( 
.A(n_1362),
.B(n_837),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1499),
.B(n_1547),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1548),
.B(n_1419),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1504),
.B(n_1422),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1486),
.A2(n_1260),
.B(n_1357),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1489),
.A2(n_1397),
.B(n_1327),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1588),
.A2(n_1390),
.B(n_1372),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1492),
.B(n_1424),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1623),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1462),
.A2(n_1430),
.B(n_1425),
.Y(n_1669)
);

A2O1A1Ixp33_ASAP7_75t_L g1670 ( 
.A1(n_1580),
.A2(n_1432),
.B(n_1438),
.C(n_1431),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1603),
.B(n_1444),
.Y(n_1671)
);

AND2x6_ASAP7_75t_L g1672 ( 
.A(n_1536),
.B(n_1447),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1477),
.B(n_1448),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1493),
.A2(n_1001),
.B(n_999),
.Y(n_1674)
);

AND2x2_ASAP7_75t_SL g1675 ( 
.A(n_1551),
.B(n_759),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1657),
.A2(n_1299),
.B(n_768),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1637),
.B(n_716),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1496),
.A2(n_1001),
.B(n_999),
.Y(n_1678)
);

NAND2x1p5_ASAP7_75t_L g1679 ( 
.A(n_1483),
.B(n_1299),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1458),
.A2(n_849),
.B1(n_852),
.B2(n_838),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1574),
.B(n_1299),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1652),
.B(n_760),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1628),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1567),
.A2(n_1001),
.B(n_999),
.Y(n_1684)
);

BUFx6f_ASAP7_75t_L g1685 ( 
.A(n_1536),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1565),
.B(n_770),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1539),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1463),
.B(n_771),
.Y(n_1688)
);

O2A1O1Ixp5_ASAP7_75t_L g1689 ( 
.A1(n_1586),
.A2(n_780),
.B(n_791),
.C(n_773),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1553),
.B(n_795),
.Y(n_1690)
);

BUFx12f_ASAP7_75t_L g1691 ( 
.A(n_1482),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1497),
.A2(n_1001),
.B(n_999),
.Y(n_1692)
);

A2O1A1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1629),
.A2(n_806),
.B(n_812),
.C(n_800),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1572),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1530),
.A2(n_724),
.B1(n_727),
.B2(n_720),
.Y(n_1695)
);

CKINVDCx8_ASAP7_75t_R g1696 ( 
.A(n_1481),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1564),
.A2(n_1003),
.B(n_1002),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1560),
.Y(n_1698)
);

INVx4_ASAP7_75t_L g1699 ( 
.A(n_1525),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1501),
.A2(n_1003),
.B(n_1002),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1472),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1490),
.A2(n_816),
.B(n_814),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1571),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1581),
.A2(n_1003),
.B(n_1002),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1545),
.B(n_827),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1554),
.B(n_929),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1597),
.A2(n_735),
.B1(n_737),
.B2(n_732),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1458),
.A2(n_834),
.B(n_840),
.C(n_830),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1527),
.B(n_841),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1546),
.A2(n_849),
.B1(n_852),
.B2(n_838),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1606),
.B(n_739),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_SL g1712 ( 
.A(n_1488),
.B(n_856),
.Y(n_1712)
);

BUFx3_ASAP7_75t_L g1713 ( 
.A(n_1520),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1575),
.B(n_743),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1584),
.A2(n_1509),
.B1(n_1563),
.B2(n_1478),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1464),
.B(n_844),
.Y(n_1716)
);

O2A1O1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1495),
.A2(n_846),
.B(n_848),
.C(n_845),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1511),
.B(n_748),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_L g1719 ( 
.A(n_1483),
.B(n_1531),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1595),
.A2(n_854),
.B(n_929),
.Y(n_1720)
);

AOI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1498),
.A2(n_948),
.B(n_932),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1491),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1494),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1558),
.B(n_856),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1591),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1464),
.B(n_749),
.Y(n_1726)
);

AND2x6_ASAP7_75t_L g1727 ( 
.A(n_1536),
.B(n_932),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1465),
.B(n_1605),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1467),
.B(n_750),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1528),
.B(n_751),
.Y(n_1730)
);

AOI21x1_ASAP7_75t_L g1731 ( 
.A1(n_1617),
.A2(n_950),
.B(n_948),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1471),
.A2(n_1003),
.B(n_1002),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1467),
.B(n_754),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1471),
.A2(n_1014),
.B(n_1003),
.Y(n_1734)
);

INVx11_ASAP7_75t_L g1735 ( 
.A(n_1577),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1503),
.B(n_755),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1543),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1543),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1505),
.A2(n_1014),
.B(n_1003),
.Y(n_1739)
);

AOI21x1_ASAP7_75t_L g1740 ( 
.A1(n_1617),
.A2(n_1643),
.B(n_1642),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_SL g1741 ( 
.A(n_1656),
.B(n_763),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1593),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1502),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1569),
.B(n_950),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1584),
.A2(n_776),
.B1(n_777),
.B2(n_766),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1598),
.A2(n_781),
.B1(n_782),
.B2(n_778),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1524),
.B(n_784),
.Y(n_1747)
);

AO21x1_ASAP7_75t_L g1748 ( 
.A1(n_1563),
.A2(n_955),
.B(n_952),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1470),
.A2(n_1460),
.B(n_1459),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1645),
.A2(n_955),
.B(n_956),
.C(n_952),
.Y(n_1750)
);

BUFx4f_ASAP7_75t_L g1751 ( 
.A(n_1481),
.Y(n_1751)
);

A2O1A1Ixp33_ASAP7_75t_L g1752 ( 
.A1(n_1455),
.A2(n_786),
.B(n_788),
.C(n_785),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1507),
.A2(n_1018),
.B(n_1014),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1594),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1510),
.B(n_789),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1569),
.B(n_956),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1508),
.B(n_792),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1600),
.B(n_794),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1568),
.B(n_957),
.Y(n_1759)
);

O2A1O1Ixp5_ASAP7_75t_L g1760 ( 
.A1(n_1611),
.A2(n_958),
.B(n_959),
.C(n_957),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1518),
.B(n_796),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1550),
.B(n_798),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1534),
.B(n_803),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1610),
.A2(n_1018),
.B(n_1014),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1608),
.A2(n_807),
.B(n_808),
.C(n_805),
.Y(n_1765)
);

INVx2_ASAP7_75t_SL g1766 ( 
.A(n_1538),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1556),
.B(n_818),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1610),
.A2(n_1018),
.B(n_1014),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1523),
.B(n_819),
.Y(n_1769)
);

BUFx4f_ASAP7_75t_L g1770 ( 
.A(n_1481),
.Y(n_1770)
);

O2A1O1Ixp5_ASAP7_75t_L g1771 ( 
.A1(n_1592),
.A2(n_961),
.B(n_1120),
.C(n_1074),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1544),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1619),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1523),
.B(n_820),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1600),
.B(n_1579),
.Y(n_1775)
);

NOR2x1_ASAP7_75t_L g1776 ( 
.A(n_1531),
.B(n_961),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1601),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1474),
.A2(n_1655),
.B(n_1623),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1578),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1579),
.B(n_821),
.Y(n_1780)
);

AOI21xp5_ASAP7_75t_L g1781 ( 
.A1(n_1474),
.A2(n_1018),
.B(n_1014),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1459),
.B(n_822),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1630),
.Y(n_1783)
);

OAI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1461),
.A2(n_829),
.B(n_825),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1461),
.B(n_1607),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1590),
.B(n_831),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1624),
.B(n_833),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1609),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1623),
.A2(n_1020),
.B(n_1018),
.Y(n_1789)
);

INVx4_ASAP7_75t_L g1790 ( 
.A(n_1525),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1602),
.B(n_1616),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1604),
.B(n_835),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1513),
.A2(n_1020),
.B(n_1018),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1612),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1639),
.A2(n_1020),
.B(n_1074),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1625),
.B(n_836),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1639),
.A2(n_1020),
.B(n_1074),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1614),
.B(n_860),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1522),
.B(n_1599),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1640),
.B(n_2),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1457),
.B(n_2),
.Y(n_1801)
);

BUFx3_ASAP7_75t_L g1802 ( 
.A(n_1583),
.Y(n_1802)
);

O2A1O1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1589),
.A2(n_5),
.B(n_3),
.C(n_4),
.Y(n_1803)
);

AND2x4_ASAP7_75t_L g1804 ( 
.A(n_1484),
.B(n_483),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1646),
.A2(n_990),
.B1(n_992),
.B2(n_988),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1542),
.B(n_1631),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1466),
.B(n_3),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1469),
.B(n_4),
.Y(n_1808)
);

INVx4_ASAP7_75t_L g1809 ( 
.A(n_1525),
.Y(n_1809)
);

INVx6_ASAP7_75t_L g1810 ( 
.A(n_1538),
.Y(n_1810)
);

BUFx10_ASAP7_75t_L g1811 ( 
.A(n_1484),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1485),
.A2(n_1020),
.B(n_1120),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1473),
.B(n_5),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1475),
.B(n_6),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1456),
.A2(n_1020),
.B(n_1120),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1519),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1480),
.B(n_6),
.Y(n_1817)
);

O2A1O1Ixp5_ASAP7_75t_L g1818 ( 
.A1(n_1576),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_1818)
);

O2A1O1Ixp5_ASAP7_75t_L g1819 ( 
.A1(n_1476),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1521),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1561),
.A2(n_990),
.B(n_988),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1618),
.A2(n_990),
.B(n_988),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1561),
.A2(n_992),
.B(n_990),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1651),
.B(n_992),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1487),
.B(n_10),
.Y(n_1825)
);

O2A1O1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1632),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1512),
.B(n_1516),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1570),
.A2(n_1000),
.B(n_992),
.Y(n_1828)
);

AND2x2_ASAP7_75t_SL g1829 ( 
.A(n_1484),
.B(n_11),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1633),
.B(n_12),
.Y(n_1830)
);

AOI21xp5_ASAP7_75t_L g1831 ( 
.A1(n_1570),
.A2(n_1000),
.B(n_992),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1641),
.B(n_14),
.Y(n_1832)
);

OAI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1618),
.A2(n_1009),
.B(n_1000),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1544),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1573),
.A2(n_1009),
.B(n_1000),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1644),
.B(n_14),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1648),
.B(n_485),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1573),
.A2(n_1009),
.B(n_1000),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1577),
.B(n_1009),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1653),
.B(n_15),
.Y(n_1840)
);

BUFx12f_ASAP7_75t_L g1841 ( 
.A(n_1537),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1654),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1526),
.Y(n_1843)
);

AOI21xp5_ASAP7_75t_L g1844 ( 
.A1(n_1582),
.A2(n_1012),
.B(n_1009),
.Y(n_1844)
);

OAI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1620),
.A2(n_1013),
.B(n_1012),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1585),
.A2(n_1013),
.B(n_1012),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1587),
.A2(n_1013),
.B(n_1012),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1535),
.B(n_15),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1526),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1515),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_R g1851 ( 
.A(n_1696),
.B(n_1658),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1711),
.A2(n_1506),
.B1(n_1500),
.B2(n_1562),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1671),
.B(n_1613),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1701),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1714),
.B(n_1787),
.Y(n_1855)
);

AOI22x1_ASAP7_75t_L g1856 ( 
.A1(n_1702),
.A2(n_1468),
.B1(n_1649),
.B2(n_1638),
.Y(n_1856)
);

O2A1O1Ixp33_ASAP7_75t_SL g1857 ( 
.A1(n_1752),
.A2(n_1479),
.B(n_1533),
.C(n_1532),
.Y(n_1857)
);

NOR2xp33_ASAP7_75t_L g1858 ( 
.A(n_1747),
.B(n_1615),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1682),
.A2(n_1675),
.B(n_1695),
.Y(n_1859)
);

OAI321xp33_ASAP7_75t_L g1860 ( 
.A1(n_1803),
.A2(n_1636),
.A3(n_1514),
.B1(n_1626),
.B2(n_1596),
.C(n_1566),
.Y(n_1860)
);

NOR2xp67_ASAP7_75t_SL g1861 ( 
.A(n_1691),
.B(n_1620),
.Y(n_1861)
);

O2A1O1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1693),
.A2(n_1529),
.B(n_1517),
.C(n_1540),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_SL g1863 ( 
.A(n_1799),
.B(n_1659),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1699),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1666),
.A2(n_1541),
.B(n_1540),
.Y(n_1865)
);

AOI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1731),
.A2(n_1650),
.B(n_1647),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1791),
.A2(n_1552),
.B1(n_1555),
.B2(n_1541),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1661),
.A2(n_1552),
.B1(n_1559),
.B2(n_1555),
.Y(n_1868)
);

BUFx2_ASAP7_75t_L g1869 ( 
.A(n_1713),
.Y(n_1869)
);

AND2x2_ASAP7_75t_SL g1870 ( 
.A(n_1829),
.B(n_1549),
.Y(n_1870)
);

NOR2xp33_ASAP7_75t_L g1871 ( 
.A(n_1741),
.B(n_1622),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1792),
.A2(n_1622),
.B1(n_1557),
.B2(n_1627),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1685),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1665),
.A2(n_1650),
.B(n_1647),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1722),
.Y(n_1875)
);

INVx4_ASAP7_75t_L g1876 ( 
.A(n_1699),
.Y(n_1876)
);

O2A1O1Ixp5_ASAP7_75t_L g1877 ( 
.A1(n_1702),
.A2(n_1634),
.B(n_1635),
.C(n_1627),
.Y(n_1877)
);

AOI21x1_ASAP7_75t_L g1878 ( 
.A1(n_1740),
.A2(n_1635),
.B(n_1634),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1790),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1664),
.A2(n_1013),
.B(n_1012),
.Y(n_1880)
);

INVx6_ASAP7_75t_L g1881 ( 
.A(n_1811),
.Y(n_1881)
);

OAI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1786),
.A2(n_1798),
.B(n_1667),
.Y(n_1882)
);

OAI22x1_ASAP7_75t_L g1883 ( 
.A1(n_1762),
.A2(n_1806),
.B1(n_1804),
.B2(n_1842),
.Y(n_1883)
);

AND2x2_ASAP7_75t_SL g1884 ( 
.A(n_1751),
.B(n_16),
.Y(n_1884)
);

OR2x6_ASAP7_75t_L g1885 ( 
.A(n_1810),
.B(n_1013),
.Y(n_1885)
);

A2O1A1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1717),
.A2(n_1017),
.B(n_1021),
.C(n_1016),
.Y(n_1886)
);

OAI22xp5_ASAP7_75t_L g1887 ( 
.A1(n_1673),
.A2(n_1017),
.B1(n_1021),
.B2(n_1016),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1723),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1743),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1694),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1741),
.B(n_1016),
.Y(n_1891)
);

AOI21xp5_ASAP7_75t_L g1892 ( 
.A1(n_1664),
.A2(n_1017),
.B(n_1016),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1834),
.B(n_487),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1660),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_SL g1895 ( 
.A(n_1662),
.B(n_1016),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1683),
.Y(n_1896)
);

NAND2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1790),
.B(n_1017),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1663),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1773),
.Y(n_1899)
);

CKINVDCx6p67_ASAP7_75t_R g1900 ( 
.A(n_1841),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1796),
.B(n_488),
.Y(n_1901)
);

NOR2xp67_ASAP7_75t_L g1902 ( 
.A(n_1834),
.B(n_491),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1718),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1685),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1822),
.A2(n_1024),
.B(n_1021),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1822),
.A2(n_1024),
.B(n_1021),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1785),
.B(n_1759),
.Y(n_1907)
);

A2O1A1Ixp33_ASAP7_75t_L g1908 ( 
.A1(n_1784),
.A2(n_1715),
.B(n_1826),
.C(n_1708),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1837),
.B(n_1024),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1833),
.A2(n_1024),
.B(n_603),
.Y(n_1910)
);

OAI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1688),
.A2(n_1778),
.B(n_1677),
.Y(n_1911)
);

O2A1O1Ixp33_ASAP7_75t_L g1912 ( 
.A1(n_1715),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1744),
.B(n_17),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1736),
.B(n_18),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1755),
.A2(n_1024),
.B1(n_21),
.B2(n_19),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1758),
.A2(n_22),
.B1(n_19),
.B2(n_20),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_SL g1917 ( 
.A(n_1837),
.B(n_20),
.Y(n_1917)
);

AOI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1845),
.A2(n_589),
.B(n_586),
.Y(n_1918)
);

OAI21xp5_ASAP7_75t_L g1919 ( 
.A1(n_1784),
.A2(n_22),
.B(n_23),
.Y(n_1919)
);

AOI33xp33_ASAP7_75t_L g1920 ( 
.A1(n_1707),
.A2(n_26),
.A3(n_28),
.B1(n_24),
.B2(n_25),
.B3(n_27),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1726),
.B(n_24),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1783),
.Y(n_1922)
);

AOI21xp5_ASAP7_75t_L g1923 ( 
.A1(n_1845),
.A2(n_599),
.B(n_598),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1809),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1749),
.A2(n_602),
.B(n_600),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1681),
.A2(n_27),
.B1(n_25),
.B2(n_26),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1728),
.B(n_495),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1729),
.B(n_1733),
.Y(n_1928)
);

INVx4_ASAP7_75t_L g1929 ( 
.A(n_1809),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1749),
.A2(n_609),
.B(n_498),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1687),
.Y(n_1931)
);

O2A1O1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1680),
.A2(n_1710),
.B(n_1724),
.C(n_1765),
.Y(n_1932)
);

INVx6_ASAP7_75t_L g1933 ( 
.A(n_1811),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1782),
.B(n_28),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1670),
.A2(n_580),
.B(n_579),
.Y(n_1935)
);

O2A1O1Ixp33_ASAP7_75t_L g1936 ( 
.A1(n_1680),
.A2(n_32),
.B(n_29),
.C(n_30),
.Y(n_1936)
);

AO22x1_ASAP7_75t_L g1937 ( 
.A1(n_1804),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_1937)
);

INVx4_ASAP7_75t_L g1938 ( 
.A(n_1685),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1843),
.A2(n_1849),
.B(n_1815),
.Y(n_1939)
);

NOR2x1_ASAP7_75t_L g1940 ( 
.A(n_1719),
.B(n_497),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1850),
.B(n_34),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1698),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_SL g1943 ( 
.A(n_1848),
.B(n_34),
.Y(n_1943)
);

NOR2xp67_ASAP7_75t_L g1944 ( 
.A(n_1769),
.B(n_499),
.Y(n_1944)
);

AND2x4_ASAP7_75t_L g1945 ( 
.A(n_1668),
.B(n_501),
.Y(n_1945)
);

O2A1O1Ixp5_ASAP7_75t_SL g1946 ( 
.A1(n_1720),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1686),
.B(n_35),
.Y(n_1947)
);

AOI21xp5_ASAP7_75t_L g1948 ( 
.A1(n_1674),
.A2(n_608),
.B(n_606),
.Y(n_1948)
);

INVx2_ASAP7_75t_SL g1949 ( 
.A(n_1751),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1710),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_1950)
);

INVx1_ASAP7_75t_SL g1951 ( 
.A(n_1779),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1678),
.A2(n_605),
.B(n_503),
.Y(n_1952)
);

XOR2xp5_ASAP7_75t_L g1953 ( 
.A(n_1772),
.B(n_502),
.Y(n_1953)
);

A2O1A1Ixp33_ASAP7_75t_L g1954 ( 
.A1(n_1676),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_1954)
);

O2A1O1Ixp33_ASAP7_75t_L g1955 ( 
.A1(n_1745),
.A2(n_43),
.B(n_40),
.C(n_42),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1703),
.Y(n_1956)
);

AND2x6_ASAP7_75t_L g1957 ( 
.A(n_1668),
.B(n_505),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1725),
.B(n_42),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1716),
.B(n_43),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1706),
.B(n_44),
.Y(n_1960)
);

AOI21xp5_ASAP7_75t_L g1961 ( 
.A1(n_1669),
.A2(n_507),
.B(n_506),
.Y(n_1961)
);

AND2x4_ASAP7_75t_L g1962 ( 
.A(n_1737),
.B(n_508),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1756),
.B(n_1742),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1754),
.B(n_44),
.Y(n_1964)
);

NOR3xp33_ASAP7_75t_L g1965 ( 
.A(n_1745),
.B(n_45),
.C(n_46),
.Y(n_1965)
);

NAND2xp33_ASAP7_75t_L g1966 ( 
.A(n_1672),
.B(n_45),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1780),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1967)
);

NOR2x1_ASAP7_75t_L g1968 ( 
.A(n_1802),
.B(n_1800),
.Y(n_1968)
);

AOI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1676),
.A2(n_604),
.B(n_513),
.Y(n_1969)
);

NOR2xp33_ASAP7_75t_L g1970 ( 
.A(n_1746),
.B(n_510),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1774),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1738),
.B(n_514),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1777),
.B(n_52),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1770),
.Y(n_1974)
);

OAI21xp5_ASAP7_75t_L g1975 ( 
.A1(n_1689),
.A2(n_53),
.B(n_54),
.Y(n_1975)
);

O2A1O1Ixp33_ASAP7_75t_L g1976 ( 
.A1(n_1712),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1788),
.Y(n_1977)
);

AOI22xp5_ASAP7_75t_L g1978 ( 
.A1(n_1730),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_1978)
);

CKINVDCx8_ASAP7_75t_R g1979 ( 
.A(n_1727),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1794),
.B(n_58),
.Y(n_1980)
);

OAI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1757),
.A2(n_1761),
.B1(n_1767),
.B2(n_1763),
.Y(n_1981)
);

BUFx2_ASAP7_75t_L g1982 ( 
.A(n_1770),
.Y(n_1982)
);

BUFx12f_ASAP7_75t_L g1983 ( 
.A(n_1810),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1830),
.B(n_58),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1816),
.B(n_59),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1709),
.B(n_516),
.Y(n_1986)
);

A2O1A1Ixp33_ASAP7_75t_L g1987 ( 
.A1(n_1805),
.A2(n_62),
.B(n_59),
.C(n_60),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1819),
.A2(n_63),
.B(n_60),
.C(n_62),
.Y(n_1988)
);

INVx1_ASAP7_75t_SL g1989 ( 
.A(n_1690),
.Y(n_1989)
);

OAI22xp5_ASAP7_75t_SL g1990 ( 
.A1(n_1766),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1820),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1832),
.B(n_65),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1732),
.A2(n_518),
.B(n_517),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1818),
.A2(n_68),
.B(n_66),
.C(n_67),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1705),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1827),
.B(n_66),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1836),
.B(n_67),
.Y(n_1997)
);

CKINVDCx8_ASAP7_75t_R g1998 ( 
.A(n_1727),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1734),
.A2(n_521),
.B(n_520),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1840),
.A2(n_1775),
.B1(n_1807),
.B2(n_1801),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1808),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1821),
.A2(n_523),
.B(n_522),
.Y(n_2002)
);

NOR2xp67_ASAP7_75t_L g2003 ( 
.A(n_1813),
.B(n_524),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1814),
.B(n_68),
.Y(n_2004)
);

AOI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1823),
.A2(n_529),
.B(n_528),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1817),
.B(n_1825),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1824),
.A2(n_72),
.B1(n_69),
.B2(n_70),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1828),
.A2(n_531),
.B(n_530),
.Y(n_2008)
);

NOR2xp33_ASAP7_75t_L g2009 ( 
.A(n_1839),
.B(n_533),
.Y(n_2009)
);

O2A1O1Ixp33_ASAP7_75t_L g2010 ( 
.A1(n_1720),
.A2(n_72),
.B(n_69),
.C(n_70),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1776),
.B(n_73),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1727),
.B(n_74),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_R g2013 ( 
.A(n_1727),
.B(n_534),
.Y(n_2013)
);

BUFx2_ASAP7_75t_L g2014 ( 
.A(n_1672),
.Y(n_2014)
);

AO22x1_ASAP7_75t_L g2015 ( 
.A1(n_1672),
.A2(n_78),
.B1(n_75),
.B2(n_77),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1672),
.B(n_1750),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1831),
.A2(n_596),
.B(n_536),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1748),
.B(n_77),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1679),
.B(n_79),
.Y(n_2019)
);

CKINVDCx11_ASAP7_75t_R g2020 ( 
.A(n_1735),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1835),
.A2(n_537),
.B(n_535),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1721),
.B(n_538),
.Y(n_2022)
);

NOR2xp33_ASAP7_75t_L g2023 ( 
.A(n_1679),
.B(n_540),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1907),
.B(n_1838),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1869),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1859),
.A2(n_1760),
.B1(n_1847),
.B2(n_1846),
.C(n_1844),
.Y(n_2026)
);

INVx2_ASAP7_75t_SL g2027 ( 
.A(n_1881),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1928),
.B(n_79),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1854),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1898),
.B(n_80),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1855),
.A2(n_1768),
.B1(n_1764),
.B2(n_1789),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1903),
.B(n_541),
.Y(n_2032)
);

A2O1A1Ixp33_ASAP7_75t_L g2033 ( 
.A1(n_1932),
.A2(n_1771),
.B(n_1753),
.C(n_1739),
.Y(n_2033)
);

A2O1A1Ixp33_ASAP7_75t_L g2034 ( 
.A1(n_1908),
.A2(n_1692),
.B(n_1697),
.C(n_1704),
.Y(n_2034)
);

INVx3_ASAP7_75t_L g2035 ( 
.A(n_1873),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1852),
.A2(n_1700),
.B1(n_1684),
.B2(n_1812),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1882),
.B(n_1781),
.Y(n_2037)
);

AOI21xp5_ASAP7_75t_L g2038 ( 
.A1(n_1911),
.A2(n_1795),
.B(n_1797),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1894),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1875),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2001),
.B(n_80),
.Y(n_2041)
);

OAI22xp5_ASAP7_75t_SL g2042 ( 
.A1(n_1990),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_1870),
.B(n_542),
.Y(n_2043)
);

OA21x2_ASAP7_75t_L g2044 ( 
.A1(n_1874),
.A2(n_1793),
.B(n_81),
.Y(n_2044)
);

OAI21x1_ASAP7_75t_L g2045 ( 
.A1(n_1878),
.A2(n_546),
.B(n_543),
.Y(n_2045)
);

AOI21xp5_ASAP7_75t_L g2046 ( 
.A1(n_1966),
.A2(n_548),
.B(n_547),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2006),
.B(n_83),
.Y(n_2047)
);

INVx2_ASAP7_75t_SL g2048 ( 
.A(n_1881),
.Y(n_2048)
);

INVx1_ASAP7_75t_SL g2049 ( 
.A(n_1989),
.Y(n_2049)
);

OAI21x1_ASAP7_75t_L g2050 ( 
.A1(n_1865),
.A2(n_551),
.B(n_549),
.Y(n_2050)
);

NOR2xp67_ASAP7_75t_L g2051 ( 
.A(n_2000),
.B(n_552),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1910),
.A2(n_560),
.B(n_555),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1995),
.B(n_85),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1888),
.Y(n_2054)
);

OAI21x1_ASAP7_75t_L g2055 ( 
.A1(n_1961),
.A2(n_1892),
.B(n_1880),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1981),
.B(n_86),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1871),
.B(n_87),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_1873),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1969),
.A2(n_563),
.B(n_562),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1873),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1889),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1896),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1866),
.A2(n_566),
.B(n_565),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_L g2064 ( 
.A1(n_1905),
.A2(n_568),
.B(n_567),
.Y(n_2064)
);

NAND2xp33_ASAP7_75t_L g2065 ( 
.A(n_1919),
.B(n_87),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1920),
.B(n_89),
.Y(n_2066)
);

OAI21x1_ASAP7_75t_L g2067 ( 
.A1(n_1906),
.A2(n_570),
.B(n_569),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1968),
.B(n_572),
.Y(n_2068)
);

AO22x2_ASAP7_75t_L g2069 ( 
.A1(n_1965),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1939),
.A2(n_575),
.B(n_574),
.Y(n_2070)
);

INVx3_ASAP7_75t_L g2071 ( 
.A(n_1904),
.Y(n_2071)
);

OAI21x1_ASAP7_75t_L g2072 ( 
.A1(n_1877),
.A2(n_577),
.B(n_576),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1883),
.B(n_581),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1963),
.B(n_90),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1901),
.B(n_582),
.Y(n_2075)
);

OAI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1948),
.A2(n_584),
.B(n_583),
.Y(n_2076)
);

OAI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1925),
.A2(n_91),
.B(n_92),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1978),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1930),
.A2(n_591),
.B(n_585),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1853),
.B(n_93),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1931),
.B(n_94),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_1952),
.A2(n_1999),
.B(n_1993),
.Y(n_2082)
);

OAI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_1935),
.A2(n_95),
.B(n_96),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_1996),
.B(n_95),
.Y(n_2084)
);

O2A1O1Ixp5_ASAP7_75t_L g2085 ( 
.A1(n_1975),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_1909),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_2086)
);

INVx1_ASAP7_75t_SL g2087 ( 
.A(n_1899),
.Y(n_2087)
);

INVx1_ASAP7_75t_SL g2088 ( 
.A(n_1922),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1933),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1942),
.B(n_100),
.Y(n_2090)
);

AOI21xp5_ASAP7_75t_L g2091 ( 
.A1(n_1918),
.A2(n_594),
.B(n_100),
.Y(n_2091)
);

OAI21x1_ASAP7_75t_L g2092 ( 
.A1(n_2002),
.A2(n_101),
.B(n_102),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1986),
.B(n_101),
.Y(n_2093)
);

AND2x4_ASAP7_75t_SL g2094 ( 
.A(n_1876),
.B(n_102),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1956),
.Y(n_2095)
);

AND3x4_ASAP7_75t_L g2096 ( 
.A(n_1962),
.B(n_103),
.C(n_104),
.Y(n_2096)
);

OA22x2_ASAP7_75t_L g2097 ( 
.A1(n_1917),
.A2(n_106),
.B1(n_103),
.B2(n_105),
.Y(n_2097)
);

BUFx10_ASAP7_75t_L g2098 ( 
.A(n_1933),
.Y(n_2098)
);

AO21x1_ASAP7_75t_L g2099 ( 
.A1(n_1912),
.A2(n_106),
.B(n_107),
.Y(n_2099)
);

OAI21x1_ASAP7_75t_L g2100 ( 
.A1(n_2005),
.A2(n_107),
.B(n_108),
.Y(n_2100)
);

INVx2_ASAP7_75t_L g2101 ( 
.A(n_1977),
.Y(n_2101)
);

BUFx4_ASAP7_75t_SL g2102 ( 
.A(n_1974),
.Y(n_2102)
);

BUFx6f_ASAP7_75t_L g2103 ( 
.A(n_1904),
.Y(n_2103)
);

AOI21xp5_ASAP7_75t_L g2104 ( 
.A1(n_1923),
.A2(n_109),
.B(n_110),
.Y(n_2104)
);

AOI221xp5_ASAP7_75t_L g2105 ( 
.A1(n_1936),
.A2(n_2010),
.B1(n_1955),
.B2(n_1971),
.C(n_1915),
.Y(n_2105)
);

OAI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_1954),
.A2(n_109),
.B(n_111),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1991),
.B(n_482),
.Y(n_2107)
);

INVx3_ASAP7_75t_L g2108 ( 
.A(n_1904),
.Y(n_2108)
);

NAND3xp33_ASAP7_75t_L g2109 ( 
.A(n_1916),
.B(n_112),
.C(n_113),
.Y(n_2109)
);

AO21x1_ASAP7_75t_L g2110 ( 
.A1(n_2018),
.A2(n_113),
.B(n_116),
.Y(n_2110)
);

AO31x2_ASAP7_75t_L g2111 ( 
.A1(n_1868),
.A2(n_118),
.A3(n_116),
.B(n_117),
.Y(n_2111)
);

AO31x2_ASAP7_75t_L g2112 ( 
.A1(n_1886),
.A2(n_119),
.A3(n_117),
.B(n_118),
.Y(n_2112)
);

BUFx6f_ASAP7_75t_L g2113 ( 
.A(n_1982),
.Y(n_2113)
);

INVx1_ASAP7_75t_SL g2114 ( 
.A(n_1890),
.Y(n_2114)
);

AOI21x1_ASAP7_75t_L g2115 ( 
.A1(n_1861),
.A2(n_120),
.B(n_121),
.Y(n_2115)
);

OAI21x1_ASAP7_75t_L g2116 ( 
.A1(n_2008),
.A2(n_122),
.B(n_124),
.Y(n_2116)
);

OAI21x1_ASAP7_75t_L g2117 ( 
.A1(n_2017),
.A2(n_122),
.B(n_125),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_L g2118 ( 
.A1(n_2021),
.A2(n_125),
.B(n_127),
.Y(n_2118)
);

AOI21x1_ASAP7_75t_L g2119 ( 
.A1(n_1891),
.A2(n_127),
.B(n_128),
.Y(n_2119)
);

AOI21xp5_ASAP7_75t_L g2120 ( 
.A1(n_1857),
.A2(n_129),
.B(n_130),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1959),
.B(n_481),
.Y(n_2121)
);

OAI21x1_ASAP7_75t_L g2122 ( 
.A1(n_1867),
.A2(n_129),
.B(n_130),
.Y(n_2122)
);

NOR4xp25_ASAP7_75t_L g2123 ( 
.A(n_1987),
.B(n_1976),
.C(n_1988),
.D(n_1994),
.Y(n_2123)
);

AND2x4_ASAP7_75t_L g2124 ( 
.A(n_2014),
.B(n_131),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1973),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1985),
.Y(n_2126)
);

BUFx10_ASAP7_75t_L g2127 ( 
.A(n_1858),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1941),
.B(n_481),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_L g2129 ( 
.A1(n_1887),
.A2(n_131),
.B(n_133),
.Y(n_2129)
);

INVxp67_ASAP7_75t_SL g2130 ( 
.A(n_1895),
.Y(n_2130)
);

OAI21x1_ASAP7_75t_L g2131 ( 
.A1(n_1862),
.A2(n_134),
.B(n_135),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1934),
.B(n_134),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1921),
.B(n_480),
.Y(n_2133)
);

OAI21x1_ASAP7_75t_L g2134 ( 
.A1(n_1946),
.A2(n_135),
.B(n_136),
.Y(n_2134)
);

INVx1_ASAP7_75t_SL g2135 ( 
.A(n_1951),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_1860),
.A2(n_136),
.B(n_137),
.Y(n_2136)
);

AOI21xp5_ASAP7_75t_L g2137 ( 
.A1(n_2016),
.A2(n_137),
.B(n_138),
.Y(n_2137)
);

AOI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_1872),
.A2(n_138),
.B(n_139),
.Y(n_2138)
);

OAI21x1_ASAP7_75t_SL g2139 ( 
.A1(n_1856),
.A2(n_140),
.B(n_141),
.Y(n_2139)
);

OAI321xp33_ASAP7_75t_L g2140 ( 
.A1(n_2077),
.A2(n_1950),
.A3(n_2007),
.B1(n_1967),
.B2(n_1970),
.C(n_1926),
.Y(n_2140)
);

AOI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_2065),
.A2(n_2015),
.B(n_2019),
.Y(n_2141)
);

A2O1A1Ixp33_ASAP7_75t_L g2142 ( 
.A1(n_2077),
.A2(n_1927),
.B(n_2009),
.C(n_1884),
.Y(n_2142)
);

BUFx2_ASAP7_75t_L g2143 ( 
.A(n_2025),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2061),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2049),
.B(n_1914),
.Y(n_2145)
);

OAI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_2104),
.A2(n_1943),
.B(n_1984),
.Y(n_2146)
);

NOR2xp67_ASAP7_75t_SL g2147 ( 
.A(n_2109),
.B(n_1979),
.Y(n_2147)
);

INVx3_ASAP7_75t_SL g2148 ( 
.A(n_2098),
.Y(n_2148)
);

BUFx3_ASAP7_75t_L g2149 ( 
.A(n_2098),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2087),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2056),
.B(n_1937),
.C(n_1992),
.Y(n_2151)
);

NOR2xp33_ASAP7_75t_L g2152 ( 
.A(n_2127),
.B(n_1863),
.Y(n_2152)
);

AOI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_2083),
.A2(n_2022),
.B(n_2023),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2126),
.B(n_1913),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2087),
.B(n_1885),
.Y(n_2155)
);

NAND2x1_ASAP7_75t_L g2156 ( 
.A(n_2095),
.B(n_2101),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2088),
.Y(n_2157)
);

OAI22xp5_ASAP7_75t_L g2158 ( 
.A1(n_2078),
.A2(n_1998),
.B1(n_1997),
.B2(n_2004),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_SL g2159 ( 
.A(n_2049),
.B(n_2013),
.Y(n_2159)
);

AOI22xp5_ASAP7_75t_L g2160 ( 
.A1(n_2042),
.A2(n_2011),
.B1(n_1947),
.B2(n_1964),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2029),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2088),
.Y(n_2162)
);

INVx2_ASAP7_75t_SL g2163 ( 
.A(n_2102),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_2038),
.A2(n_2022),
.B(n_1940),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2040),
.B(n_2054),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_2046),
.A2(n_2051),
.B(n_2082),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2125),
.B(n_1960),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2039),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2114),
.B(n_1980),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2114),
.B(n_2012),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2062),
.Y(n_2171)
);

A2O1A1Ixp33_ASAP7_75t_L g2172 ( 
.A1(n_2106),
.A2(n_2003),
.B(n_1944),
.C(n_1902),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_2058),
.Y(n_2173)
);

INVx3_ASAP7_75t_SL g2174 ( 
.A(n_2127),
.Y(n_2174)
);

A2O1A1Ixp33_ASAP7_75t_SL g2175 ( 
.A1(n_2136),
.A2(n_1864),
.B(n_1924),
.C(n_1879),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_2113),
.Y(n_2176)
);

BUFx3_ASAP7_75t_L g2177 ( 
.A(n_2027),
.Y(n_2177)
);

AOI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_2042),
.A2(n_1958),
.B1(n_1972),
.B2(n_1962),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2111),
.Y(n_2179)
);

AOI22xp5_ASAP7_75t_L g2180 ( 
.A1(n_2078),
.A2(n_1972),
.B1(n_1893),
.B2(n_1953),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_2051),
.A2(n_2052),
.B(n_2059),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_2120),
.A2(n_1945),
.B(n_1897),
.Y(n_2182)
);

INVx1_ASAP7_75t_SL g2183 ( 
.A(n_2135),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2113),
.B(n_1885),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2035),
.Y(n_2185)
);

AOI21xp5_ASAP7_75t_L g2186 ( 
.A1(n_2091),
.A2(n_1945),
.B(n_1893),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2079),
.A2(n_1879),
.B(n_1864),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2111),
.Y(n_2188)
);

O2A1O1Ixp5_ASAP7_75t_L g2189 ( 
.A1(n_2106),
.A2(n_1924),
.B(n_1929),
.C(n_1876),
.Y(n_2189)
);

INVx3_ASAP7_75t_SL g2190 ( 
.A(n_2113),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2135),
.B(n_1949),
.Y(n_2191)
);

A2O1A1Ixp33_ASAP7_75t_SL g2192 ( 
.A1(n_2138),
.A2(n_1957),
.B(n_1851),
.C(n_1900),
.Y(n_2192)
);

CKINVDCx6p67_ASAP7_75t_R g2193 ( 
.A(n_2058),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2028),
.B(n_1957),
.Y(n_2194)
);

BUFx4_ASAP7_75t_SL g2195 ( 
.A(n_2084),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2024),
.B(n_1957),
.Y(n_2196)
);

BUFx2_ASAP7_75t_L g2197 ( 
.A(n_2035),
.Y(n_2197)
);

BUFx2_ASAP7_75t_SL g2198 ( 
.A(n_2048),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2060),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2111),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2032),
.B(n_1983),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_2060),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2057),
.B(n_1957),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2080),
.B(n_1938),
.Y(n_2204)
);

BUFx6f_ASAP7_75t_L g2205 ( 
.A(n_2058),
.Y(n_2205)
);

NAND2xp33_ASAP7_75t_L g2206 ( 
.A(n_2109),
.B(n_2020),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_R g2207 ( 
.A(n_2089),
.B(n_1929),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2047),
.B(n_1938),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2093),
.B(n_140),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_2130),
.B(n_141),
.Y(n_2210)
);

NAND2xp33_ASAP7_75t_L g2211 ( 
.A(n_2066),
.B(n_142),
.Y(n_2211)
);

BUFx6f_ASAP7_75t_L g2212 ( 
.A(n_2103),
.Y(n_2212)
);

A2O1A1Ixp33_ASAP7_75t_L g2213 ( 
.A1(n_2105),
.A2(n_144),
.B(n_142),
.C(n_143),
.Y(n_2213)
);

AOI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_2037),
.A2(n_2031),
.B(n_2036),
.Y(n_2214)
);

OA21x2_ASAP7_75t_L g2215 ( 
.A1(n_2072),
.A2(n_143),
.B(n_144),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_2071),
.Y(n_2216)
);

OR2x6_ASAP7_75t_L g2217 ( 
.A(n_2073),
.B(n_145),
.Y(n_2217)
);

AOI21xp5_ASAP7_75t_L g2218 ( 
.A1(n_2055),
.A2(n_145),
.B(n_147),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_2148),
.Y(n_2219)
);

AOI22xp33_ASAP7_75t_L g2220 ( 
.A1(n_2206),
.A2(n_2099),
.B1(n_2069),
.B2(n_2110),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2150),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_L g2222 ( 
.A1(n_2142),
.A2(n_2096),
.B1(n_2069),
.B2(n_2097),
.Y(n_2222)
);

AOI22xp33_ASAP7_75t_SL g2223 ( 
.A1(n_2158),
.A2(n_2139),
.B1(n_2137),
.B2(n_2122),
.Y(n_2223)
);

AOI22xp33_ASAP7_75t_L g2224 ( 
.A1(n_2211),
.A2(n_2132),
.B1(n_2133),
.B2(n_2121),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_SL g2225 ( 
.A1(n_2151),
.A2(n_2131),
.B1(n_2043),
.B2(n_2086),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_2156),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2161),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2180),
.A2(n_2124),
.B1(n_2128),
.B2(n_2075),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2170),
.B(n_2030),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_2185),
.Y(n_2230)
);

CKINVDCx8_ASAP7_75t_R g2231 ( 
.A(n_2198),
.Y(n_2231)
);

OAI22xp33_ASAP7_75t_SL g2232 ( 
.A1(n_2217),
.A2(n_2068),
.B1(n_2115),
.B2(n_2041),
.Y(n_2232)
);

OAI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_2180),
.A2(n_2053),
.B1(n_2119),
.B2(n_2074),
.Y(n_2233)
);

BUFx12f_ASAP7_75t_L g2234 ( 
.A(n_2163),
.Y(n_2234)
);

CKINVDCx11_ASAP7_75t_R g2235 ( 
.A(n_2190),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2144),
.Y(n_2236)
);

CKINVDCx20_ASAP7_75t_R g2237 ( 
.A(n_2174),
.Y(n_2237)
);

AOI22xp33_ASAP7_75t_SL g2238 ( 
.A1(n_2151),
.A2(n_2209),
.B1(n_2141),
.B2(n_2153),
.Y(n_2238)
);

BUFx12f_ASAP7_75t_L g2239 ( 
.A(n_2149),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2165),
.Y(n_2240)
);

INVx2_ASAP7_75t_L g2241 ( 
.A(n_2157),
.Y(n_2241)
);

CKINVDCx5p33_ASAP7_75t_R g2242 ( 
.A(n_2207),
.Y(n_2242)
);

BUFx6f_ASAP7_75t_L g2243 ( 
.A(n_2205),
.Y(n_2243)
);

CKINVDCx5p33_ASAP7_75t_R g2244 ( 
.A(n_2143),
.Y(n_2244)
);

BUFx6f_ASAP7_75t_L g2245 ( 
.A(n_2205),
.Y(n_2245)
);

INVx1_ASAP7_75t_SL g2246 ( 
.A(n_2183),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2183),
.B(n_2081),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_2205),
.Y(n_2248)
);

INVx3_ASAP7_75t_L g2249 ( 
.A(n_2199),
.Y(n_2249)
);

BUFx12f_ASAP7_75t_L g2250 ( 
.A(n_2210),
.Y(n_2250)
);

AOI22xp33_ASAP7_75t_L g2251 ( 
.A1(n_2147),
.A2(n_2124),
.B1(n_2100),
.B2(n_2116),
.Y(n_2251)
);

AOI22xp33_ASAP7_75t_SL g2252 ( 
.A1(n_2146),
.A2(n_2217),
.B1(n_2210),
.B2(n_2186),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2162),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2168),
.Y(n_2254)
);

AOI22xp33_ASAP7_75t_L g2255 ( 
.A1(n_2217),
.A2(n_2092),
.B1(n_2118),
.B2(n_2117),
.Y(n_2255)
);

INVx1_ASAP7_75t_SL g2256 ( 
.A(n_2177),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2171),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2176),
.B(n_2071),
.Y(n_2258)
);

INVx1_ASAP7_75t_SL g2259 ( 
.A(n_2191),
.Y(n_2259)
);

AOI22xp33_ASAP7_75t_SL g2260 ( 
.A1(n_2203),
.A2(n_2094),
.B1(n_2129),
.B2(n_2134),
.Y(n_2260)
);

INVx4_ASAP7_75t_L g2261 ( 
.A(n_2212),
.Y(n_2261)
);

AOI22xp33_ASAP7_75t_SL g2262 ( 
.A1(n_2214),
.A2(n_2085),
.B1(n_2123),
.B2(n_2044),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2160),
.A2(n_2090),
.B1(n_2107),
.B2(n_2026),
.Y(n_2263)
);

BUFx10_ASAP7_75t_L g2264 ( 
.A(n_2201),
.Y(n_2264)
);

AOI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2196),
.A2(n_2076),
.B1(n_2050),
.B2(n_2070),
.Y(n_2265)
);

INVx3_ASAP7_75t_L g2266 ( 
.A(n_2202),
.Y(n_2266)
);

OAI21xp33_ASAP7_75t_SL g2267 ( 
.A1(n_2159),
.A2(n_2194),
.B(n_2160),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2221),
.B(n_2179),
.Y(n_2268)
);

BUFx3_ASAP7_75t_L g2269 ( 
.A(n_2235),
.Y(n_2269)
);

AND2x6_ASAP7_75t_L g2270 ( 
.A(n_2226),
.B(n_2155),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2246),
.B(n_2145),
.Y(n_2271)
);

OR2x6_ASAP7_75t_L g2272 ( 
.A(n_2226),
.B(n_2164),
.Y(n_2272)
);

O2A1O1Ixp5_ASAP7_75t_L g2273 ( 
.A1(n_2222),
.A2(n_2218),
.B(n_2213),
.C(n_2181),
.Y(n_2273)
);

AOI21xp5_ASAP7_75t_L g2274 ( 
.A1(n_2238),
.A2(n_2166),
.B(n_2140),
.Y(n_2274)
);

O2A1O1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_2233),
.A2(n_2192),
.B(n_2172),
.C(n_2175),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2240),
.B(n_2188),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2238),
.A2(n_2178),
.B1(n_2182),
.B2(n_2152),
.Y(n_2277)
);

OAI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2220),
.A2(n_2178),
.B1(n_2204),
.B2(n_2208),
.Y(n_2278)
);

A2O1A1Ixp33_ASAP7_75t_L g2279 ( 
.A1(n_2267),
.A2(n_2252),
.B(n_2224),
.C(n_2189),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2259),
.B(n_2200),
.Y(n_2280)
);

AOI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2262),
.A2(n_2187),
.B(n_2034),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2254),
.Y(n_2282)
);

AND2x2_ASAP7_75t_L g2283 ( 
.A(n_2236),
.B(n_2197),
.Y(n_2283)
);

NOR2x1_ASAP7_75t_SL g2284 ( 
.A(n_2241),
.B(n_2253),
.Y(n_2284)
);

AOI211xp5_ASAP7_75t_L g2285 ( 
.A1(n_2233),
.A2(n_2123),
.B(n_2169),
.C(n_2167),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2257),
.Y(n_2286)
);

AND2x2_ASAP7_75t_L g2287 ( 
.A(n_2258),
.B(n_2154),
.Y(n_2287)
);

AND2x2_ASAP7_75t_L g2288 ( 
.A(n_2227),
.B(n_2155),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2230),
.B(n_2216),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2230),
.B(n_2173),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2249),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2247),
.B(n_2044),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_2249),
.B(n_2173),
.Y(n_2293)
);

O2A1O1Ixp33_ASAP7_75t_L g2294 ( 
.A1(n_2232),
.A2(n_2033),
.B(n_2184),
.C(n_2108),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_2229),
.B(n_2112),
.Y(n_2295)
);

AOI211xp5_ASAP7_75t_SL g2296 ( 
.A1(n_2274),
.A2(n_2228),
.B(n_2237),
.C(n_2252),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2280),
.B(n_2266),
.Y(n_2297)
);

CKINVDCx5p33_ASAP7_75t_R g2298 ( 
.A(n_2269),
.Y(n_2298)
);

BUFx2_ASAP7_75t_L g2299 ( 
.A(n_2272),
.Y(n_2299)
);

CKINVDCx5p33_ASAP7_75t_R g2300 ( 
.A(n_2269),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2284),
.Y(n_2301)
);

BUFx10_ASAP7_75t_L g2302 ( 
.A(n_2272),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2276),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_R g2304 ( 
.A(n_2270),
.B(n_2231),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2276),
.Y(n_2305)
);

INVx3_ASAP7_75t_L g2306 ( 
.A(n_2272),
.Y(n_2306)
);

NOR2xp33_ASAP7_75t_L g2307 ( 
.A(n_2298),
.B(n_2219),
.Y(n_2307)
);

BUFx3_ASAP7_75t_L g2308 ( 
.A(n_2299),
.Y(n_2308)
);

AND2x2_ASAP7_75t_L g2309 ( 
.A(n_2299),
.B(n_2272),
.Y(n_2309)
);

OA21x2_ASAP7_75t_L g2310 ( 
.A1(n_2299),
.A2(n_2281),
.B(n_2279),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2306),
.B(n_2270),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2303),
.Y(n_2312)
);

OA21x2_ASAP7_75t_L g2313 ( 
.A1(n_2301),
.A2(n_2279),
.B(n_2273),
.Y(n_2313)
);

OR2x6_ASAP7_75t_L g2314 ( 
.A(n_2301),
.B(n_2275),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2312),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2312),
.Y(n_2316)
);

NAND2x1p5_ASAP7_75t_L g2317 ( 
.A(n_2310),
.B(n_2306),
.Y(n_2317)
);

AND2x4_ASAP7_75t_SL g2318 ( 
.A(n_2311),
.B(n_2219),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2312),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_2308),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2310),
.B(n_2306),
.Y(n_2321)
);

BUFx2_ASAP7_75t_SL g2322 ( 
.A(n_2308),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2308),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_2308),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_2318),
.Y(n_2325)
);

INVx3_ASAP7_75t_SL g2326 ( 
.A(n_2320),
.Y(n_2326)
);

OAI31xp33_ASAP7_75t_L g2327 ( 
.A1(n_2317),
.A2(n_2296),
.A3(n_2277),
.B(n_2310),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2318),
.B(n_2313),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2315),
.Y(n_2329)
);

INVx3_ASAP7_75t_L g2330 ( 
.A(n_2317),
.Y(n_2330)
);

BUFx2_ASAP7_75t_L g2331 ( 
.A(n_2320),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2324),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2321),
.A2(n_2310),
.B1(n_2313),
.B2(n_2314),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2324),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2322),
.Y(n_2335)
);

OAI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2322),
.A2(n_2310),
.B1(n_2314),
.B2(n_2313),
.Y(n_2336)
);

OR2x2_ASAP7_75t_L g2337 ( 
.A(n_2335),
.B(n_2323),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2330),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2331),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_2330),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2327),
.B(n_2336),
.Y(n_2341)
);

NAND2x1p5_ASAP7_75t_L g2342 ( 
.A(n_2325),
.B(n_2310),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2331),
.Y(n_2343)
);

OR2x2_ASAP7_75t_L g2344 ( 
.A(n_2335),
.B(n_2314),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2330),
.Y(n_2345)
);

INVx1_ASAP7_75t_SL g2346 ( 
.A(n_2344),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2341),
.B(n_2326),
.Y(n_2347)
);

INVx3_ASAP7_75t_L g2348 ( 
.A(n_2340),
.Y(n_2348)
);

OR2x2_ASAP7_75t_L g2349 ( 
.A(n_2337),
.B(n_2326),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2348),
.B(n_2325),
.Y(n_2350)
);

OR2x2_ASAP7_75t_L g2351 ( 
.A(n_2347),
.B(n_2339),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2349),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2346),
.Y(n_2353)
);

AOI32xp33_ASAP7_75t_L g2354 ( 
.A1(n_2350),
.A2(n_2333),
.A3(n_2321),
.B1(n_2343),
.B2(n_2339),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2350),
.Y(n_2355)
);

INVx1_ASAP7_75t_SL g2356 ( 
.A(n_2351),
.Y(n_2356)
);

OAI21xp33_ASAP7_75t_SL g2357 ( 
.A1(n_2353),
.A2(n_2328),
.B(n_2343),
.Y(n_2357)
);

AOI222xp33_ASAP7_75t_L g2358 ( 
.A1(n_2352),
.A2(n_2326),
.B1(n_2334),
.B2(n_2330),
.C1(n_2328),
.C2(n_2329),
.Y(n_2358)
);

NAND3xp33_ASAP7_75t_L g2359 ( 
.A(n_2350),
.B(n_2345),
.C(n_2338),
.Y(n_2359)
);

AO21x2_ASAP7_75t_L g2360 ( 
.A1(n_2355),
.A2(n_2329),
.B(n_2319),
.Y(n_2360)
);

OR2x2_ASAP7_75t_L g2361 ( 
.A(n_2356),
.B(n_2334),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2359),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_2358),
.Y(n_2363)
);

NOR2xp33_ASAP7_75t_L g2364 ( 
.A(n_2357),
.B(n_2300),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2354),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2355),
.B(n_2332),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_2355),
.B(n_2342),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2355),
.B(n_2332),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2355),
.B(n_2307),
.Y(n_2369)
);

A2O1A1Ixp33_ASAP7_75t_L g2370 ( 
.A1(n_2365),
.A2(n_2340),
.B(n_2332),
.C(n_2296),
.Y(n_2370)
);

OAI211xp5_ASAP7_75t_SL g2371 ( 
.A1(n_2365),
.A2(n_2332),
.B(n_2307),
.C(n_2285),
.Y(n_2371)
);

OAI21xp5_ASAP7_75t_SL g2372 ( 
.A1(n_2364),
.A2(n_2309),
.B(n_2219),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2369),
.B(n_2234),
.Y(n_2373)
);

AOI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2363),
.A2(n_2314),
.B1(n_2313),
.B2(n_2309),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2361),
.Y(n_2375)
);

HB1xp67_ASAP7_75t_L g2376 ( 
.A(n_2360),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2368),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2366),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2367),
.B(n_2314),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2362),
.A2(n_2314),
.B(n_2313),
.Y(n_2380)
);

INVx2_ASAP7_75t_SL g2381 ( 
.A(n_2360),
.Y(n_2381)
);

INVx1_ASAP7_75t_SL g2382 ( 
.A(n_2361),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2376),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2381),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2375),
.Y(n_2385)
);

AOI221xp5_ASAP7_75t_L g2386 ( 
.A1(n_2370),
.A2(n_2316),
.B1(n_2309),
.B2(n_2306),
.C(n_2219),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2382),
.B(n_2314),
.Y(n_2387)
);

OR2x2_ASAP7_75t_L g2388 ( 
.A(n_2377),
.B(n_2314),
.Y(n_2388)
);

OAI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2374),
.A2(n_2313),
.B1(n_2306),
.B2(n_2301),
.Y(n_2389)
);

XNOR2xp5_ASAP7_75t_L g2390 ( 
.A(n_2379),
.B(n_2242),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2378),
.Y(n_2391)
);

AOI21xp33_ASAP7_75t_L g2392 ( 
.A1(n_2373),
.A2(n_2372),
.B(n_2371),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2380),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_2380),
.A2(n_2309),
.B1(n_2311),
.B2(n_2239),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2376),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2371),
.A2(n_2311),
.B1(n_2302),
.B2(n_2264),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2382),
.B(n_2256),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2393),
.Y(n_2398)
);

OR2x2_ASAP7_75t_L g2399 ( 
.A(n_2397),
.B(n_2388),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_2384),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2385),
.B(n_2244),
.Y(n_2401)
);

HB1xp67_ASAP7_75t_L g2402 ( 
.A(n_2387),
.Y(n_2402)
);

NOR2xp33_ASAP7_75t_L g2403 ( 
.A(n_2390),
.B(n_2392),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_SL g2404 ( 
.A(n_2389),
.B(n_2311),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2383),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_L g2406 ( 
.A(n_2394),
.B(n_2311),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2395),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2391),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2386),
.B(n_2311),
.Y(n_2409)
);

OAI222xp33_ASAP7_75t_L g2410 ( 
.A1(n_2396),
.A2(n_2224),
.B1(n_2223),
.B2(n_2225),
.C1(n_2278),
.C2(n_2262),
.Y(n_2410)
);

AOI22xp5_ASAP7_75t_L g2411 ( 
.A1(n_2396),
.A2(n_2264),
.B1(n_2302),
.B2(n_2250),
.Y(n_2411)
);

O2A1O1Ixp5_ASAP7_75t_L g2412 ( 
.A1(n_2404),
.A2(n_2400),
.B(n_2398),
.C(n_2405),
.Y(n_2412)
);

OAI211xp5_ASAP7_75t_L g2413 ( 
.A1(n_2403),
.A2(n_2304),
.B(n_2223),
.C(n_2225),
.Y(n_2413)
);

NOR3xp33_ASAP7_75t_L g2414 ( 
.A(n_2402),
.B(n_2195),
.C(n_2294),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2401),
.B(n_2271),
.Y(n_2415)
);

NOR3xp33_ASAP7_75t_L g2416 ( 
.A(n_2399),
.B(n_2260),
.C(n_2295),
.Y(n_2416)
);

INVx1_ASAP7_75t_SL g2417 ( 
.A(n_2408),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2407),
.B(n_2302),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2411),
.B(n_2302),
.Y(n_2419)
);

NOR4xp25_ASAP7_75t_L g2420 ( 
.A(n_2406),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2409),
.B(n_2302),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_L g2422 ( 
.A(n_2410),
.B(n_2282),
.Y(n_2422)
);

AND4x1_ASAP7_75t_L g2423 ( 
.A(n_2403),
.B(n_2263),
.C(n_150),
.D(n_148),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_2400),
.Y(n_2424)
);

OA22x2_ASAP7_75t_L g2425 ( 
.A1(n_2411),
.A2(n_2303),
.B1(n_2305),
.B2(n_2261),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2401),
.Y(n_2426)
);

NOR3xp33_ASAP7_75t_L g2427 ( 
.A(n_2403),
.B(n_2260),
.C(n_149),
.Y(n_2427)
);

AOI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2401),
.A2(n_2263),
.B(n_2292),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2401),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_2400),
.B(n_2297),
.Y(n_2430)
);

NAND4xp25_ASAP7_75t_L g2431 ( 
.A(n_2403),
.B(n_2251),
.C(n_2255),
.D(n_2292),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2401),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2401),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2420),
.B(n_151),
.Y(n_2434)
);

OAI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_2424),
.A2(n_2305),
.B1(n_2297),
.B2(n_2193),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2423),
.B(n_151),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2417),
.B(n_152),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2430),
.B(n_2418),
.Y(n_2438)
);

AOI321xp33_ASAP7_75t_L g2439 ( 
.A1(n_2419),
.A2(n_2251),
.A3(n_2184),
.B1(n_154),
.B2(n_156),
.C(n_152),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2421),
.B(n_153),
.Y(n_2440)
);

AOI31xp67_ASAP7_75t_SL g2441 ( 
.A1(n_2422),
.A2(n_2304),
.A3(n_155),
.B(n_153),
.Y(n_2441)
);

OAI211xp5_ASAP7_75t_SL g2442 ( 
.A1(n_2412),
.A2(n_157),
.B(n_154),
.C(n_155),
.Y(n_2442)
);

NAND3xp33_ASAP7_75t_L g2443 ( 
.A(n_2426),
.B(n_158),
.C(n_159),
.Y(n_2443)
);

NOR2x1_ASAP7_75t_L g2444 ( 
.A(n_2429),
.B(n_158),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2414),
.B(n_159),
.Y(n_2445)
);

NOR2x1_ASAP7_75t_L g2446 ( 
.A(n_2432),
.B(n_160),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2415),
.B(n_2433),
.Y(n_2447)
);

NOR2xp33_ASAP7_75t_L g2448 ( 
.A(n_2425),
.B(n_160),
.Y(n_2448)
);

NAND4xp25_ASAP7_75t_SL g2449 ( 
.A(n_2427),
.B(n_2297),
.C(n_2280),
.D(n_2291),
.Y(n_2449)
);

INVxp67_ASAP7_75t_SL g2450 ( 
.A(n_2428),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2416),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_SL g2452 ( 
.A(n_2413),
.B(n_2103),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2431),
.Y(n_2453)
);

INVxp67_ASAP7_75t_L g2454 ( 
.A(n_2418),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2419),
.A2(n_161),
.B(n_162),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2424),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2430),
.Y(n_2457)
);

NOR3x1_ASAP7_75t_L g2458 ( 
.A(n_2424),
.B(n_161),
.C(n_162),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2430),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2430),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2430),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_2420),
.B(n_163),
.Y(n_2462)
);

OR2x2_ASAP7_75t_L g2463 ( 
.A(n_2420),
.B(n_163),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2420),
.B(n_2103),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2420),
.B(n_164),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2420),
.B(n_164),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2430),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2424),
.B(n_165),
.Y(n_2468)
);

AOI221xp5_ASAP7_75t_L g2469 ( 
.A1(n_2420),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.C(n_168),
.Y(n_2469)
);

NOR4xp25_ASAP7_75t_L g2470 ( 
.A(n_2417),
.B(n_170),
.C(n_166),
.D(n_169),
.Y(n_2470)
);

AOI311xp33_ASAP7_75t_L g2471 ( 
.A1(n_2440),
.A2(n_2451),
.A3(n_2448),
.B(n_2453),
.C(n_2457),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_L g2472 ( 
.A(n_2468),
.B(n_170),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_SL g2473 ( 
.A(n_2436),
.B(n_2261),
.Y(n_2473)
);

NAND4xp25_ASAP7_75t_L g2474 ( 
.A(n_2439),
.B(n_173),
.C(n_171),
.D(n_172),
.Y(n_2474)
);

NOR3xp33_ASAP7_75t_L g2475 ( 
.A(n_2445),
.B(n_171),
.C(n_172),
.Y(n_2475)
);

NAND3xp33_ASAP7_75t_SL g2476 ( 
.A(n_2469),
.B(n_174),
.C(n_175),
.Y(n_2476)
);

AOI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2456),
.A2(n_2449),
.B1(n_2442),
.B2(n_2450),
.Y(n_2477)
);

INVxp67_ASAP7_75t_L g2478 ( 
.A(n_2444),
.Y(n_2478)
);

AOI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2459),
.A2(n_2270),
.B1(n_2283),
.B2(n_2245),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2463),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2434),
.Y(n_2481)
);

NAND2xp5_ASAP7_75t_L g2482 ( 
.A(n_2470),
.B(n_175),
.Y(n_2482)
);

NOR2x1_ASAP7_75t_L g2483 ( 
.A(n_2446),
.B(n_176),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2470),
.B(n_177),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2458),
.B(n_177),
.Y(n_2485)
);

O2A1O1Ixp33_ASAP7_75t_L g2486 ( 
.A1(n_2462),
.A2(n_181),
.B(n_178),
.C(n_179),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2465),
.B(n_178),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2466),
.Y(n_2488)
);

INVxp67_ASAP7_75t_L g2489 ( 
.A(n_2437),
.Y(n_2489)
);

OAI322xp33_ASAP7_75t_L g2490 ( 
.A1(n_2452),
.A2(n_179),
.A3(n_181),
.B1(n_182),
.B2(n_183),
.C1(n_184),
.C2(n_185),
.Y(n_2490)
);

NAND3xp33_ASAP7_75t_L g2491 ( 
.A(n_2455),
.B(n_182),
.C(n_184),
.Y(n_2491)
);

NOR2x1_ASAP7_75t_L g2492 ( 
.A(n_2443),
.B(n_185),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2464),
.Y(n_2493)
);

NAND3xp33_ASAP7_75t_L g2494 ( 
.A(n_2460),
.B(n_186),
.C(n_187),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2461),
.B(n_188),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2467),
.B(n_188),
.Y(n_2496)
);

NOR3x1_ASAP7_75t_L g2497 ( 
.A(n_2438),
.B(n_190),
.C(n_191),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2447),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2454),
.Y(n_2499)
);

NOR2x1_ASAP7_75t_L g2500 ( 
.A(n_2441),
.B(n_190),
.Y(n_2500)
);

AOI221xp5_ASAP7_75t_L g2501 ( 
.A1(n_2435),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.C(n_194),
.Y(n_2501)
);

NOR3xp33_ASAP7_75t_L g2502 ( 
.A(n_2440),
.B(n_192),
.C(n_193),
.Y(n_2502)
);

OAI21xp5_ASAP7_75t_L g2503 ( 
.A1(n_2455),
.A2(n_2063),
.B(n_2064),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2470),
.B(n_2243),
.Y(n_2504)
);

NAND3xp33_ASAP7_75t_L g2505 ( 
.A(n_2469),
.B(n_194),
.C(n_195),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2468),
.B(n_195),
.Y(n_2506)
);

NOR2x1_ASAP7_75t_L g2507 ( 
.A(n_2444),
.B(n_196),
.Y(n_2507)
);

OAI211xp5_ASAP7_75t_L g2508 ( 
.A1(n_2469),
.A2(n_198),
.B(n_196),
.C(n_197),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2482),
.Y(n_2509)
);

NOR3xp33_ASAP7_75t_L g2510 ( 
.A(n_2487),
.B(n_197),
.C(n_199),
.Y(n_2510)
);

OAI211xp5_ASAP7_75t_L g2511 ( 
.A1(n_2477),
.A2(n_201),
.B(n_199),
.C(n_200),
.Y(n_2511)
);

INVxp67_ASAP7_75t_SL g2512 ( 
.A(n_2483),
.Y(n_2512)
);

NAND4xp25_ASAP7_75t_L g2513 ( 
.A(n_2471),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_2513)
);

NAND4xp25_ASAP7_75t_L g2514 ( 
.A(n_2473),
.B(n_204),
.C(n_202),
.D(n_203),
.Y(n_2514)
);

NAND5xp2_ASAP7_75t_L g2515 ( 
.A(n_2499),
.B(n_207),
.C(n_205),
.D(n_206),
.E(n_208),
.Y(n_2515)
);

NOR2xp33_ASAP7_75t_L g2516 ( 
.A(n_2474),
.B(n_2485),
.Y(n_2516)
);

OAI321xp33_ASAP7_75t_L g2517 ( 
.A1(n_2493),
.A2(n_2268),
.A3(n_2248),
.B1(n_2245),
.B2(n_2243),
.C(n_210),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_L g2518 ( 
.A(n_2501),
.B(n_2475),
.C(n_2478),
.Y(n_2518)
);

NAND4xp25_ASAP7_75t_L g2519 ( 
.A(n_2500),
.B(n_208),
.C(n_205),
.D(n_207),
.Y(n_2519)
);

NAND4xp25_ASAP7_75t_L g2520 ( 
.A(n_2505),
.B(n_211),
.C(n_209),
.D(n_210),
.Y(n_2520)
);

AND4x1_ASAP7_75t_L g2521 ( 
.A(n_2497),
.B(n_213),
.C(n_209),
.D(n_212),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_2507),
.B(n_212),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2484),
.Y(n_2523)
);

AOI211x1_ASAP7_75t_L g2524 ( 
.A1(n_2504),
.A2(n_215),
.B(n_213),
.C(n_214),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2495),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_2502),
.B(n_214),
.Y(n_2526)
);

NOR3xp33_ASAP7_75t_SL g2527 ( 
.A(n_2476),
.B(n_215),
.C(n_216),
.Y(n_2527)
);

OAI22xp5_ASAP7_75t_L g2528 ( 
.A1(n_2491),
.A2(n_2245),
.B1(n_2248),
.B2(n_2243),
.Y(n_2528)
);

NOR4xp25_ASAP7_75t_L g2529 ( 
.A(n_2486),
.B(n_218),
.C(n_216),
.D(n_217),
.Y(n_2529)
);

OR2x2_ASAP7_75t_L g2530 ( 
.A(n_2496),
.B(n_218),
.Y(n_2530)
);

NOR5xp2_ASAP7_75t_L g2531 ( 
.A(n_2489),
.B(n_222),
.C(n_219),
.D(n_220),
.E(n_223),
.Y(n_2531)
);

AOI221xp5_ASAP7_75t_L g2532 ( 
.A1(n_2480),
.A2(n_225),
.B1(n_220),
.B2(n_222),
.C(n_226),
.Y(n_2532)
);

AOI211x1_ASAP7_75t_SL g2533 ( 
.A1(n_2498),
.A2(n_228),
.B(n_225),
.C(n_227),
.Y(n_2533)
);

AOI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_2472),
.A2(n_2506),
.B(n_2508),
.Y(n_2534)
);

OAI211xp5_ASAP7_75t_SL g2535 ( 
.A1(n_2481),
.A2(n_230),
.B(n_227),
.C(n_229),
.Y(n_2535)
);

NOR2xp33_ASAP7_75t_SL g2536 ( 
.A(n_2490),
.B(n_229),
.Y(n_2536)
);

NOR3xp33_ASAP7_75t_SL g2537 ( 
.A(n_2488),
.B(n_2494),
.C(n_2492),
.Y(n_2537)
);

NOR3xp33_ASAP7_75t_L g2538 ( 
.A(n_2503),
.B(n_230),
.C(n_231),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2479),
.Y(n_2539)
);

AND2x2_ASAP7_75t_SL g2540 ( 
.A(n_2497),
.B(n_231),
.Y(n_2540)
);

NAND3xp33_ASAP7_75t_L g2541 ( 
.A(n_2501),
.B(n_232),
.C(n_233),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2493),
.Y(n_2542)
);

NAND4xp75_ASAP7_75t_L g2543 ( 
.A(n_2483),
.B(n_235),
.C(n_233),
.D(n_234),
.Y(n_2543)
);

NAND4xp75_ASAP7_75t_L g2544 ( 
.A(n_2483),
.B(n_238),
.C(n_236),
.D(n_237),
.Y(n_2544)
);

OAI211xp5_ASAP7_75t_L g2545 ( 
.A1(n_2477),
.A2(n_239),
.B(n_236),
.C(n_238),
.Y(n_2545)
);

AOI221xp5_ASAP7_75t_L g2546 ( 
.A1(n_2486),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.C(n_242),
.Y(n_2546)
);

OAI21xp5_ASAP7_75t_SL g2547 ( 
.A1(n_2477),
.A2(n_241),
.B(n_242),
.Y(n_2547)
);

NOR3xp33_ASAP7_75t_L g2548 ( 
.A(n_2487),
.B(n_243),
.C(n_244),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2474),
.B(n_243),
.Y(n_2549)
);

NAND3xp33_ASAP7_75t_L g2550 ( 
.A(n_2501),
.B(n_244),
.C(n_245),
.Y(n_2550)
);

OAI211xp5_ASAP7_75t_SL g2551 ( 
.A1(n_2477),
.A2(n_247),
.B(n_245),
.C(n_246),
.Y(n_2551)
);

NOR2xp67_ASAP7_75t_L g2552 ( 
.A(n_2474),
.B(n_246),
.Y(n_2552)
);

NOR2x1_ASAP7_75t_L g2553 ( 
.A(n_2483),
.B(n_247),
.Y(n_2553)
);

NAND3xp33_ASAP7_75t_SL g2554 ( 
.A(n_2482),
.B(n_248),
.C(n_249),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2483),
.B(n_248),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2483),
.B(n_249),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2482),
.Y(n_2557)
);

NOR4xp25_ASAP7_75t_L g2558 ( 
.A(n_2476),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2558)
);

AOI21xp33_ASAP7_75t_SL g2559 ( 
.A1(n_2482),
.A2(n_250),
.B(n_251),
.Y(n_2559)
);

NAND4xp75_ASAP7_75t_L g2560 ( 
.A(n_2483),
.B(n_254),
.C(n_252),
.D(n_253),
.Y(n_2560)
);

OAI211xp5_ASAP7_75t_SL g2561 ( 
.A1(n_2477),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_2561)
);

AND2x2_ASAP7_75t_L g2562 ( 
.A(n_2500),
.B(n_2287),
.Y(n_2562)
);

INVxp67_ASAP7_75t_SL g2563 ( 
.A(n_2483),
.Y(n_2563)
);

NAND2xp5_ASAP7_75t_L g2564 ( 
.A(n_2483),
.B(n_256),
.Y(n_2564)
);

NAND4xp25_ASAP7_75t_L g2565 ( 
.A(n_2471),
.B(n_259),
.C(n_257),
.D(n_258),
.Y(n_2565)
);

NAND4xp25_ASAP7_75t_L g2566 ( 
.A(n_2471),
.B(n_259),
.C(n_257),
.D(n_258),
.Y(n_2566)
);

AOI221x1_ASAP7_75t_L g2567 ( 
.A1(n_2493),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.C(n_264),
.Y(n_2567)
);

NAND3xp33_ASAP7_75t_L g2568 ( 
.A(n_2501),
.B(n_261),
.C(n_262),
.Y(n_2568)
);

OAI21xp33_ASAP7_75t_SL g2569 ( 
.A1(n_2504),
.A2(n_2287),
.B(n_2283),
.Y(n_2569)
);

OAI22xp33_ASAP7_75t_L g2570 ( 
.A1(n_2473),
.A2(n_2245),
.B1(n_2248),
.B2(n_2243),
.Y(n_2570)
);

OAI322xp33_ASAP7_75t_L g2571 ( 
.A1(n_2536),
.A2(n_263),
.A3(n_264),
.B1(n_265),
.B2(n_266),
.C1(n_267),
.C2(n_268),
.Y(n_2571)
);

XNOR2x1_ASAP7_75t_L g2572 ( 
.A(n_2543),
.B(n_265),
.Y(n_2572)
);

INVxp33_ASAP7_75t_L g2573 ( 
.A(n_2519),
.Y(n_2573)
);

NOR2x1p5_ASAP7_75t_L g2574 ( 
.A(n_2544),
.B(n_267),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2562),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2553),
.Y(n_2576)
);

NOR2xp33_ASAP7_75t_L g2577 ( 
.A(n_2515),
.B(n_269),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_R g2578 ( 
.A(n_2554),
.B(n_269),
.Y(n_2578)
);

HB1xp67_ASAP7_75t_L g2579 ( 
.A(n_2560),
.Y(n_2579)
);

NOR4xp75_ASAP7_75t_L g2580 ( 
.A(n_2542),
.B(n_272),
.C(n_270),
.D(n_271),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2540),
.Y(n_2581)
);

BUFx4f_ASAP7_75t_SL g2582 ( 
.A(n_2542),
.Y(n_2582)
);

AOI331xp33_ASAP7_75t_L g2583 ( 
.A1(n_2516),
.A2(n_272),
.A3(n_273),
.B1(n_275),
.B2(n_277),
.B3(n_278),
.C1(n_279),
.Y(n_2583)
);

NOR2x1_ASAP7_75t_L g2584 ( 
.A(n_2513),
.B(n_273),
.Y(n_2584)
);

NAND3xp33_ASAP7_75t_L g2585 ( 
.A(n_2521),
.B(n_275),
.C(n_277),
.Y(n_2585)
);

INVxp67_ASAP7_75t_L g2586 ( 
.A(n_2549),
.Y(n_2586)
);

AOI32xp33_ASAP7_75t_L g2587 ( 
.A1(n_2551),
.A2(n_2108),
.A3(n_2293),
.B1(n_2290),
.B2(n_281),
.Y(n_2587)
);

OAI21xp5_ASAP7_75t_SL g2588 ( 
.A1(n_2547),
.A2(n_278),
.B(n_279),
.Y(n_2588)
);

BUFx2_ASAP7_75t_SL g2589 ( 
.A(n_2512),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_2559),
.B(n_280),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2527),
.B(n_2290),
.Y(n_2591)
);

OAI211xp5_ASAP7_75t_SL g2592 ( 
.A1(n_2537),
.A2(n_282),
.B(n_280),
.C(n_281),
.Y(n_2592)
);

AOI21xp5_ASAP7_75t_L g2593 ( 
.A1(n_2563),
.A2(n_2555),
.B(n_2522),
.Y(n_2593)
);

AOI221xp5_ASAP7_75t_L g2594 ( 
.A1(n_2558),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.C(n_286),
.Y(n_2594)
);

AOI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2552),
.A2(n_2270),
.B1(n_2248),
.B2(n_2293),
.Y(n_2595)
);

CKINVDCx20_ASAP7_75t_R g2596 ( 
.A(n_2509),
.Y(n_2596)
);

OAI322xp33_ASAP7_75t_L g2597 ( 
.A1(n_2539),
.A2(n_283),
.A3(n_284),
.B1(n_285),
.B2(n_287),
.C1(n_288),
.C2(n_289),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2556),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2529),
.B(n_287),
.Y(n_2599)
);

OAI22xp5_ASAP7_75t_L g2600 ( 
.A1(n_2541),
.A2(n_2286),
.B1(n_2212),
.B2(n_2265),
.Y(n_2600)
);

NOR3xp33_ASAP7_75t_L g2601 ( 
.A(n_2511),
.B(n_2545),
.C(n_2565),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2510),
.B(n_290),
.Y(n_2602)
);

OAI22xp33_ASAP7_75t_L g2603 ( 
.A1(n_2566),
.A2(n_2212),
.B1(n_2266),
.B2(n_2215),
.Y(n_2603)
);

NOR4xp25_ASAP7_75t_L g2604 ( 
.A(n_2561),
.B(n_293),
.C(n_290),
.D(n_292),
.Y(n_2604)
);

AOI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2564),
.A2(n_294),
.B(n_295),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2538),
.A2(n_2270),
.B1(n_2215),
.B2(n_2288),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2530),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2523),
.Y(n_2608)
);

AOI21xp5_ASAP7_75t_L g2609 ( 
.A1(n_2526),
.A2(n_294),
.B(n_295),
.Y(n_2609)
);

OA21x2_ASAP7_75t_L g2610 ( 
.A1(n_2557),
.A2(n_2534),
.B(n_2525),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2524),
.Y(n_2611)
);

OAI21xp33_ASAP7_75t_SL g2612 ( 
.A1(n_2520),
.A2(n_296),
.B(n_297),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2548),
.B(n_296),
.Y(n_2613)
);

HB1xp67_ASAP7_75t_L g2614 ( 
.A(n_2533),
.Y(n_2614)
);

NOR2xp33_ASAP7_75t_R g2615 ( 
.A(n_2514),
.B(n_297),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2550),
.Y(n_2616)
);

OAI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2568),
.A2(n_2289),
.B1(n_2288),
.B2(n_300),
.Y(n_2617)
);

NOR2x1_ASAP7_75t_L g2618 ( 
.A(n_2535),
.B(n_298),
.Y(n_2618)
);

NAND2xp5_ASAP7_75t_L g2619 ( 
.A(n_2546),
.B(n_2532),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2528),
.Y(n_2620)
);

AO22x2_ASAP7_75t_L g2621 ( 
.A1(n_2518),
.A2(n_300),
.B1(n_298),
.B2(n_299),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2531),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2567),
.Y(n_2623)
);

OAI22xp5_ASAP7_75t_L g2624 ( 
.A1(n_2570),
.A2(n_2289),
.B1(n_302),
.B2(n_299),
.Y(n_2624)
);

AOI221xp5_ASAP7_75t_L g2625 ( 
.A1(n_2517),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.C(n_304),
.Y(n_2625)
);

NAND2xp33_ASAP7_75t_R g2626 ( 
.A(n_2569),
.B(n_301),
.Y(n_2626)
);

OAI322xp33_ASAP7_75t_SL g2627 ( 
.A1(n_2539),
.A2(n_304),
.A3(n_305),
.B1(n_306),
.B2(n_307),
.C1(n_309),
.C2(n_310),
.Y(n_2627)
);

AOI221x1_ASAP7_75t_L g2628 ( 
.A1(n_2513),
.A2(n_307),
.B1(n_309),
.B2(n_310),
.C(n_311),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2562),
.Y(n_2629)
);

OAI21xp5_ASAP7_75t_SL g2630 ( 
.A1(n_2547),
.A2(n_311),
.B(n_312),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_2562),
.B(n_314),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2562),
.Y(n_2632)
);

AOI322xp5_ASAP7_75t_L g2633 ( 
.A1(n_2562),
.A2(n_315),
.A3(n_316),
.B1(n_317),
.B2(n_318),
.C1(n_319),
.C2(n_320),
.Y(n_2633)
);

XNOR2xp5_ASAP7_75t_L g2634 ( 
.A(n_2521),
.B(n_315),
.Y(n_2634)
);

AOI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2562),
.A2(n_2270),
.B1(n_2067),
.B2(n_2045),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2591),
.B(n_317),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_2577),
.B(n_318),
.Y(n_2637)
);

NOR4xp75_ASAP7_75t_L g2638 ( 
.A(n_2631),
.B(n_320),
.C(n_321),
.D(n_322),
.Y(n_2638)
);

NAND4xp75_ASAP7_75t_L g2639 ( 
.A(n_2575),
.B(n_321),
.C(n_322),
.D(n_323),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2571),
.B(n_323),
.Y(n_2640)
);

NOR2x1_ASAP7_75t_L g2641 ( 
.A(n_2576),
.B(n_324),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2634),
.Y(n_2642)
);

NAND2x1p5_ASAP7_75t_L g2643 ( 
.A(n_2629),
.B(n_325),
.Y(n_2643)
);

NAND4xp75_ASAP7_75t_L g2644 ( 
.A(n_2632),
.B(n_326),
.C(n_327),
.D(n_328),
.Y(n_2644)
);

NAND4xp75_ASAP7_75t_L g2645 ( 
.A(n_2628),
.B(n_326),
.C(n_327),
.D(n_329),
.Y(n_2645)
);

NAND4xp75_ASAP7_75t_L g2646 ( 
.A(n_2584),
.B(n_329),
.C(n_330),
.D(n_331),
.Y(n_2646)
);

AND2x4_ASAP7_75t_L g2647 ( 
.A(n_2581),
.B(n_330),
.Y(n_2647)
);

AOI22xp5_ASAP7_75t_L g2648 ( 
.A1(n_2582),
.A2(n_331),
.B1(n_332),
.B2(n_333),
.Y(n_2648)
);

OAI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_2595),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_2649)
);

NAND2x1p5_ASAP7_75t_L g2650 ( 
.A(n_2623),
.B(n_334),
.Y(n_2650)
);

INVx3_ASAP7_75t_L g2651 ( 
.A(n_2610),
.Y(n_2651)
);

XNOR2xp5_ASAP7_75t_L g2652 ( 
.A(n_2572),
.B(n_336),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2580),
.B(n_337),
.Y(n_2653)
);

XOR2xp5_ASAP7_75t_L g2654 ( 
.A(n_2596),
.B(n_338),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2610),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2599),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2590),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2621),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2621),
.Y(n_2659)
);

OR2x2_ASAP7_75t_L g2660 ( 
.A(n_2604),
.B(n_339),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2585),
.Y(n_2661)
);

AND2x4_ASAP7_75t_L g2662 ( 
.A(n_2574),
.B(n_339),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2614),
.B(n_340),
.Y(n_2663)
);

NOR2x1p5_ASAP7_75t_L g2664 ( 
.A(n_2602),
.B(n_340),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2622),
.Y(n_2665)
);

NOR2x1_ASAP7_75t_L g2666 ( 
.A(n_2597),
.B(n_341),
.Y(n_2666)
);

NOR2xp33_ASAP7_75t_L g2667 ( 
.A(n_2592),
.B(n_342),
.Y(n_2667)
);

NOR2x1_ASAP7_75t_L g2668 ( 
.A(n_2589),
.B(n_342),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2618),
.Y(n_2669)
);

NOR2xp33_ASAP7_75t_L g2670 ( 
.A(n_2588),
.B(n_343),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2579),
.B(n_343),
.Y(n_2671)
);

NAND4xp75_ASAP7_75t_L g2672 ( 
.A(n_2593),
.B(n_2609),
.C(n_2616),
.D(n_2605),
.Y(n_2672)
);

NAND2x1p5_ASAP7_75t_SL g2673 ( 
.A(n_2620),
.B(n_344),
.Y(n_2673)
);

NOR2x1_ASAP7_75t_L g2674 ( 
.A(n_2630),
.B(n_344),
.Y(n_2674)
);

AND2x4_ASAP7_75t_L g2675 ( 
.A(n_2611),
.B(n_345),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2613),
.Y(n_2676)
);

INVx2_ASAP7_75t_SL g2677 ( 
.A(n_2578),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2613),
.Y(n_2678)
);

NAND4xp75_ASAP7_75t_L g2679 ( 
.A(n_2625),
.B(n_346),
.C(n_347),
.D(n_348),
.Y(n_2679)
);

NOR2xp33_ASAP7_75t_SL g2680 ( 
.A(n_2608),
.B(n_346),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2607),
.Y(n_2681)
);

OR2x2_ASAP7_75t_L g2682 ( 
.A(n_2624),
.B(n_347),
.Y(n_2682)
);

NOR2x1_ASAP7_75t_L g2683 ( 
.A(n_2598),
.B(n_2619),
.Y(n_2683)
);

NAND4xp75_ASAP7_75t_L g2684 ( 
.A(n_2594),
.B(n_348),
.C(n_349),
.D(n_350),
.Y(n_2684)
);

NAND4xp75_ASAP7_75t_L g2685 ( 
.A(n_2612),
.B(n_349),
.C(n_350),
.D(n_351),
.Y(n_2685)
);

AOI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2601),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_L g2687 ( 
.A(n_2633),
.B(n_352),
.Y(n_2687)
);

NAND4xp75_ASAP7_75t_L g2688 ( 
.A(n_2573),
.B(n_353),
.C(n_354),
.D(n_355),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2626),
.Y(n_2689)
);

INVxp33_ASAP7_75t_SL g2690 ( 
.A(n_2615),
.Y(n_2690)
);

NAND3xp33_ASAP7_75t_SL g2691 ( 
.A(n_2650),
.B(n_2586),
.C(n_2587),
.Y(n_2691)
);

NAND5xp2_ASAP7_75t_L g2692 ( 
.A(n_2665),
.B(n_2663),
.C(n_2690),
.D(n_2642),
.E(n_2636),
.Y(n_2692)
);

NAND2x1p5_ASAP7_75t_L g2693 ( 
.A(n_2668),
.B(n_2583),
.Y(n_2693)
);

OR2x2_ASAP7_75t_L g2694 ( 
.A(n_2673),
.B(n_2617),
.Y(n_2694)
);

NOR4xp25_ASAP7_75t_L g2695 ( 
.A(n_2658),
.B(n_2659),
.C(n_2669),
.D(n_2671),
.Y(n_2695)
);

BUFx2_ASAP7_75t_L g2696 ( 
.A(n_2641),
.Y(n_2696)
);

HB1xp67_ASAP7_75t_L g2697 ( 
.A(n_2638),
.Y(n_2697)
);

NAND3xp33_ASAP7_75t_SL g2698 ( 
.A(n_2643),
.B(n_2600),
.C(n_2606),
.Y(n_2698)
);

NAND2xp5_ASAP7_75t_SL g2699 ( 
.A(n_2653),
.B(n_2603),
.Y(n_2699)
);

NOR3xp33_ASAP7_75t_SL g2700 ( 
.A(n_2672),
.B(n_2627),
.C(n_355),
.Y(n_2700)
);

NAND3xp33_ASAP7_75t_SL g2701 ( 
.A(n_2637),
.B(n_2635),
.C(n_356),
.Y(n_2701)
);

NOR4xp25_ASAP7_75t_L g2702 ( 
.A(n_2661),
.B(n_357),
.C(n_358),
.D(n_359),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2675),
.B(n_360),
.Y(n_2703)
);

HB1xp67_ASAP7_75t_L g2704 ( 
.A(n_2645),
.Y(n_2704)
);

NAND3xp33_ASAP7_75t_SL g2705 ( 
.A(n_2687),
.B(n_360),
.C(n_361),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2654),
.Y(n_2706)
);

XNOR2xp5_ASAP7_75t_L g2707 ( 
.A(n_2652),
.B(n_361),
.Y(n_2707)
);

NAND4xp25_ASAP7_75t_L g2708 ( 
.A(n_2667),
.B(n_362),
.C(n_363),
.D(n_365),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_L g2709 ( 
.A(n_2646),
.B(n_362),
.Y(n_2709)
);

NOR5xp2_ASAP7_75t_L g2710 ( 
.A(n_2689),
.B(n_363),
.C(n_365),
.D(n_366),
.E(n_367),
.Y(n_2710)
);

AOI211x1_ASAP7_75t_L g2711 ( 
.A1(n_2649),
.A2(n_368),
.B(n_369),
.C(n_370),
.Y(n_2711)
);

A2O1A1Ixp33_ASAP7_75t_L g2712 ( 
.A1(n_2640),
.A2(n_368),
.B(n_371),
.C(n_372),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2660),
.Y(n_2713)
);

AND3x2_ASAP7_75t_L g2714 ( 
.A(n_2680),
.B(n_371),
.C(n_372),
.Y(n_2714)
);

NOR2x2_ASAP7_75t_L g2715 ( 
.A(n_2685),
.B(n_373),
.Y(n_2715)
);

OR2x6_ASAP7_75t_L g2716 ( 
.A(n_2662),
.B(n_374),
.Y(n_2716)
);

AND5x1_ASAP7_75t_L g2717 ( 
.A(n_2670),
.B(n_374),
.C(n_375),
.D(n_376),
.E(n_377),
.Y(n_2717)
);

NOR3xp33_ASAP7_75t_SL g2718 ( 
.A(n_2652),
.B(n_376),
.C(n_377),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2684),
.Y(n_2719)
);

NOR3xp33_ASAP7_75t_L g2720 ( 
.A(n_2681),
.B(n_2683),
.C(n_2655),
.Y(n_2720)
);

NAND4xp75_ASAP7_75t_L g2721 ( 
.A(n_2666),
.B(n_378),
.C(n_379),
.D(n_380),
.Y(n_2721)
);

NOR3x1_ASAP7_75t_L g2722 ( 
.A(n_2679),
.B(n_381),
.C(n_382),
.Y(n_2722)
);

OA22x2_ASAP7_75t_L g2723 ( 
.A1(n_2686),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_2647),
.B(n_383),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2684),
.B(n_384),
.Y(n_2725)
);

NOR2x1p5_ASAP7_75t_L g2726 ( 
.A(n_2639),
.B(n_385),
.Y(n_2726)
);

NOR3xp33_ASAP7_75t_SL g2727 ( 
.A(n_2676),
.B(n_385),
.C(n_386),
.Y(n_2727)
);

NAND5xp2_ASAP7_75t_L g2728 ( 
.A(n_2656),
.B(n_386),
.C(n_387),
.D(n_388),
.E(n_389),
.Y(n_2728)
);

NOR2x1p5_ASAP7_75t_L g2729 ( 
.A(n_2644),
.B(n_389),
.Y(n_2729)
);

NOR4xp25_ASAP7_75t_L g2730 ( 
.A(n_2651),
.B(n_390),
.C(n_391),
.D(n_392),
.Y(n_2730)
);

NOR3xp33_ASAP7_75t_L g2731 ( 
.A(n_2678),
.B(n_390),
.C(n_392),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2674),
.B(n_393),
.Y(n_2732)
);

OR3x1_ASAP7_75t_L g2733 ( 
.A(n_2657),
.B(n_393),
.C(n_394),
.Y(n_2733)
);

BUFx6f_ASAP7_75t_L g2734 ( 
.A(n_2696),
.Y(n_2734)
);

INVxp67_ASAP7_75t_L g2735 ( 
.A(n_2728),
.Y(n_2735)
);

BUFx6f_ASAP7_75t_L g2736 ( 
.A(n_2713),
.Y(n_2736)
);

BUFx2_ASAP7_75t_L g2737 ( 
.A(n_2716),
.Y(n_2737)
);

HB1xp67_ASAP7_75t_L g2738 ( 
.A(n_2733),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2707),
.Y(n_2739)
);

HB1xp67_ASAP7_75t_L g2740 ( 
.A(n_2716),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2717),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2703),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2714),
.Y(n_2743)
);

BUFx12f_ASAP7_75t_L g2744 ( 
.A(n_2694),
.Y(n_2744)
);

HB1xp67_ASAP7_75t_L g2745 ( 
.A(n_2726),
.Y(n_2745)
);

HB1xp67_ASAP7_75t_L g2746 ( 
.A(n_2729),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2715),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2724),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2704),
.Y(n_2749)
);

AOI21xp33_ASAP7_75t_L g2750 ( 
.A1(n_2709),
.A2(n_2677),
.B(n_2682),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2725),
.Y(n_2751)
);

NOR2xp33_ASAP7_75t_L g2752 ( 
.A(n_2708),
.B(n_2688),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2727),
.B(n_2664),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2730),
.B(n_2648),
.Y(n_2754)
);

XOR2xp5_ASAP7_75t_L g2755 ( 
.A(n_2721),
.B(n_394),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2723),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2732),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_2718),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2706),
.Y(n_2759)
);

INVxp33_ASAP7_75t_L g2760 ( 
.A(n_2697),
.Y(n_2760)
);

CKINVDCx6p67_ASAP7_75t_R g2761 ( 
.A(n_2719),
.Y(n_2761)
);

BUFx10_ASAP7_75t_L g2762 ( 
.A(n_2695),
.Y(n_2762)
);

AOI32xp33_ASAP7_75t_L g2763 ( 
.A1(n_2760),
.A2(n_2720),
.A3(n_2699),
.B1(n_2731),
.B2(n_2722),
.Y(n_2763)
);

OAI322xp33_ASAP7_75t_L g2764 ( 
.A1(n_2755),
.A2(n_2693),
.A3(n_2692),
.B1(n_2700),
.B2(n_2705),
.C1(n_2691),
.C2(n_2698),
.Y(n_2764)
);

AOI322xp5_ASAP7_75t_L g2765 ( 
.A1(n_2752),
.A2(n_2701),
.A3(n_2712),
.B1(n_2711),
.B2(n_2710),
.C1(n_2702),
.C2(n_401),
.Y(n_2765)
);

NOR2x1_ASAP7_75t_L g2766 ( 
.A(n_2737),
.B(n_395),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2762),
.Y(n_2767)
);

AOI32xp33_ASAP7_75t_L g2768 ( 
.A1(n_2756),
.A2(n_396),
.A3(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_2768)
);

OAI322xp33_ASAP7_75t_L g2769 ( 
.A1(n_2735),
.A2(n_396),
.A3(n_398),
.B1(n_399),
.B2(n_400),
.C1(n_402),
.C2(n_403),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2741),
.Y(n_2770)
);

AOI22xp5_ASAP7_75t_L g2771 ( 
.A1(n_2749),
.A2(n_403),
.B1(n_404),
.B2(n_405),
.Y(n_2771)
);

OAI211xp5_ASAP7_75t_L g2772 ( 
.A1(n_2750),
.A2(n_404),
.B(n_406),
.C(n_407),
.Y(n_2772)
);

OAI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2761),
.A2(n_406),
.B1(n_408),
.B2(n_409),
.Y(n_2773)
);

AOI322xp5_ASAP7_75t_L g2774 ( 
.A1(n_2738),
.A2(n_408),
.A3(n_409),
.B1(n_410),
.B2(n_411),
.C1(n_412),
.C2(n_413),
.Y(n_2774)
);

AOI22xp5_ASAP7_75t_L g2775 ( 
.A1(n_2744),
.A2(n_410),
.B1(n_411),
.B2(n_412),
.Y(n_2775)
);

OAI322xp33_ASAP7_75t_L g2776 ( 
.A1(n_2743),
.A2(n_414),
.A3(n_415),
.B1(n_416),
.B2(n_417),
.C1(n_418),
.C2(n_419),
.Y(n_2776)
);

AOI222xp33_ASAP7_75t_L g2777 ( 
.A1(n_2758),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.C1(n_418),
.C2(n_419),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2734),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.Y(n_2778)
);

OAI211xp5_ASAP7_75t_SL g2779 ( 
.A1(n_2751),
.A2(n_420),
.B(n_422),
.C(n_423),
.Y(n_2779)
);

AOI322xp5_ASAP7_75t_L g2780 ( 
.A1(n_2740),
.A2(n_2746),
.A3(n_2745),
.B1(n_2747),
.B2(n_2757),
.C1(n_2753),
.C2(n_2739),
.Y(n_2780)
);

OAI221xp5_ASAP7_75t_L g2781 ( 
.A1(n_2754),
.A2(n_423),
.B1(n_424),
.B2(n_425),
.C(n_427),
.Y(n_2781)
);

OAI211xp5_ASAP7_75t_L g2782 ( 
.A1(n_2759),
.A2(n_425),
.B(n_429),
.C(n_430),
.Y(n_2782)
);

OA22x2_ASAP7_75t_L g2783 ( 
.A1(n_2767),
.A2(n_2742),
.B1(n_2748),
.B2(n_2734),
.Y(n_2783)
);

AOI22xp5_ASAP7_75t_L g2784 ( 
.A1(n_2770),
.A2(n_2736),
.B1(n_2766),
.B2(n_2779),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2764),
.Y(n_2785)
);

AOI22x1_ASAP7_75t_SL g2786 ( 
.A1(n_2777),
.A2(n_2736),
.B1(n_431),
.B2(n_433),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2772),
.Y(n_2787)
);

CKINVDCx20_ASAP7_75t_R g2788 ( 
.A(n_2775),
.Y(n_2788)
);

AO22x2_ASAP7_75t_L g2789 ( 
.A1(n_2782),
.A2(n_430),
.B1(n_431),
.B2(n_433),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2773),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2776),
.Y(n_2791)
);

O2A1O1Ixp33_ASAP7_75t_L g2792 ( 
.A1(n_2781),
.A2(n_435),
.B(n_436),
.C(n_437),
.Y(n_2792)
);

AO22x2_ASAP7_75t_L g2793 ( 
.A1(n_2763),
.A2(n_435),
.B1(n_436),
.B2(n_437),
.Y(n_2793)
);

AOI22xp5_ASAP7_75t_L g2794 ( 
.A1(n_2771),
.A2(n_438),
.B1(n_439),
.B2(n_440),
.Y(n_2794)
);

XNOR2xp5_ASAP7_75t_L g2795 ( 
.A(n_2786),
.B(n_2778),
.Y(n_2795)
);

NAND3xp33_ASAP7_75t_L g2796 ( 
.A(n_2784),
.B(n_2780),
.C(n_2765),
.Y(n_2796)
);

NOR2x1p5_ASAP7_75t_L g2797 ( 
.A(n_2791),
.B(n_2768),
.Y(n_2797)
);

NOR3x2_ASAP7_75t_L g2798 ( 
.A(n_2783),
.B(n_2769),
.C(n_2774),
.Y(n_2798)
);

OAI222xp33_ASAP7_75t_L g2799 ( 
.A1(n_2785),
.A2(n_438),
.B1(n_439),
.B2(n_441),
.C1(n_442),
.C2(n_443),
.Y(n_2799)
);

AOI21xp5_ASAP7_75t_L g2800 ( 
.A1(n_2787),
.A2(n_2790),
.B(n_2792),
.Y(n_2800)
);

NAND3xp33_ASAP7_75t_L g2801 ( 
.A(n_2794),
.B(n_441),
.C(n_442),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2789),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_2802),
.B(n_2793),
.Y(n_2803)
);

AOI21xp5_ASAP7_75t_L g2804 ( 
.A1(n_2800),
.A2(n_2788),
.B(n_445),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_SL g2805 ( 
.A1(n_2795),
.A2(n_443),
.B1(n_445),
.B2(n_447),
.Y(n_2805)
);

AOI21xp5_ASAP7_75t_L g2806 ( 
.A1(n_2796),
.A2(n_2801),
.B(n_2799),
.Y(n_2806)
);

XNOR2xp5_ASAP7_75t_L g2807 ( 
.A(n_2798),
.B(n_447),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2797),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2807),
.Y(n_2809)
);

AOI21xp33_ASAP7_75t_SL g2810 ( 
.A1(n_2808),
.A2(n_448),
.B(n_449),
.Y(n_2810)
);

OAI22x1_ASAP7_75t_SL g2811 ( 
.A1(n_2806),
.A2(n_448),
.B1(n_450),
.B2(n_451),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2804),
.B(n_451),
.Y(n_2812)
);

OAI22x1_ASAP7_75t_SL g2813 ( 
.A1(n_2803),
.A2(n_452),
.B1(n_453),
.B2(n_454),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2812),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2809),
.B(n_2805),
.Y(n_2815)
);

AOI221xp5_ASAP7_75t_L g2816 ( 
.A1(n_2814),
.A2(n_2810),
.B1(n_2811),
.B2(n_2813),
.C(n_458),
.Y(n_2816)
);

AOI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2816),
.A2(n_2815),
.B1(n_456),
.B2(n_457),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2816),
.A2(n_454),
.B1(n_458),
.B2(n_459),
.Y(n_2818)
);

NAND3xp33_ASAP7_75t_L g2819 ( 
.A(n_2817),
.B(n_459),
.C(n_460),
.Y(n_2819)
);

AOI21xp5_ASAP7_75t_L g2820 ( 
.A1(n_2819),
.A2(n_2818),
.B(n_462),
.Y(n_2820)
);

AOI221x1_ASAP7_75t_L g2821 ( 
.A1(n_2820),
.A2(n_461),
.B1(n_462),
.B2(n_463),
.C(n_464),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2821),
.A2(n_461),
.B(n_463),
.Y(n_2822)
);

AOI211xp5_ASAP7_75t_L g2823 ( 
.A1(n_2822),
.A2(n_464),
.B(n_465),
.C(n_466),
.Y(n_2823)
);


endmodule