module real_aes_180_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_756;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g550 ( .A(n_0), .B(n_176), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_1), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_2), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g134 ( .A(n_3), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_4), .B(n_512), .Y(n_511) );
NAND2xp33_ASAP7_75t_SL g593 ( .A(n_5), .B(n_163), .Y(n_593) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_6), .B(n_143), .Y(n_167) );
INVx1_ASAP7_75t_L g586 ( .A(n_7), .Y(n_586) );
INVx1_ASAP7_75t_L g189 ( .A(n_8), .Y(n_189) );
CKINVDCx16_ASAP7_75t_R g819 ( .A(n_9), .Y(n_819) );
CKINVDCx5p33_ASAP7_75t_R g205 ( .A(n_10), .Y(n_205) );
AND2x2_ASAP7_75t_L g509 ( .A(n_11), .B(n_220), .Y(n_509) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_13), .Y(n_109) );
INVx1_ASAP7_75t_L g177 ( .A(n_14), .Y(n_177) );
AOI221x1_ASAP7_75t_L g589 ( .A1(n_15), .A2(n_194), .B1(n_514), .B2(n_590), .C(n_592), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_16), .B(n_512), .Y(n_573) );
INVx1_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
INVx1_ASAP7_75t_L g174 ( .A(n_18), .Y(n_174) );
INVx1_ASAP7_75t_SL g249 ( .A(n_19), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_20), .B(n_154), .Y(n_153) );
AOI33xp33_ASAP7_75t_L g226 ( .A1(n_21), .A2(n_50), .A3(n_131), .B1(n_149), .B2(n_227), .B3(n_228), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_22), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_23), .B(n_176), .Y(n_516) );
AOI221xp5_ASAP7_75t_SL g560 ( .A1(n_24), .A2(n_39), .B1(n_512), .B2(n_514), .C(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g198 ( .A(n_25), .Y(n_198) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_26), .A2(n_89), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g144 ( .A(n_26), .B(n_89), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_27), .B(n_179), .Y(n_577) );
INVxp67_ASAP7_75t_L g588 ( .A(n_28), .Y(n_588) );
AND2x2_ASAP7_75t_L g535 ( .A(n_29), .B(n_219), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_30), .B(n_187), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_31), .A2(n_514), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_32), .B(n_179), .Y(n_562) );
AND2x2_ASAP7_75t_L g137 ( .A(n_33), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g148 ( .A(n_33), .Y(n_148) );
AND2x2_ASAP7_75t_L g163 ( .A(n_33), .B(n_134), .Y(n_163) );
OR2x6_ASAP7_75t_L g111 ( .A(n_34), .B(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_35), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_36), .B(n_187), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_37), .A2(n_128), .B1(n_140), .B2(n_143), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_38), .B(n_160), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_40), .A2(n_80), .B1(n_146), .B2(n_514), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_41), .B(n_154), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_42), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_43), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_44), .B(n_176), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_45), .B(n_165), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_46), .B(n_154), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_47), .Y(n_139) );
AND2x2_ASAP7_75t_L g553 ( .A(n_48), .B(n_219), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_49), .B(n_219), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_51), .B(n_154), .Y(n_217) );
INVx1_ASAP7_75t_L g132 ( .A(n_52), .Y(n_132) );
INVx1_ASAP7_75t_L g156 ( .A(n_52), .Y(n_156) );
AND2x2_ASAP7_75t_L g218 ( .A(n_53), .B(n_219), .Y(n_218) );
AOI221xp5_ASAP7_75t_L g186 ( .A1(n_54), .A2(n_73), .B1(n_146), .B2(n_187), .C(n_188), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_55), .B(n_187), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_56), .B(n_512), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_57), .B(n_140), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g237 ( .A1(n_58), .A2(n_146), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g526 ( .A(n_59), .B(n_219), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_60), .B(n_179), .Y(n_551) );
INVx1_ASAP7_75t_L g170 ( .A(n_61), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_62), .B(n_176), .Y(n_524) );
AND2x2_ASAP7_75t_SL g578 ( .A(n_63), .B(n_220), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_64), .A2(n_514), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g216 ( .A(n_65), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_66), .B(n_179), .Y(n_517) );
AND2x2_ASAP7_75t_SL g542 ( .A(n_67), .B(n_165), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_68), .A2(n_146), .B(n_215), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_69), .A2(n_87), .B1(n_494), .B2(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_69), .Y(n_801) );
INVx1_ASAP7_75t_L g138 ( .A(n_70), .Y(n_138) );
INVx1_ASAP7_75t_L g158 ( .A(n_70), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_71), .B(n_187), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_72), .Y(n_115) );
AND2x2_ASAP7_75t_L g251 ( .A(n_74), .B(n_194), .Y(n_251) );
INVx1_ASAP7_75t_L g171 ( .A(n_75), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_76), .A2(n_146), .B(n_248), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g145 ( .A1(n_77), .A2(n_146), .B(n_152), .C(n_164), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_78), .B(n_512), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_79), .A2(n_83), .B1(n_187), .B2(n_512), .Y(n_540) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
AND2x2_ASAP7_75t_SL g235 ( .A(n_82), .B(n_194), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_84), .A2(n_146), .B1(n_224), .B2(n_225), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_85), .B(n_176), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_86), .B(n_176), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g120 ( .A(n_87), .B(n_121), .C(n_348), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_87), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_88), .A2(n_514), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g239 ( .A(n_90), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_91), .B(n_179), .Y(n_523) );
AND2x2_ASAP7_75t_L g230 ( .A(n_92), .B(n_194), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g195 ( .A1(n_93), .A2(n_196), .B(n_197), .C(n_199), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_94), .B(n_512), .Y(n_552) );
INVxp67_ASAP7_75t_L g591 ( .A(n_95), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_96), .B(n_179), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_97), .A2(n_514), .B(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g106 ( .A(n_98), .Y(n_106) );
BUFx2_ASAP7_75t_SL g796 ( .A(n_98), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_99), .B(n_154), .Y(n_240) );
AOI21xp33_ASAP7_75t_SL g100 ( .A1(n_101), .A2(n_813), .B(n_820), .Y(n_100) );
OA21x2_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_116), .B(n_794), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g102 ( .A(n_103), .B(n_107), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_107), .A2(n_799), .B(n_802), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_107), .B(n_811), .Y(n_810) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_115), .Y(n_107) );
BUFx2_ASAP7_75t_R g812 ( .A(n_108), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x6_ASAP7_75t_SL g501 ( .A(n_109), .B(n_111), .Y(n_501) );
OR2x6_ASAP7_75t_SL g785 ( .A(n_109), .B(n_110), .Y(n_785) );
OR2x2_ASAP7_75t_L g793 ( .A(n_109), .B(n_111), .Y(n_793) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OAI21xp5_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_786), .B(n_787), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_498), .B1(n_502), .B2(n_783), .Y(n_118) );
AO22x2_ASAP7_75t_L g788 ( .A1(n_119), .A2(n_499), .B1(n_502), .B2(n_784), .Y(n_788) );
AOI211x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_390), .B(n_491), .C(n_495), .Y(n_119) );
INVxp67_ASAP7_75t_L g493 ( .A(n_121), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_121), .B(n_435), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_295), .C(n_328), .Y(n_121) );
AOI211xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_252), .B(n_261), .C(n_285), .Y(n_122) );
OAI21xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_181), .B(n_231), .Y(n_123) );
OR2x2_ASAP7_75t_L g305 ( .A(n_124), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g433 ( .A(n_124), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g417 ( .A(n_125), .B(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_125), .A2(n_438), .B1(n_441), .B2(n_442), .Y(n_437) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_166), .Y(n_125) );
INVx1_ASAP7_75t_L g284 ( .A(n_126), .Y(n_284) );
AND2x4_ASAP7_75t_L g301 ( .A(n_126), .B(n_282), .Y(n_301) );
INVx2_ASAP7_75t_L g323 ( .A(n_126), .Y(n_323) );
AND2x2_ASAP7_75t_L g371 ( .A(n_126), .B(n_234), .Y(n_371) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_126), .Y(n_385) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_145), .Y(n_126) );
NOR3xp33_ASAP7_75t_L g128 ( .A(n_129), .B(n_135), .C(n_139), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g187 ( .A(n_130), .B(n_136), .Y(n_187) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
OR2x6_ASAP7_75t_L g161 ( .A(n_131), .B(n_150), .Y(n_161) );
INVxp33_ASAP7_75t_L g227 ( .A(n_131), .Y(n_227) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g151 ( .A(n_132), .B(n_134), .Y(n_151) );
AND2x4_ASAP7_75t_L g179 ( .A(n_132), .B(n_157), .Y(n_179) );
HB1xp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x6_ASAP7_75t_L g514 ( .A(n_137), .B(n_151), .Y(n_514) );
INVx2_ASAP7_75t_L g150 ( .A(n_138), .Y(n_150) );
AND2x6_ASAP7_75t_L g176 ( .A(n_138), .B(n_155), .Y(n_176) );
INVx4_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_140), .B(n_204), .Y(n_203) );
AOI21x1_ASAP7_75t_L g546 ( .A1(n_140), .A2(n_547), .B(n_553), .Y(n_546) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx4f_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
AND2x4_ASAP7_75t_L g143 ( .A(n_142), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_SL g220 ( .A(n_142), .B(n_144), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_143), .B(n_162), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_143), .A2(n_237), .B(n_241), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_143), .A2(n_511), .B(n_513), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_143), .B(n_586), .Y(n_585) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_143), .B(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_143), .B(n_591), .Y(n_590) );
NOR3xp33_ASAP7_75t_L g592 ( .A(n_143), .B(n_172), .C(n_593), .Y(n_592) );
INVxp67_ASAP7_75t_L g206 ( .A(n_146), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_146), .A2(n_187), .B1(n_585), .B2(n_587), .Y(n_584) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NOR2x1p5_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
INVx1_ASAP7_75t_L g228 ( .A(n_149), .Y(n_228) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_159), .B(n_162), .Y(n_152) );
INVx1_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
AND2x4_ASAP7_75t_L g512 ( .A(n_154), .B(n_163), .Y(n_512) );
AND2x4_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI22xp5_ASAP7_75t_L g169 ( .A1(n_161), .A2(n_170), .B1(n_171), .B2(n_172), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_SL g188 ( .A1(n_161), .A2(n_162), .B(n_189), .C(n_190), .Y(n_188) );
INVxp67_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g215 ( .A1(n_161), .A2(n_162), .B(n_216), .C(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_161), .A2(n_162), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g248 ( .A1(n_161), .A2(n_162), .B(n_249), .C(n_250), .Y(n_248) );
INVx1_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_162), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_162), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_162), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_162), .A2(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_162), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_162), .A2(n_576), .B(n_577), .Y(n_575) );
INVx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_163), .Y(n_199) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_222), .B(n_230), .Y(n_221) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_164), .A2(n_222), .B(n_230), .Y(n_266) );
AOI21x1_ASAP7_75t_L g538 ( .A1(n_164), .A2(n_539), .B(n_542), .Y(n_538) );
INVx2_ASAP7_75t_SL g164 ( .A(n_165), .Y(n_164) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_165), .A2(n_186), .B(n_191), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_165), .A2(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g242 ( .A(n_166), .B(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g271 ( .A(n_166), .Y(n_271) );
INVx3_ASAP7_75t_L g282 ( .A(n_166), .Y(n_282) );
AND2x4_ASAP7_75t_L g166 ( .A(n_167), .B(n_168), .Y(n_166) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_173), .B(n_180), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_172), .B(n_198), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B1(n_177), .B2(n_178), .Y(n_173) );
INVxp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVxp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_181), .A2(n_366), .B1(n_368), .B2(n_370), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_181), .B(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_183), .B(n_209), .Y(n_182) );
INVx3_ASAP7_75t_L g255 ( .A(n_183), .Y(n_255) );
AND2x2_ASAP7_75t_L g263 ( .A(n_183), .B(n_264), .Y(n_263) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_183), .Y(n_293) );
NAND2x1_ASAP7_75t_SL g382 ( .A(n_183), .B(n_254), .Y(n_382) );
AND2x4_ASAP7_75t_L g183 ( .A(n_184), .B(n_192), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g260 ( .A(n_185), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_185), .B(n_266), .Y(n_278) );
AND2x2_ASAP7_75t_L g291 ( .A(n_185), .B(n_192), .Y(n_291) );
AND2x4_ASAP7_75t_L g298 ( .A(n_185), .B(n_299), .Y(n_298) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_185), .Y(n_347) );
INVx1_ASAP7_75t_L g357 ( .A(n_185), .Y(n_357) );
INVxp67_ASAP7_75t_L g440 ( .A(n_185), .Y(n_440) );
INVx1_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
INVx1_ASAP7_75t_L g258 ( .A(n_192), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_192), .B(n_268), .Y(n_277) );
INVx2_ASAP7_75t_L g345 ( .A(n_192), .Y(n_345) );
INVx1_ASAP7_75t_L g388 ( .A(n_192), .Y(n_388) );
OR2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B1(n_200), .B2(n_201), .Y(n_193) );
INVx3_ASAP7_75t_L g201 ( .A(n_194), .Y(n_201) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_201), .A2(n_212), .B(n_218), .Y(n_211) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_201), .A2(n_212), .B(n_218), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_206), .B1(n_207), .B2(n_208), .Y(n_202) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g314 ( .A(n_209), .B(n_291), .Y(n_314) );
AND2x2_ASAP7_75t_L g463 ( .A(n_209), .B(n_387), .Y(n_463) );
AND2x2_ASAP7_75t_L g469 ( .A(n_209), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_209), .B(n_430), .Y(n_480) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NOR2x1_ASAP7_75t_L g259 ( .A(n_211), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g406 ( .A(n_211), .B(n_345), .Y(n_406) );
AND2x2_ASAP7_75t_L g410 ( .A(n_211), .B(n_265), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g244 ( .A(n_219), .Y(n_244) );
OA21x2_ASAP7_75t_L g559 ( .A1(n_219), .A2(n_560), .B(n_564), .Y(n_559) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g254 ( .A(n_221), .Y(n_254) );
INVx2_ASAP7_75t_L g299 ( .A(n_221), .Y(n_299) );
AND2x2_ASAP7_75t_L g344 ( .A(n_221), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_223), .B(n_229), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_242), .Y(n_232) );
OR2x6_ASAP7_75t_L g412 ( .A(n_233), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g416 ( .A(n_233), .B(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx4_ASAP7_75t_L g275 ( .A(n_234), .Y(n_275) );
AND2x4_ASAP7_75t_L g283 ( .A(n_234), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g318 ( .A(n_234), .B(n_243), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_234), .B(n_341), .Y(n_364) );
AND2x2_ASAP7_75t_L g380 ( .A(n_234), .B(n_271), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_234), .B(n_336), .Y(n_434) );
INVx2_ASAP7_75t_L g449 ( .A(n_234), .Y(n_449) );
OR2x6_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g294 ( .A(n_242), .B(n_283), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_242), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_SL g398 ( .A(n_242), .B(n_321), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_242), .B(n_334), .Y(n_427) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_243), .Y(n_273) );
AND2x2_ASAP7_75t_L g281 ( .A(n_243), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_243), .Y(n_304) );
INVx2_ASAP7_75t_L g307 ( .A(n_243), .Y(n_307) );
INVx1_ASAP7_75t_L g340 ( .A(n_243), .Y(n_340) );
INVx1_ASAP7_75t_L g418 ( .A(n_243), .Y(n_418) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_245), .B(n_251), .Y(n_243) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_244), .A2(n_520), .B(n_526), .Y(n_519) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_244), .A2(n_529), .B(n_535), .Y(n_528) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_244), .A2(n_529), .B(n_535), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_253), .B(n_256), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_254), .B(n_257), .Y(n_330) );
AND4x1_ASAP7_75t_SL g420 ( .A(n_254), .B(n_395), .C(n_421), .D(n_423), .Y(n_420) );
OR2x2_ASAP7_75t_L g474 ( .A(n_254), .B(n_475), .Y(n_474) );
OR2x2_ASAP7_75t_L g366 ( .A(n_255), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
AND2x2_ASAP7_75t_L g309 ( .A(n_258), .B(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_258), .B(n_267), .Y(n_432) );
AND2x2_ASAP7_75t_L g378 ( .A(n_259), .B(n_344), .Y(n_378) );
OAI32xp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_269), .A3(n_274), .B1(n_276), .B2(n_279), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g429 ( .A(n_264), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g442 ( .A(n_264), .B(n_360), .Y(n_442) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g405 ( .A(n_265), .Y(n_405) );
AND2x2_ASAP7_75t_L g439 ( .A(n_265), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_266), .B(n_268), .Y(n_367) );
INVx3_ASAP7_75t_L g290 ( .A(n_267), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_267), .B(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_268), .Y(n_327) );
AND2x2_ASAP7_75t_L g346 ( .A(n_268), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g374 ( .A(n_270), .Y(n_374) );
NAND2x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g320 ( .A(n_271), .Y(n_320) );
NOR2x1_ASAP7_75t_L g487 ( .A(n_271), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_274), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g312 ( .A(n_275), .B(n_280), .Y(n_312) );
AND2x4_ASAP7_75t_L g334 ( .A(n_275), .B(n_284), .Y(n_334) );
AND2x4_ASAP7_75t_SL g384 ( .A(n_275), .B(n_385), .Y(n_384) );
NOR2x1_ASAP7_75t_L g396 ( .A(n_275), .B(n_352), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_276), .A2(n_472), .B1(n_474), .B2(n_476), .Y(n_471) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx2_ASAP7_75t_SL g484 ( .A(n_277), .Y(n_484) );
INVx2_ASAP7_75t_L g310 ( .A(n_278), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_281), .B(n_287), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_281), .A2(n_483), .B1(n_486), .B2(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g341 ( .A(n_282), .Y(n_341) );
AND2x2_ASAP7_75t_L g414 ( .A(n_282), .B(n_323), .Y(n_414) );
INVx2_ASAP7_75t_L g287 ( .A(n_283), .Y(n_287) );
OAI21xp5_ASAP7_75t_SL g285 ( .A1(n_286), .A2(n_288), .B(n_292), .Y(n_285) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_289), .A2(n_444), .B1(n_447), .B2(n_448), .Y(n_443) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_290), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_290), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g459 ( .A(n_290), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NOR3xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_311), .C(n_315), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B1(n_305), .B2(n_308), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g325 ( .A(n_298), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g386 ( .A(n_298), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g399 ( .A(n_298), .B(n_388), .Y(n_399) );
AND2x2_ASAP7_75t_L g447 ( .A(n_298), .B(n_406), .Y(n_447) );
AND2x2_ASAP7_75t_L g483 ( .A(n_298), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx4_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
AND2x2_ASAP7_75t_L g448 ( .A(n_301), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g453 ( .A(n_304), .Y(n_453) );
AND2x2_ASAP7_75t_L g461 ( .A(n_304), .B(n_414), .Y(n_461) );
INVx1_ASAP7_75t_L g363 ( .A(n_306), .Y(n_363) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_309), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_310), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B(n_324), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_317), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
AOI21xp33_ASAP7_75t_SL g328 ( .A1(n_320), .A2(n_329), .B(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_L g369 ( .A(n_320), .B(n_334), .Y(n_369) );
AND2x4_ASAP7_75t_L g338 ( .A(n_321), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_SL g426 ( .A(n_321), .B(n_418), .Y(n_426) );
INVx2_ASAP7_75t_SL g454 ( .A(n_321), .Y(n_454) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AOI21xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_337), .B(n_342), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_334), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_334), .B(n_339), .Y(n_482) );
AND2x2_ASAP7_75t_L g379 ( .A(n_335), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g383 ( .A(n_335), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g422 ( .A(n_335), .Y(n_422) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_335), .B(n_352), .Y(n_441) );
INVx1_ASAP7_75t_L g470 ( .A(n_335), .Y(n_470) );
INVx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_SL g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_340), .B(n_414), .Y(n_446) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g354 ( .A(n_344), .Y(n_354) );
AND2x2_ASAP7_75t_L g360 ( .A(n_345), .B(n_357), .Y(n_360) );
INVxp67_ASAP7_75t_L g496 ( .A(n_348), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_348), .B(n_391), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_375), .Y(n_348) );
NOR3xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_365), .C(n_372), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B1(n_358), .B2(n_361), .Y(n_350) );
INVx2_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
NAND2xp5_ASAP7_75t_R g407 ( .A(n_352), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx3_ASAP7_75t_L g403 ( .A(n_356), .Y(n_403) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g455 ( .A(n_359), .Y(n_455) );
INVx2_ASAP7_75t_L g475 ( .A(n_360), .Y(n_475) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_362), .A2(n_479), .B1(n_481), .B2(n_483), .Y(n_478) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g372 ( .A(n_366), .B(n_371), .C(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI222xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_381), .B2(n_383), .C1(n_386), .C2(n_389), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_380), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g408 ( .A(n_384), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_384), .B(n_453), .Y(n_476) );
INVx1_ASAP7_75t_L g430 ( .A(n_387), .Y(n_430) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_387), .A2(n_466), .B(n_467), .Y(n_465) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g409 ( .A(n_388), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_435), .Y(n_390) );
INVxp67_ASAP7_75t_L g497 ( .A(n_391), .Y(n_497) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_400), .C(n_419), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_401), .A2(n_407), .B1(n_409), .B2(n_411), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx2_ASAP7_75t_L g468 ( .A(n_403), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g404 ( .A(n_405), .B(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g438 ( .A(n_406), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_415), .A2(n_457), .B1(n_460), .B2(n_462), .Y(n_456) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g486 ( .A(n_418), .B(n_487), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_424), .C(n_431), .Y(n_419) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x2_ASAP7_75t_L g473 ( .A(n_422), .B(n_448), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_427), .B(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVxp67_ASAP7_75t_L g492 ( .A(n_435), .Y(n_492) );
NAND4xp75_ASAP7_75t_L g435 ( .A(n_436), .B(n_450), .C(n_464), .D(n_477), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_443), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g490 ( .A(n_439), .B(n_484), .Y(n_490) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g488 ( .A(n_449), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_455), .B(n_456), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_454), .B(n_468), .Y(n_467) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_469), .B(n_471), .Y(n_464) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_485), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
AOI21xp5_ASAP7_75t_SL g495 ( .A1(n_494), .A2(n_496), .B(n_497), .Y(n_495) );
INVx4_ASAP7_75t_SL g498 ( .A(n_499), .Y(n_498) );
INVx3_ASAP7_75t_SL g499 ( .A(n_500), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_501), .Y(n_500) );
INVx3_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_713), .Y(n_503) );
NOR4xp25_ASAP7_75t_SL g504 ( .A(n_505), .B(n_606), .C(n_650), .D(n_677), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_569), .B1(n_579), .B2(n_594), .C(n_596), .Y(n_505) );
AOI32xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_536), .A3(n_543), .B1(n_554), .B2(n_565), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_507), .B(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_507), .A2(n_719), .B1(n_777), .B2(n_780), .Y(n_776) );
AND2x4_ASAP7_75t_SL g507 ( .A(n_508), .B(n_518), .Y(n_507) );
INVx5_ASAP7_75t_L g568 ( .A(n_508), .Y(n_568) );
OR2x2_ASAP7_75t_L g595 ( .A(n_508), .B(n_567), .Y(n_595) );
AND2x4_ASAP7_75t_L g597 ( .A(n_508), .B(n_528), .Y(n_597) );
INVx2_ASAP7_75t_L g612 ( .A(n_508), .Y(n_612) );
OR2x2_ASAP7_75t_L g624 ( .A(n_508), .B(n_537), .Y(n_624) );
AND2x2_ASAP7_75t_L g631 ( .A(n_508), .B(n_527), .Y(n_631) );
AND2x2_ASAP7_75t_SL g673 ( .A(n_508), .B(n_556), .Y(n_673) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_508), .Y(n_730) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
INVx3_ASAP7_75t_SL g625 ( .A(n_518), .Y(n_625) );
AND2x2_ASAP7_75t_L g644 ( .A(n_518), .B(n_568), .Y(n_644) );
AOI32xp33_ASAP7_75t_L g759 ( .A1(n_518), .A2(n_630), .A3(n_660), .B1(n_690), .B2(n_725), .Y(n_759) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
AND2x2_ASAP7_75t_L g599 ( .A(n_519), .B(n_537), .Y(n_599) );
OR2x2_ASAP7_75t_L g615 ( .A(n_519), .B(n_528), .Y(n_615) );
INVx1_ASAP7_75t_L g638 ( .A(n_519), .Y(n_638) );
INVx2_ASAP7_75t_L g654 ( .A(n_519), .Y(n_654) );
AND2x2_ASAP7_75t_L g691 ( .A(n_519), .B(n_556), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_519), .B(n_528), .Y(n_710) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_519), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g746 ( .A(n_528), .B(n_537), .Y(n_746) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_528), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_534), .Y(n_529) );
OR2x2_ASAP7_75t_L g594 ( .A(n_536), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g600 ( .A(n_536), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g613 ( .A(n_536), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g775 ( .A(n_536), .B(n_644), .Y(n_775) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g704 ( .A(n_537), .B(n_654), .Y(n_704) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_538), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_543), .B(n_671), .Y(n_773) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_544), .B(n_721), .Y(n_720) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g558 ( .A(n_545), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g580 ( .A(n_545), .Y(n_580) );
AND2x2_ASAP7_75t_L g604 ( .A(n_545), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_545), .B(n_582), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_545), .B(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g662 ( .A(n_545), .Y(n_662) );
OR2x2_ASAP7_75t_L g681 ( .A(n_545), .B(n_608), .Y(n_681) );
INVx1_ASAP7_75t_L g688 ( .A(n_545), .Y(n_688) );
NOR2xp33_ASAP7_75t_R g740 ( .A(n_545), .B(n_571), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_545), .B(n_583), .Y(n_744) );
INVx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_552), .Y(n_547) );
AOI32xp33_ASAP7_75t_L g767 ( .A1(n_554), .A2(n_603), .A3(n_768), .B1(n_769), .B2(n_770), .Y(n_767) );
INVx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
INVx2_ASAP7_75t_L g634 ( .A(n_556), .Y(n_634) );
AND2x4_ASAP7_75t_L g653 ( .A(n_556), .B(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_556), .B(n_625), .Y(n_682) );
OR2x2_ASAP7_75t_L g736 ( .A(n_556), .B(n_737), .Y(n_736) );
OR2x2_ASAP7_75t_L g694 ( .A(n_557), .B(n_695), .Y(n_694) );
OR2x2_ASAP7_75t_L g752 ( .A(n_557), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_558), .B(n_571), .Y(n_718) );
AND2x2_ASAP7_75t_L g755 ( .A(n_558), .B(n_721), .Y(n_755) );
INVx2_ASAP7_75t_L g605 ( .A(n_559), .Y(n_605) );
INVx2_ASAP7_75t_L g608 ( .A(n_559), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_559), .B(n_571), .Y(n_628) );
INVx1_ASAP7_75t_L g659 ( .A(n_559), .Y(n_659) );
OR2x2_ASAP7_75t_L g685 ( .A(n_559), .B(n_571), .Y(n_685) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_559), .Y(n_737) );
BUFx3_ASAP7_75t_L g766 ( .A(n_559), .Y(n_766) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g635 ( .A(n_566), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_566), .B(n_653), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_566), .B(n_724), .Y(n_723) );
AND2x4_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_567), .B(n_638), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g667 ( .A1(n_567), .A2(n_634), .B(n_652), .Y(n_667) );
OAI32xp33_ASAP7_75t_L g689 ( .A1(n_568), .A2(n_690), .A3(n_692), .B1(n_694), .B2(n_696), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_568), .B(n_653), .Y(n_762) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g695 ( .A(n_570), .Y(n_695) );
NOR2x1p5_ASAP7_75t_L g765 ( .A(n_570), .B(n_766), .Y(n_765) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x4_ASAP7_75t_L g581 ( .A(n_571), .B(n_582), .Y(n_581) );
AND2x4_ASAP7_75t_SL g603 ( .A(n_571), .B(n_583), .Y(n_603) );
OR2x2_ASAP7_75t_L g607 ( .A(n_571), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g642 ( .A(n_571), .Y(n_642) );
AND2x2_ASAP7_75t_L g660 ( .A(n_571), .B(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g671 ( .A(n_571), .B(n_583), .Y(n_671) );
OR2x2_ASAP7_75t_L g733 ( .A(n_571), .B(n_734), .Y(n_733) );
OR2x2_ASAP7_75t_L g750 ( .A(n_571), .B(n_681), .Y(n_750) );
INVx1_ASAP7_75t_L g782 ( .A(n_571), .Y(n_782) );
OR2x6_ASAP7_75t_L g571 ( .A(n_572), .B(n_578), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_580), .B(n_659), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_581), .B(n_693), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g697 ( .A1(n_581), .A2(n_698), .B1(n_703), .B2(n_705), .C1(n_708), .C2(n_711), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_581), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g725 ( .A(n_581), .B(n_604), .Y(n_725) );
AND2x2_ASAP7_75t_L g687 ( .A(n_582), .B(n_688), .Y(n_687) );
OR2x2_ASAP7_75t_L g702 ( .A(n_582), .B(n_607), .Y(n_702) );
INVx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_583), .B(n_608), .Y(n_640) );
AND2x4_ASAP7_75t_L g661 ( .A(n_583), .B(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g721 ( .A(n_583), .B(n_642), .Y(n_721) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
INVx1_ASAP7_75t_SL g601 ( .A(n_595), .Y(n_601) );
NAND2xp33_ASAP7_75t_SL g770 ( .A(n_595), .B(n_625), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .C(n_602), .Y(n_596) );
INVx2_ASAP7_75t_SL g647 ( .A(n_597), .Y(n_647) );
AND2x2_ASAP7_75t_L g651 ( .A(n_598), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_599), .B(n_647), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_599), .A2(n_637), .B(n_673), .C(n_674), .Y(n_672) );
AND2x2_ASAP7_75t_L g749 ( .A(n_599), .B(n_730), .Y(n_749) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x4_ASAP7_75t_L g648 ( .A(n_603), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g753 ( .A(n_603), .Y(n_753) );
OAI211xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_609), .B(n_616), .C(n_643), .Y(n_606) );
INVx2_ASAP7_75t_L g618 ( .A(n_607), .Y(n_618) );
OR2x2_ASAP7_75t_L g665 ( .A(n_607), .B(n_666), .Y(n_665) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_608), .Y(n_649) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_611), .B(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g703 ( .A(n_611), .B(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_611), .B(n_691), .Y(n_757) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g715 ( .A1(n_613), .A2(n_716), .B1(n_717), .B2(n_719), .C1(n_722), .C2(n_725), .Y(n_715) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_614), .A2(n_679), .B1(n_682), .B2(n_683), .C(n_689), .Y(n_678) );
AND2x2_ASAP7_75t_L g716 ( .A(n_614), .B(n_673), .Y(n_716) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp33_ASAP7_75t_SL g629 ( .A(n_615), .B(n_630), .Y(n_629) );
AOI221x1_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_621), .B1(n_626), .B2(n_629), .C(n_632), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
AND2x2_ASAP7_75t_L g769 ( .A(n_619), .B(n_707), .Y(n_769) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g627 ( .A(n_620), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
OAI32xp33_ASAP7_75t_L g735 ( .A1(n_625), .A2(n_666), .A3(n_736), .B1(n_738), .B2(n_742), .Y(n_735) );
OAI21xp33_ASAP7_75t_SL g754 ( .A1(n_626), .A2(n_755), .B(n_756), .Y(n_754) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B(n_639), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
OR2x2_ASAP7_75t_L g636 ( .A(n_634), .B(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g709 ( .A(n_634), .B(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_638), .A2(n_664), .B1(n_667), .B2(n_668), .C(n_672), .Y(n_663) );
INVx1_ASAP7_75t_L g739 ( .A(n_638), .Y(n_739) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_638), .Y(n_745) );
OR2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_647), .B(n_712), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_655), .B(n_663), .Y(n_650) );
HB1xp67_ASAP7_75t_L g724 ( .A(n_654), .Y(n_724) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_660), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_657), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g676 ( .A(n_659), .Y(n_676) );
INVx1_ASAP7_75t_L g666 ( .A(n_661), .Y(n_666) );
AND2x2_ASAP7_75t_SL g675 ( .A(n_661), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_661), .B(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_661), .B(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
OR2x2_ASAP7_75t_L g680 ( .A(n_671), .B(n_681), .Y(n_680) );
INVx2_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_676), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_678), .B(n_697), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g693 ( .A(n_681), .Y(n_693) );
INVx1_ASAP7_75t_SL g683 ( .A(n_684), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_SL g707 ( .A(n_685), .Y(n_707) );
INVx1_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_687), .B(n_765), .Y(n_764) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_688), .Y(n_701) );
BUFx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_699), .B(n_702), .Y(n_698) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g712 ( .A(n_704), .Y(n_712) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g731 ( .A(n_710), .Y(n_731) );
NOR4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_747), .C(n_758), .D(n_771), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_726), .Y(n_714) );
O2A1O1Ixp33_ASAP7_75t_L g726 ( .A1(n_716), .A2(n_727), .B(n_732), .C(n_735), .Y(n_726) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_729), .B(n_731), .Y(n_728) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_729), .A2(n_739), .B(n_740), .C(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
OAI21xp33_ASAP7_75t_SL g742 ( .A1(n_743), .A2(n_745), .B(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_SL g777 ( .A(n_746), .B(n_778), .Y(n_777) );
OAI221xp5_ASAP7_75t_SL g747 ( .A1(n_748), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_754), .Y(n_747) );
INVx1_ASAP7_75t_SL g751 ( .A(n_749), .Y(n_751) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND3xp33_ASAP7_75t_SL g758 ( .A(n_759), .B(n_760), .C(n_767), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_763), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_774), .B(n_776), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVxp33_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_784), .Y(n_783) );
CKINVDCx11_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_786), .A2(n_788), .B(n_789), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx3_ASAP7_75t_L g816 ( .A(n_793), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
INVx1_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
OAI21x1_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_807), .B(n_810), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2x1_ASAP7_75t_L g807 ( .A(n_800), .B(n_808), .Y(n_807) );
INVxp67_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_L g809 ( .A(n_804), .Y(n_809) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_SL g811 ( .A(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx2_ASAP7_75t_SL g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g822 ( .A(n_815), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g815 ( .A(n_816), .B(n_817), .Y(n_815) );
INVx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
endmodule