module fake_jpeg_31840_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_34),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_33),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

A2O1A1O1Ixp25_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_33),
.B(n_24),
.C(n_18),
.D(n_29),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_29),
.B(n_21),
.C(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_31),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_67),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_43),
.A2(n_28),
.B1(n_32),
.B2(n_27),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_65),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_28),
.B1(n_32),
.B2(n_27),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_19),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_31),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_71),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_75),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_32),
.B1(n_27),
.B2(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_40),
.A2(n_25),
.B1(n_23),
.B2(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_44),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_21),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_23),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_90),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_83),
.B(n_86),
.Y(n_128)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_73),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_51),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

OA21x2_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_41),
.B(n_46),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_62),
.B1(n_79),
.B2(n_55),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_51),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_97),
.C(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_46),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_38),
.B1(n_36),
.B2(n_20),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_102),
.B1(n_6),
.B2(n_7),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_38),
.B1(n_20),
.B2(n_2),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_59),
.B1(n_70),
.B2(n_55),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_80),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_20),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_20),
.C(n_3),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_SL g109 ( 
.A1(n_66),
.A2(n_0),
.B(n_4),
.C(n_6),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_4),
.B(n_6),
.Y(n_115)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_110),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_119),
.B1(n_106),
.B2(n_101),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_115),
.A2(n_89),
.B(n_82),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_90),
.B1(n_88),
.B2(n_84),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_124),
.B1(n_133),
.B2(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_15),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_16),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_127),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_95),
.C(n_87),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_86),
.B(n_12),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_11),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_134),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_59),
.C(n_68),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_101),
.B1(n_109),
.B2(n_83),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_11),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_135),
.B(n_128),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_136),
.A2(n_155),
.B1(n_120),
.B2(n_125),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_138),
.B(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_148),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_93),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_91),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_147),
.B(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_99),
.Y(n_147)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_121),
.CI(n_126),
.CON(n_148),
.SN(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_152),
.B(n_156),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_113),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_131),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_141),
.C(n_148),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_124),
.A2(n_98),
.B1(n_110),
.B2(n_89),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_98),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_115),
.B1(n_111),
.B2(n_119),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_149),
.B1(n_132),
.B2(n_68),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_165),
.C(n_157),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_112),
.B(n_111),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_163),
.A2(n_164),
.B(n_173),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_112),
.B(n_111),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_135),
.C(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_166),
.B(n_151),
.Y(n_176)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_140),
.A2(n_156),
.B1(n_155),
.B2(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_167),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_130),
.B1(n_103),
.B2(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_147),
.A2(n_141),
.B(n_137),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_183),
.B1(n_185),
.B2(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_184),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_173),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_153),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_159),
.C(n_158),
.Y(n_199)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_132),
.B1(n_85),
.B2(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_132),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_104),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_199),
.C(n_179),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_198),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_170),
.B(n_163),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_196),
.B(n_197),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_170),
.B(n_162),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_182),
.A2(n_162),
.B(n_169),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g198 ( 
.A(n_180),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_196),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_177),
.C(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_206),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_175),
.C(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_195),
.B(n_174),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_207),
.B(n_189),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_183),
.C(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_174),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_212),
.C(n_171),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_189),
.C(n_181),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_213),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_167),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_205),
.B(n_181),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_214),
.A2(n_212),
.B(n_8),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_216),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_217),
.B(n_208),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_218),
.A2(n_220),
.B1(n_7),
.B2(n_8),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_7),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_222),
.B(n_8),
.Y(n_223)
);

AOI221xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_9),
.B1(n_58),
.B2(n_62),
.C(n_215),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_62),
.Y(n_225)
);


endmodule