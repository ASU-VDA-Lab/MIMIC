module real_jpeg_8428_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_2),
.A2(n_21),
.B1(n_22),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_3),
.A2(n_21),
.B1(n_22),
.B2(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_10),
.A2(n_21),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_10),
.B(n_21),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_10),
.A2(n_58),
.B1(n_95),
.B2(n_96),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_47),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_73),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_65),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_65),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_51),
.B2(n_64),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_26),
.B1(n_29),
.B2(n_34),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_20),
.A2(n_26),
.B1(n_29),
.B2(n_69),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_27),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_21),
.A2(n_22),
.B1(n_42),
.B2(n_43),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_21),
.B(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_22),
.A2(n_37),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_26),
.A2(n_29),
.B1(n_69),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_27),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_27),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_29),
.B(n_40),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_30),
.B(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_30),
.B(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_30),
.B(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_31),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_45),
.B2(n_46),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_40),
.CON(n_37),
.SN(n_37)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_42),
.B(n_44),
.C(n_45),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_42),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_40),
.B(n_96),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_60),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_58),
.A2(n_79),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_59),
.A2(n_60),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.CI(n_70),
.CON(n_65),
.SN(n_65)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_103),
.B(n_106),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_91),
.B(n_102),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_81),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_90),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_90),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_97),
.B(n_101),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_93),
.B(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_104),
.B(n_105),
.Y(n_106)
);


endmodule