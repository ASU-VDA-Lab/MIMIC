module fake_jpeg_19626_n_29 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_15;

AOI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_12),
.A2(n_8),
.B1(n_7),
.B2(n_13),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_5),
.Y(n_17)
);

AOI32xp33_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_11),
.A3(n_10),
.B1(n_9),
.B2(n_3),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_15),
.B(n_6),
.C(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_19),
.A2(n_20),
.B1(n_14),
.B2(n_17),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_14),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_15),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_24),
.B(n_20),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_16),
.B(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_16),
.Y(n_28)
);

OA21x2_ASAP7_75t_L g29 ( 
.A1(n_28),
.A2(n_24),
.B(n_6),
.Y(n_29)
);


endmodule