module real_jpeg_19131_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_17;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_73;
wire n_65;
wire n_35;
wire n_33;
wire n_50;
wire n_38;
wire n_29;
wire n_55;
wire n_69;
wire n_49;
wire n_10;
wire n_58;
wire n_31;
wire n_52;
wire n_67;
wire n_63;
wire n_12;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_72;
wire n_28;
wire n_44;
wire n_60;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_11;
wire n_14;
wire n_71;
wire n_51;
wire n_45;
wire n_25;
wire n_47;
wire n_61;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_70;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_56;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_0),
.B(n_4),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_7),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_8),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_1),
.A2(n_14),
.B1(n_15),
.B2(n_23),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g56 ( 
.A(n_3),
.B(n_57),
.CON(n_56),
.SN(n_56)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_42),
.Y(n_46)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_7),
.Y(n_61)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_50),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_29),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_27),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_24),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_19),
.B(n_21),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_18),
.Y(n_16)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_20),
.B(n_21),
.C(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_17),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_25),
.A2(n_26),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_26),
.B(n_41),
.C(n_42),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_68),
.B(n_73),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_52),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g31 ( 
.A1(n_32),
.A2(n_43),
.B(n_51),
.Y(n_31)
);

NOR3xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_53),
.C(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_38),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.C(n_37),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_48),
.C(n_50),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_47),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_63),
.B(n_67),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_59),
.Y(n_55)
);

BUFx24_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);


endmodule