module fake_jpeg_2400_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_6),
.B(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_2),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_18),
.B(n_13),
.C(n_19),
.Y(n_36)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_2),
.B(n_3),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_25),
.B(n_26),
.Y(n_35)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_4),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_9),
.A2(n_12),
.B1(n_13),
.B2(n_11),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_13),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_29),
.Y(n_44)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_11),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_34),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_14),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_35),
.B(n_30),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_26),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_34),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.C(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_44),
.B(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_28),
.B(n_32),
.C(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_52),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_51),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_53),
.B(n_48),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_56),
.C(n_55),
.Y(n_58)
);


endmodule