module real_jpeg_26237_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_83;
wire n_166;
wire n_176;
wire n_286;
wire n_300;
wire n_292;
wire n_249;
wire n_215;
wire n_221;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_299;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_290;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_285;
wire n_45;
wire n_172;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_300),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_2),
.B(n_301),
.Y(n_300)
);

BUFx8_ASAP7_75t_L g73 ( 
.A(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_4),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_9),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_6),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_6),
.A2(n_44),
.B1(n_73),
.B2(n_74),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_6),
.B(n_29),
.C(n_32),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_6),
.B(n_30),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_6),
.B(n_51),
.C(n_54),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_70),
.C(n_73),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_6),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_6),
.B(n_101),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_6),
.B(n_63),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_60),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_8),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_8),
.A2(n_60),
.B1(n_73),
.B2(n_74),
.Y(n_190)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_10),
.A2(n_21),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_10),
.A2(n_35),
.B1(n_54),
.B2(n_55),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_35),
.B1(n_73),
.B2(n_74),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_11),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_11),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_11),
.A2(n_24),
.B1(n_54),
.B2(n_55),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_11),
.A2(n_24),
.B1(n_73),
.B2(n_74),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_13),
.Y(n_127)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_293),
.B(n_297),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_76),
.B(n_292),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_18),
.B(n_38),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_18),
.B(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_18),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_25),
.B1(n_30),
.B2(n_34),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_41),
.B(n_42),
.Y(n_40)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_23),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_25),
.A2(n_30),
.B1(n_43),
.B2(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_27),
.B(n_186),
.Y(n_185)
);

AO22x1_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_32),
.B(n_220),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_34),
.B(n_296),
.Y(n_295)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_39),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_39),
.B(n_290),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_45),
.CI(n_56),
.CON(n_39),
.SN(n_39)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_42),
.B(n_59),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_53),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_48),
.A2(n_53),
.B(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_49),
.A2(n_63),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_49),
.B(n_106),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OA22x2_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_53),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_105),
.B(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_54),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_54),
.B(n_233),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_64),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_SL g123 ( 
.A(n_57),
.B(n_124),
.C(n_131),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_57),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_57),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_57),
.A2(n_131),
.B1(n_132),
.B2(n_145),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_57),
.A2(n_103),
.B1(n_145),
.B2(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_57),
.B(n_103),
.C(n_183),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_61),
.A2(n_64),
.B1(n_113),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_61),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_109),
.C(n_114),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_75),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_66),
.B(n_91),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_68),
.A2(n_91),
.B1(n_101),
.B2(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_72),
.A2(n_90),
.B(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_73),
.B(n_238),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_289),
.B(n_291),
.Y(n_76)
);

OAI211xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_133),
.B(n_147),
.C(n_288),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_118),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_79),
.B(n_118),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_96),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_98),
.C(n_107),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_92),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_81),
.A2(n_92),
.B1(n_93),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_81),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_81),
.A2(n_88),
.B1(n_121),
.B2(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

INVxp33_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_83),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_86),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_85),
.A2(n_126),
.B(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_87),
.B(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_88),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_94),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_107),
.B2(n_108),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_99),
.B(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_103),
.B(n_204),
.C(n_206),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_103),
.A2(n_194),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_109),
.A2(n_110),
.B1(n_141),
.B2(n_146),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_109),
.B(n_131),
.C(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_109),
.A2(n_110),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_109),
.A2(n_110),
.B1(n_165),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_157),
.C(n_165),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_110),
.B(n_137),
.C(n_141),
.Y(n_290)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_123),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_122),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_125),
.A2(n_128),
.B1(n_129),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_125),
.Y(n_279)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_128),
.A2(n_129),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_128),
.A2(n_129),
.B1(n_217),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_129),
.B(n_211),
.C(n_217),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_129),
.B(n_188),
.C(n_250),
.Y(n_254)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_131),
.A2(n_132),
.B1(n_179),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_131),
.A2(n_132),
.B1(n_163),
.B2(n_176),
.Y(n_256)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_132),
.B(n_163),
.C(n_257),
.Y(n_260)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_148),
.C(n_149),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_135),
.B(n_136),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_169),
.B(n_287),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_167),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_151),
.B(n_167),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_152),
.B(n_154),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_156),
.B(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_157),
.A2(n_158),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_163),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_159),
.A2(n_163),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_161),
.A2(n_190),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_163),
.A2(n_176),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_163),
.B(n_234),
.Y(n_246)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_165),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_282),
.B(n_286),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_207),
.B(n_268),
.C(n_281),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_196),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_172),
.B(n_196),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_182),
.B2(n_195),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_175),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_175),
.B(n_181),
.C(n_195),
.Y(n_269)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_187),
.A2(n_188),
.B1(n_248),
.B2(n_249),
.Y(n_247)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_188),
.B(n_242),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_202),
.C(n_203),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_197),
.A2(n_198),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_203),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_206),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_204),
.B(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_267),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_226),
.B(n_266),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_223),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_210),
.B(n_223),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_212),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_216),
.B(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_217),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_259),
.B(n_265),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_253),
.B(n_258),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_245),
.B(n_252),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_235),
.B(n_244),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_232),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_241),
.B(n_243),
.Y(n_235)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_246),
.B(n_247),
.Y(n_252)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_250),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_261),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_262),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_270),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_280),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_277),
.B2(n_278),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_278),
.C(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);


endmodule