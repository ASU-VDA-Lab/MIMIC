module fake_jpeg_3208_n_195 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_195);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_195;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_41),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_59),
.Y(n_83)
);

BUFx16f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_78),
.Y(n_81)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_68),
.B1(n_56),
.B2(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_87),
.B1(n_75),
.B2(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_73),
.A2(n_57),
.B1(n_53),
.B2(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_94),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_102),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_50),
.B(n_62),
.C(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_71),
.B1(n_75),
.B2(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_99),
.A2(n_91),
.B1(n_88),
.B2(n_55),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_61),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_75),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_101),
.B(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_81),
.B(n_69),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_52),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_105),
.Y(n_112)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_78),
.B1(n_53),
.B2(n_57),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_92),
.B1(n_91),
.B2(n_101),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_63),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_94),
.B1(n_100),
.B2(n_98),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_117),
.B1(n_120),
.B2(n_124),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_2),
.Y(n_142)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_95),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_65),
.B1(n_60),
.B2(n_66),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_21),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_65),
.B(n_2),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_3),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_0),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_22),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_144),
.Y(n_162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_109),
.B(n_111),
.C(n_110),
.D(n_126),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_10),
.B(n_11),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_146),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_20),
.B1(n_47),
.B2(n_46),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_136),
.B1(n_145),
.B2(n_6),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_49),
.B1(n_45),
.B2(n_43),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_42),
.C(n_39),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_148),
.C(n_19),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_3),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_115),
.B(n_4),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_4),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_5),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_27),
.C(n_26),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_24),
.Y(n_149)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_23),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_129),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_154),
.Y(n_167)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_165),
.B1(n_152),
.B2(n_164),
.C(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_157),
.B(n_160),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_139),
.Y(n_158)
);

AOI21x1_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_143),
.B(n_148),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_131),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_163),
.C(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_164),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_8),
.C(n_9),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_166),
.A2(n_140),
.B1(n_15),
.B2(n_16),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_152),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_174),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_136),
.C(n_134),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_158),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_162),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_156),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_175),
.B(n_176),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_183),
.C(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_179),
.Y(n_187)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

AOI31xp67_ASAP7_75t_L g185 ( 
.A1(n_180),
.A2(n_150),
.A3(n_170),
.B(n_172),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_184),
.B(n_185),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_168),
.C(n_150),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_178),
.C(n_181),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_190),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_187),
.A2(n_177),
.B1(n_182),
.B2(n_155),
.Y(n_190)
);

AOI21x1_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_188),
.B(n_174),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_13),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_13),
.B(n_17),
.Y(n_194)
);

XNOR2x2_ASAP7_75t_SL g195 ( 
.A(n_194),
.B(n_18),
.Y(n_195)
);


endmodule