module fake_ariane_1472_n_644 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_644);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_644;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_610;
wire n_205;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_139;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_166;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_330;
wire n_400;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_588;
wire n_638;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_617;
wire n_616;
wire n_630;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_641;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_544;
wire n_540;
wire n_216;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_375;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_531;

BUFx3_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_53),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_83),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_38),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_12),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_13),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_21),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_43),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_26),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_70),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_69),
.Y(n_149)
);

BUFx10_ASAP7_75t_L g150 ( 
.A(n_103),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_60),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_44),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_9),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_86),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_87),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_24),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_81),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_5),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_62),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_47),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_55),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_32),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_57),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_75),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_108),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_106),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_25),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_19),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_80),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_27),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_30),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_65),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_63),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_109),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_15),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_50),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_124),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_28),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_48),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_33),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_128),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_77),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_20),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_82),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_76),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_104),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_131),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_107),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_133),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_135),
.A2(n_0),
.B(n_1),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_2),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

OAI21x1_ASAP7_75t_L g211 ( 
.A1(n_144),
.A2(n_68),
.B(n_126),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_151),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_143),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_162),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_151),
.Y(n_217)
);

AOI22x1_ASAP7_75t_SL g218 ( 
.A1(n_195),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_146),
.Y(n_219)
);

AND2x4_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_7),
.Y(n_220)
);

OAI22x1_ASAP7_75t_SL g221 ( 
.A1(n_156),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_136),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_151),
.Y(n_224)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_142),
.A2(n_11),
.B(n_12),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_176),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

AND2x4_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_11),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_150),
.Y(n_229)
);

OAI22x1_ASAP7_75t_R g230 ( 
.A1(n_200),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_230)
);

AND2x4_ASAP7_75t_L g231 ( 
.A(n_144),
.B(n_14),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_150),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_147),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_169),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_152),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_153),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_147),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_189),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

OA21x2_ASAP7_75t_L g245 ( 
.A1(n_170),
.A2(n_23),
.B(n_29),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_171),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_175),
.B(n_34),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_179),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_243),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

NOR2xp67_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_137),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_243),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_138),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_168),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_234),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_213),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_210),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_229),
.Y(n_268)
);

NAND2xp33_ASAP7_75t_R g269 ( 
.A(n_232),
.B(n_186),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_237),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_R g273 ( 
.A(n_222),
.B(n_140),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_219),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_227),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_231),
.B(n_201),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_223),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_219),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_230),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_240),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_204),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_236),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_204),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_206),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_206),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_235),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_235),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_208),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_208),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_236),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_210),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_218),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_R g300 ( 
.A(n_244),
.B(n_145),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_220),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_252),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_251),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_247),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_257),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_286),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_281),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_249),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_209),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_247),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_277),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_284),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_220),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_256),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_244),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_270),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_274),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_287),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_301),
.B(n_231),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_261),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_263),
.Y(n_328)
);

AO221x1_ASAP7_75t_L g329 ( 
.A1(n_269),
.A2(n_215),
.B1(n_221),
.B2(n_241),
.C(n_193),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_269),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_247),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_273),
.B(n_228),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_209),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_273),
.B(n_228),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_276),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_266),
.Y(n_338)
);

NAND2x1_ASAP7_75t_L g339 ( 
.A(n_266),
.B(n_233),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_294),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_278),
.B(n_239),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_279),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_264),
.B(n_239),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_268),
.B(n_246),
.Y(n_347)
);

NOR3xp33_ASAP7_75t_SL g348 ( 
.A(n_262),
.B(n_185),
.C(n_154),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_271),
.B(n_246),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_300),
.B(n_236),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_300),
.B(n_253),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_298),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_260),
.B(n_203),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_254),
.B(n_216),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_272),
.B(n_149),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_292),
.B(n_238),
.Y(n_357)
);

OR2x2_ASAP7_75t_SL g358 ( 
.A(n_283),
.B(n_207),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_255),
.B(n_238),
.Y(n_359)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_250),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_250),
.Y(n_361)
);

AO221x1_ASAP7_75t_L g362 ( 
.A1(n_299),
.A2(n_196),
.B1(n_198),
.B2(n_238),
.C(n_207),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_274),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_252),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_281),
.Y(n_365)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_282),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_251),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_319),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_310),
.B(n_155),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_307),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_334),
.A2(n_238),
.B1(n_225),
.B2(n_207),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_302),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_318),
.A2(n_225),
.B1(n_177),
.B2(n_245),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_311),
.B(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_306),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_333),
.A2(n_245),
.B1(n_184),
.B2(n_183),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_331),
.B(n_158),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_364),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_305),
.B(n_160),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_303),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_321),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_L g383 ( 
.A(n_366),
.B(n_161),
.Y(n_383)
);

BUFx8_ASAP7_75t_SL g384 ( 
.A(n_322),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_163),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_362),
.A2(n_245),
.B1(n_190),
.B2(n_188),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_324),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_314),
.B(n_164),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_320),
.Y(n_389)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_316),
.B(n_211),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_314),
.B(n_166),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_332),
.B(n_167),
.Y(n_393)
);

OR2x6_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_210),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_325),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_315),
.B(n_172),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_335),
.A2(n_192),
.B(n_174),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_365),
.B(n_173),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_309),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_332),
.B(n_178),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_330),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_348),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_329),
.A2(n_197),
.B1(n_187),
.B2(n_194),
.Y(n_405)
);

A2O1A1Ixp33_ASAP7_75t_L g406 ( 
.A1(n_312),
.A2(n_199),
.B(n_182),
.C(n_212),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_342),
.B(n_224),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_340),
.B(n_224),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g409 ( 
.A(n_351),
.B(n_224),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_355),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_367),
.Y(n_411)
);

OR2x2_ASAP7_75t_SL g412 ( 
.A(n_357),
.B(n_224),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_338),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g415 ( 
.A1(n_323),
.A2(n_217),
.B(n_212),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_326),
.A2(n_217),
.B1(n_212),
.B2(n_37),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_357),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_340),
.B(n_217),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_347),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_360),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_344),
.B(n_217),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_350),
.A2(n_212),
.B(n_36),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g425 ( 
.A(n_359),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_358),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_341),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_353),
.B(n_127),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_366),
.B(n_41),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_313),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_343),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_304),
.Y(n_432)
);

O2A1O1Ixp33_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_354),
.B(n_317),
.C(n_356),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_410),
.Y(n_434)
);

A2O1A1Ixp33_ASAP7_75t_L g435 ( 
.A1(n_428),
.A2(n_339),
.B(n_349),
.C(n_344),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_427),
.B(n_363),
.Y(n_436)
);

O2A1O1Ixp33_ASAP7_75t_L g437 ( 
.A1(n_389),
.A2(n_345),
.B(n_366),
.C(n_363),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_372),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_363),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g440 ( 
.A1(n_383),
.A2(n_337),
.B(n_336),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_SL g441 ( 
.A(n_404),
.B(n_366),
.C(n_337),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_380),
.A2(n_337),
.B(n_336),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_374),
.B(n_366),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_375),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_426),
.A2(n_336),
.B1(n_328),
.B2(n_46),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_420),
.B(n_328),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_384),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_377),
.A2(n_328),
.B(n_45),
.C(n_49),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_429),
.A2(n_42),
.B(n_51),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_414),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_379),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_385),
.A2(n_52),
.B(n_56),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_382),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_388),
.A2(n_58),
.B(n_59),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_392),
.A2(n_401),
.B1(n_393),
.B2(n_418),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_377),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_67),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_SL g462 ( 
.A1(n_370),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_462)
);

OR2x2_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_79),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_408),
.A2(n_85),
.B(n_88),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_408),
.A2(n_89),
.B(n_91),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_405),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_387),
.B(n_92),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_395),
.B(n_93),
.Y(n_469)
);

NOR3xp33_ASAP7_75t_SL g470 ( 
.A(n_369),
.B(n_94),
.C(n_95),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_416),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_419),
.A2(n_96),
.B(n_97),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_391),
.B(n_98),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_474),
.Y(n_477)
);

CKINVDCx6p67_ASAP7_75t_R g478 ( 
.A(n_448),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_458),
.Y(n_479)
);

OR3x4_ASAP7_75t_SL g480 ( 
.A(n_467),
.B(n_405),
.C(n_426),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_434),
.Y(n_481)
);

AO21x2_ASAP7_75t_L g482 ( 
.A1(n_449),
.A2(n_373),
.B(n_429),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_438),
.Y(n_483)
);

BUFx2_ASAP7_75t_R g484 ( 
.A(n_439),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_459),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_465),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

NAND2x1p5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_398),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_461),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_443),
.A2(n_457),
.B(n_468),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_445),
.A2(n_378),
.B1(n_399),
.B2(n_394),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_443),
.A2(n_373),
.B(n_417),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_446),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_453),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_468),
.A2(n_406),
.B(n_376),
.Y(n_495)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_450),
.A2(n_442),
.B(n_464),
.Y(n_496)
);

AOI22x1_ASAP7_75t_L g497 ( 
.A1(n_454),
.A2(n_430),
.B1(n_415),
.B2(n_424),
.Y(n_497)
);

AO21x2_ASAP7_75t_L g498 ( 
.A1(n_469),
.A2(n_417),
.B(n_422),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_453),
.Y(n_499)
);

BUFx5_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_371),
.B(n_386),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_461),
.Y(n_502)
);

INVx3_ASAP7_75t_SL g503 ( 
.A(n_475),
.Y(n_503)
);

OR3x4_ASAP7_75t_SL g504 ( 
.A(n_470),
.B(n_397),
.C(n_394),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_469),
.A2(n_411),
.B(n_400),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_475),
.Y(n_506)
);

AOI22xp33_ASAP7_75t_L g507 ( 
.A1(n_480),
.A2(n_460),
.B1(n_471),
.B2(n_451),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_500),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_412),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_485),
.Y(n_511)
);

CKINVDCx11_ASAP7_75t_R g512 ( 
.A(n_478),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_500),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_496),
.A2(n_472),
.B(n_456),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_502),
.A2(n_460),
.B1(n_476),
.B2(n_455),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_489),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_502),
.A2(n_452),
.B1(n_463),
.B2(n_436),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_490),
.A2(n_390),
.B(n_435),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_496),
.A2(n_440),
.B(n_437),
.Y(n_519)
);

CKINVDCx6p67_ASAP7_75t_R g520 ( 
.A(n_478),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_486),
.B(n_398),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_483),
.B(n_403),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_500),
.Y(n_523)
);

CKINVDCx11_ASAP7_75t_R g524 ( 
.A(n_503),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_499),
.B(n_447),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_500),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_480),
.A2(n_381),
.B1(n_441),
.B2(n_409),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_499),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_500),
.B(n_433),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_477),
.A2(n_493),
.B1(n_492),
.B2(n_482),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_500),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_495),
.A2(n_390),
.B(n_473),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_484),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_488),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_515),
.A2(n_491),
.B(n_488),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_509),
.B(n_503),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_511),
.B(n_477),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_521),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_510),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_493),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_500),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_R g543 ( 
.A(n_524),
.B(n_533),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_522),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_521),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_R g547 ( 
.A(n_512),
.B(n_487),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_525),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_525),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_516),
.B(n_500),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_487),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_486),
.Y(n_552)
);

NAND3xp33_ASAP7_75t_SL g553 ( 
.A(n_527),
.B(n_505),
.C(n_488),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_506),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_520),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_517),
.B(n_529),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_R g557 ( 
.A(n_513),
.B(n_506),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_523),
.B(n_506),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_518),
.A2(n_492),
.B1(n_482),
.B2(n_498),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_521),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_521),
.B(n_494),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_529),
.A2(n_482),
.B(n_492),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_518),
.A2(n_498),
.B1(n_501),
.B2(n_391),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_508),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_544),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_534),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_544),
.B(n_526),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_538),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_545),
.B(n_526),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_538),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_548),
.Y(n_571)
);

BUFx2_ASAP7_75t_L g572 ( 
.A(n_557),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_508),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_562),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_534),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_536),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_554),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_562),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_555),
.B(n_531),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_537),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_542),
.B(n_526),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_541),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_558),
.B(n_557),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_535),
.B(n_531),
.Y(n_584)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_556),
.B(n_530),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_534),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_551),
.B(n_518),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_565),
.B(n_556),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_565),
.B(n_564),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_582),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_582),
.B(n_540),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_576),
.B(n_539),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_576),
.B(n_539),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_577),
.B(n_558),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_587),
.B(n_550),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_559),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_572),
.B(n_560),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_571),
.B(n_558),
.Y(n_599)
);

OAI221xp5_ASAP7_75t_L g600 ( 
.A1(n_585),
.A2(n_559),
.B1(n_552),
.B2(n_532),
.C(n_563),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_572),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_577),
.B(n_561),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_598),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_589),
.B(n_579),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_594),
.B(n_566),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_595),
.B(n_581),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_601),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_591),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_588),
.B(n_580),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_583),
.Y(n_610)
);

NAND4xp75_ASAP7_75t_SL g611 ( 
.A(n_604),
.B(n_543),
.C(n_555),
.D(n_583),
.Y(n_611)
);

OAI322xp33_ASAP7_75t_L g612 ( 
.A1(n_609),
.A2(n_588),
.A3(n_589),
.B1(n_596),
.B2(n_599),
.C1(n_585),
.C2(n_600),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_610),
.B(n_593),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_608),
.Y(n_614)
);

AOI33xp33_ASAP7_75t_L g615 ( 
.A1(n_603),
.A2(n_592),
.A3(n_569),
.B1(n_567),
.B2(n_563),
.B3(n_590),
.Y(n_615)
);

OAI322xp33_ASAP7_75t_L g616 ( 
.A1(n_606),
.A2(n_596),
.A3(n_600),
.B1(n_573),
.B2(n_597),
.C1(n_569),
.C2(n_570),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_604),
.B(n_567),
.Y(n_617)
);

NOR2x1_ASAP7_75t_L g618 ( 
.A(n_611),
.B(n_584),
.Y(n_618)
);

OAI21xp33_ASAP7_75t_SL g619 ( 
.A1(n_611),
.A2(n_607),
.B(n_605),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_614),
.A2(n_605),
.B1(n_584),
.B2(n_553),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g621 ( 
.A(n_617),
.B(n_584),
.Y(n_621)
);

O2A1O1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_612),
.A2(n_584),
.B(n_532),
.C(n_462),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_620),
.A2(n_613),
.B1(n_616),
.B2(n_575),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_621),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_619),
.B(n_615),
.Y(n_625)
);

AOI222xp33_ASAP7_75t_L g626 ( 
.A1(n_618),
.A2(n_570),
.B1(n_578),
.B2(n_574),
.C1(n_568),
.C2(n_501),
.Y(n_626)
);

AOI221xp5_ASAP7_75t_L g627 ( 
.A1(n_622),
.A2(n_543),
.B1(n_547),
.B2(n_574),
.C(n_578),
.Y(n_627)
);

OAI21xp33_ASAP7_75t_L g628 ( 
.A1(n_625),
.A2(n_547),
.B(n_514),
.Y(n_628)
);

OAI322xp33_ASAP7_75t_L g629 ( 
.A1(n_623),
.A2(n_575),
.A3(n_566),
.B1(n_586),
.B2(n_568),
.C1(n_497),
.C2(n_504),
.Y(n_629)
);

NOR2x1_ASAP7_75t_L g630 ( 
.A(n_627),
.B(n_575),
.Y(n_630)
);

AOI211xp5_ASAP7_75t_L g631 ( 
.A1(n_628),
.A2(n_624),
.B(n_626),
.C(n_514),
.Y(n_631)
);

NOR3x1_ASAP7_75t_L g632 ( 
.A(n_629),
.B(n_519),
.C(n_504),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_631),
.B(n_630),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_633),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_634),
.Y(n_635)
);

AOI322xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_632),
.A3(n_518),
.B1(n_498),
.B2(n_407),
.C1(n_566),
.C2(n_586),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_636),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_637),
.A2(n_546),
.B1(n_586),
.B2(n_398),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_638),
.A2(n_391),
.B(n_519),
.Y(n_639)
);

HB1xp67_ASAP7_75t_L g640 ( 
.A(n_639),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_99),
.B(n_100),
.Y(n_641)
);

NAND2x1p5_ASAP7_75t_SL g642 ( 
.A(n_641),
.B(n_101),
.Y(n_642)
);

AOI221xp5_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_110),
.B1(n_111),
.B2(n_114),
.C(n_118),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_643),
.A2(n_546),
.B1(n_120),
.B2(n_123),
.Y(n_644)
);


endmodule