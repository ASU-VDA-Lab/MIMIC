module fake_jpeg_12706_n_590 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_590);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_590;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_56),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_57),
.B(n_58),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_23),
.B(n_18),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_60),
.B(n_64),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_61),
.B(n_70),
.Y(n_115)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_68),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_72),
.B(n_76),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g148 ( 
.A(n_75),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_17),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_17),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_92),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_91),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_32),
.B(n_17),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_97),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_94),
.Y(n_179)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_16),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_36),
.Y(n_157)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_29),
.Y(n_99)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_99),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g172 ( 
.A(n_102),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_22),
.Y(n_103)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_28),
.Y(n_108)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_25),
.Y(n_112)
);

INVx8_ASAP7_75t_SL g134 ( 
.A(n_112),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_100),
.A2(n_36),
.B1(n_38),
.B2(n_47),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_127),
.A2(n_51),
.B1(n_52),
.B2(n_50),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_57),
.A2(n_54),
.B(n_47),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_128),
.B(n_133),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_140),
.B(n_151),
.Y(n_234)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_149),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_83),
.Y(n_151)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_154),
.Y(n_215)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_89),
.Y(n_155)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_155),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_75),
.Y(n_180)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_74),
.Y(n_158)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

NAND2x1_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_54),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

CKINVDCx9p33_ASAP7_75t_R g165 ( 
.A(n_102),
.Y(n_165)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_61),
.B(n_37),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_166),
.B(n_49),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_94),
.Y(n_190)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_180),
.B(n_225),
.Y(n_256)
);

NAND3xp33_ASAP7_75t_L g295 ( 
.A(n_181),
.B(n_239),
.C(n_241),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_52),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_196),
.Y(n_251)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_183),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_130),
.A2(n_68),
.B1(n_108),
.B2(n_107),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_184),
.A2(n_216),
.B1(n_178),
.B2(n_160),
.Y(n_283)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_138),
.Y(n_186)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_187),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_115),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_188),
.B(n_197),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_190),
.Y(n_246)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_191),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_192),
.Y(n_299)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_51),
.Y(n_196)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_198),
.Y(n_280)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_199),
.Y(n_257)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_200),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_94),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_201),
.B(n_204),
.Y(n_275)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_202),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_125),
.B(n_38),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_143),
.Y(n_205)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_205),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_132),
.Y(n_207)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_208),
.Y(n_284)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_209),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_211),
.Y(n_282)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_212),
.Y(n_292)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_213),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_50),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_224),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_137),
.A2(n_103),
.B1(n_106),
.B2(n_77),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_148),
.B(n_111),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_217),
.B(n_221),
.Y(n_271)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

BUFx24_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_177),
.B(n_113),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_219),
.B(n_223),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_233),
.Y(n_250)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_123),
.B(n_42),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_141),
.B(n_48),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g225 ( 
.A(n_126),
.B(n_42),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_127),
.A2(n_88),
.B1(n_63),
.B2(n_79),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_226),
.A2(n_236),
.B1(n_168),
.B2(n_163),
.Y(n_274)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_174),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_229),
.Y(n_261)
);

INVx11_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_161),
.B(n_46),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_231),
.B(n_232),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_164),
.B(n_46),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_156),
.Y(n_233)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_146),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_122),
.A2(n_73),
.B1(n_78),
.B2(n_69),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_172),
.B(n_62),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_237),
.B(n_238),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_172),
.B(n_101),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_118),
.B(n_35),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_124),
.B(n_35),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_167),
.A2(n_56),
.B1(n_59),
.B2(n_30),
.Y(n_242)
);

OAI22x1_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_134),
.B1(n_156),
.B2(n_159),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g243 ( 
.A(n_146),
.B(n_96),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_217),
.C(n_210),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_245),
.B(n_265),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_167),
.C(n_148),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_247),
.B(n_254),
.C(n_294),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_249),
.A2(n_176),
.B1(n_65),
.B2(n_3),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_180),
.B(n_188),
.C(n_243),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_259),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_228),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_262),
.B(n_276),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_226),
.A2(n_91),
.B1(n_86),
.B2(n_82),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_146),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_267),
.B(n_268),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_234),
.B(n_153),
.Y(n_268)
);

O2A1O1Ixp33_ASAP7_75t_L g269 ( 
.A1(n_203),
.A2(n_153),
.B(n_116),
.C(n_138),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_269),
.A2(n_187),
.B(n_198),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_274),
.A2(n_277),
.B1(n_283),
.B2(n_53),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_184),
.A2(n_120),
.B1(n_121),
.B2(n_160),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_SL g278 ( 
.A(n_243),
.B(n_171),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_278),
.A2(n_1),
.B(n_3),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_179),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_286),
.B(n_293),
.Y(n_334)
);

OA22x2_ASAP7_75t_L g289 ( 
.A1(n_236),
.A2(n_34),
.B1(n_40),
.B2(n_49),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_297),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_212),
.B(n_185),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_291),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_193),
.B(n_121),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_230),
.B(n_222),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_240),
.B(n_99),
.Y(n_294)
);

OA22x2_ASAP7_75t_L g297 ( 
.A1(n_216),
.A2(n_40),
.B1(n_41),
.B2(n_48),
.Y(n_297)
);

AO21x2_ASAP7_75t_L g298 ( 
.A1(n_242),
.A2(n_178),
.B(n_80),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_235),
.B1(n_186),
.B2(n_199),
.Y(n_305)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

INVx13_ASAP7_75t_L g384 ( 
.A(n_300),
.Y(n_384)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_263),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_301),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_253),
.B(n_258),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_302),
.B(n_311),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_298),
.A2(n_227),
.B1(n_202),
.B2(n_221),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_303),
.A2(n_313),
.B1(n_320),
.B2(n_323),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_304),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_305),
.A2(n_313),
.B1(n_320),
.B2(n_303),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_206),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_330),
.C(n_346),
.Y(n_356)
);

AND2x2_ASAP7_75t_SL g309 ( 
.A(n_245),
.B(n_215),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_315),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_208),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_319),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_253),
.B(n_205),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_275),
.B(n_209),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_312),
.B(n_318),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_298),
.A2(n_233),
.B1(n_229),
.B2(n_211),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_257),
.Y(n_314)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_345),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_218),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_253),
.B(n_191),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_298),
.A2(n_207),
.B1(n_195),
.B2(n_192),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_322),
.A2(n_328),
.B1(n_342),
.B2(n_344),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_298),
.A2(n_256),
.B1(n_260),
.B2(n_283),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_247),
.A2(n_176),
.B1(n_53),
.B2(n_220),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_324),
.A2(n_336),
.B(n_296),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_251),
.B(n_41),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_325),
.B(n_331),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_278),
.A2(n_53),
.B(n_220),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_326),
.A2(n_248),
.B(n_296),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_264),
.B(n_0),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_246),
.B(n_0),
.Y(n_331)
);

INVx5_ASAP7_75t_SL g332 ( 
.A(n_269),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_265),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_280),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_337),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_14),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_340),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_271),
.B(n_3),
.Y(n_340)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_252),
.Y(n_341)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_271),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_265),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_252),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_266),
.B(n_279),
.Y(n_346)
);

INVx6_ASAP7_75t_SL g347 ( 
.A(n_280),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_347),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_255),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_348),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_L g349 ( 
.A1(n_297),
.A2(n_5),
.B(n_7),
.C(n_8),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_5),
.Y(n_378)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_270),
.Y(n_350)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g352 ( 
.A(n_329),
.B(n_250),
.C(n_257),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_352),
.B(n_373),
.C(n_393),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_332),
.A2(n_297),
.B1(n_289),
.B2(n_287),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_355),
.B(n_360),
.Y(n_398)
);

BUFx24_ASAP7_75t_SL g358 ( 
.A(n_327),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_327),
.Y(n_405)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_332),
.A2(n_297),
.B1(n_289),
.B2(n_287),
.Y(n_360)
);

AOI32xp33_ASAP7_75t_L g364 ( 
.A1(n_302),
.A2(n_261),
.A3(n_282),
.B1(n_249),
.B2(n_284),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_364),
.A2(n_372),
.B(n_378),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_333),
.A2(n_265),
.B1(n_289),
.B2(n_272),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_367),
.B(n_375),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_348),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_370),
.B(n_335),
.Y(n_407)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_307),
.B(n_284),
.C(n_273),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_322),
.A2(n_272),
.B1(n_244),
.B2(n_281),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_317),
.B(n_263),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_379),
.B(n_383),
.Y(n_428)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_381),
.B(n_311),
.C(n_306),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_308),
.A2(n_244),
.B1(n_281),
.B2(n_299),
.Y(n_383)
);

OAI32xp33_ASAP7_75t_L g388 ( 
.A1(n_349),
.A2(n_273),
.A3(n_288),
.B1(n_299),
.B2(n_248),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_392),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_323),
.A2(n_288),
.B1(n_9),
.B2(n_10),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_389),
.A2(n_344),
.B1(n_342),
.B2(n_340),
.Y(n_406)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_343),
.Y(n_391)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_308),
.B(n_7),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_329),
.B(n_9),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_353),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_399),
.B(n_403),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_368),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_401),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_352),
.B(n_309),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_409),
.C(n_424),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_381),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_363),
.Y(n_404)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_404),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_405),
.B(n_408),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_414),
.B1(n_321),
.B2(n_375),
.Y(n_453)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_334),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_309),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_363),
.Y(n_410)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_386),
.B(n_334),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_411),
.B(n_418),
.Y(n_463)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_412),
.Y(n_459)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_391),
.Y(n_415)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_379),
.Y(n_416)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_416),
.Y(n_439)
);

INVx13_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_417),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_351),
.B(n_325),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_369),
.A2(n_319),
.B1(n_316),
.B2(n_321),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_419),
.A2(n_374),
.B1(n_367),
.B2(n_336),
.Y(n_434)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

OA22x2_ASAP7_75t_SL g421 ( 
.A1(n_376),
.A2(n_321),
.B1(n_336),
.B2(n_316),
.Y(n_421)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_421),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_377),
.B(n_361),
.Y(n_422)
);

NOR2x1_ASAP7_75t_L g466 ( 
.A(n_422),
.B(n_430),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_377),
.B(n_335),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_429),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_373),
.B(n_310),
.C(n_316),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_368),
.A2(n_326),
.B(n_338),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_425),
.Y(n_460)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_384),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g438 ( 
.A(n_426),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_330),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_362),
.Y(n_431)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_432),
.A2(n_369),
.B1(n_416),
.B2(n_372),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_433),
.A2(n_442),
.B1(n_449),
.B2(n_406),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_434),
.A2(n_453),
.B1(n_461),
.B2(n_422),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_432),
.A2(n_389),
.B1(n_376),
.B2(n_374),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_411),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_447),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g447 ( 
.A(n_399),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_398),
.A2(n_378),
.B1(n_366),
.B2(n_354),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_398),
.A2(n_394),
.B1(n_365),
.B2(n_388),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_413),
.B(n_356),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_455),
.C(n_413),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_401),
.B(n_315),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_454),
.A2(n_397),
.B(n_427),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_409),
.B(n_346),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_392),
.Y(n_456)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_456),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_428),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_457),
.A2(n_415),
.B1(n_412),
.B2(n_400),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_419),
.A2(n_305),
.B1(n_394),
.B2(n_383),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_359),
.Y(n_462)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_462),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_410),
.Y(n_467)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_467),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_470),
.B(n_477),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_449),
.A2(n_397),
.B1(n_380),
.B2(n_396),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_471),
.A2(n_482),
.B1(n_461),
.B2(n_460),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_443),
.B(n_424),
.C(n_402),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_473),
.B(n_478),
.C(n_481),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_437),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_476),
.B(n_483),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_450),
.B(n_396),
.Y(n_477)
);

MAJx2_ASAP7_75t_L g478 ( 
.A(n_443),
.B(n_403),
.C(n_421),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_479),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_SL g480 ( 
.A(n_437),
.B(n_421),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_480),
.A2(n_494),
.B(n_466),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_425),
.C(n_362),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_463),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_439),
.B(n_404),
.Y(n_484)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_484),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g485 ( 
.A(n_445),
.Y(n_485)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_485),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_456),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_486),
.B(n_489),
.Y(n_507)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_441),
.Y(n_487)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_487),
.Y(n_496)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_438),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_440),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_490),
.A2(n_492),
.B1(n_493),
.B2(n_464),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_452),
.B(n_339),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_491),
.B(n_442),
.Y(n_503)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_441),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_454),
.A2(n_380),
.B(n_400),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_436),
.B(n_324),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_495),
.B(n_434),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_482),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_501),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_499),
.A2(n_493),
.B1(n_451),
.B2(n_465),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_470),
.B(n_436),
.C(n_460),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_503),
.B(n_395),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_439),
.C(n_446),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_504),
.B(n_505),
.Y(n_521)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_467),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_508),
.B(n_513),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_446),
.C(n_454),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_518),
.C(n_494),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_495),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_484),
.Y(n_512)
);

NAND3xp33_ASAP7_75t_SL g524 ( 
.A(n_512),
.B(n_469),
.C(n_475),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_481),
.B(n_433),
.Y(n_513)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_515),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_478),
.B(n_458),
.C(n_459),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_510),
.A2(n_480),
.B(n_474),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_522),
.A2(n_525),
.B(n_529),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_523),
.B(n_536),
.Y(n_542)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_524),
.Y(n_540)
);

A2O1A1O1Ixp25_ASAP7_75t_L g525 ( 
.A1(n_509),
.A2(n_466),
.B(n_472),
.C(n_469),
.D(n_471),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_506),
.B(n_468),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_527),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_516),
.A2(n_468),
.B1(n_472),
.B2(n_492),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_491),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_531),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_501),
.B(n_458),
.C(n_487),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_532),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_497),
.A2(n_395),
.B1(n_420),
.B2(n_438),
.Y(n_533)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_533),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_499),
.A2(n_514),
.B1(n_517),
.B2(n_508),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_534),
.B(n_537),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_535),
.B(n_503),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_514),
.A2(n_438),
.B1(n_465),
.B2(n_387),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_347),
.Y(n_538)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_538),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_511),
.C(n_500),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_541),
.B(n_542),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_513),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_543),
.B(n_545),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_536),
.B(n_511),
.C(n_500),
.Y(n_545)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_546),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_531),
.B(n_502),
.C(n_496),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_542),
.C(n_545),
.Y(n_556)
);

OA21x2_ASAP7_75t_L g551 ( 
.A1(n_534),
.A2(n_502),
.B(n_507),
.Y(n_551)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_551),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_520),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_553),
.A2(n_496),
.B1(n_519),
.B2(n_525),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_538),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g563 ( 
.A1(n_554),
.A2(n_537),
.B1(n_345),
.B2(n_387),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_558),
.Y(n_575)
);

INVx6_ASAP7_75t_L g558 ( 
.A(n_549),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_555),
.A2(n_529),
.B(n_521),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_559),
.A2(n_560),
.B(n_561),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_535),
.C(n_522),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g572 ( 
.A(n_563),
.B(n_551),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_543),
.B(n_359),
.C(n_357),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_565),
.B(n_567),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_540),
.A2(n_304),
.B1(n_357),
.B2(n_301),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_566),
.B(n_544),
.C(n_552),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_569),
.C(n_570),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_550),
.C(n_553),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_562),
.B(n_548),
.C(n_551),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_572),
.A2(n_547),
.B1(n_564),
.B2(n_539),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_547),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_573),
.B(n_565),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_574),
.A2(n_557),
.B(n_555),
.Y(n_577)
);

O2A1O1Ixp33_ASAP7_75t_SL g582 ( 
.A1(n_577),
.A2(n_561),
.B(n_539),
.C(n_567),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_578),
.B(n_579),
.C(n_559),
.Y(n_581)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_575),
.B(n_560),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_SL g583 ( 
.A(n_580),
.B(n_571),
.Y(n_583)
);

AOI322xp5_ASAP7_75t_L g584 ( 
.A1(n_581),
.A2(n_582),
.A3(n_583),
.B1(n_571),
.B2(n_577),
.C1(n_564),
.C2(n_576),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_584),
.A2(n_585),
.B(n_341),
.Y(n_586)
);

AOI322xp5_ASAP7_75t_L g585 ( 
.A1(n_583),
.A2(n_426),
.A3(n_417),
.B1(n_304),
.B2(n_546),
.C1(n_300),
.C2(n_314),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_586),
.A2(n_10),
.B(n_11),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_10),
.C(n_11),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_588),
.A2(n_14),
.B(n_10),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_589),
.B(n_12),
.Y(n_590)
);


endmodule