module real_aes_3474_n_297 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_296, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_297);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_296;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_297;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_792;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_1089;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_856;
wire n_594;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_961;
wire n_870;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_1040;
wire n_415;
wire n_572;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_1078;
wire n_495;
wire n_892;
wire n_994;
wire n_370;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_931;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_973;
wire n_1081;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_999;
wire n_913;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_501;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_303;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_1079;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1003;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_359;
wire n_717;
wire n_982;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_1088;
wire n_1055;
wire n_988;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_1097;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_1076;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_0), .A2(n_29), .B1(n_553), .B2(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_1), .Y(n_308) );
AND2x4_ASAP7_75t_L g850 ( .A(n_1), .B(n_289), .Y(n_850) );
AND2x4_ASAP7_75t_L g855 ( .A(n_1), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g615 ( .A(n_2), .Y(n_615) );
INVx1_ASAP7_75t_L g743 ( .A(n_3), .Y(n_743) );
INVx1_ASAP7_75t_SL g760 ( .A(n_4), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_5), .A2(n_85), .B1(n_556), .B2(n_558), .Y(n_555) );
AO22x1_ASAP7_75t_L g876 ( .A1(n_6), .A2(n_11), .B1(n_851), .B2(n_861), .Y(n_876) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_7), .A2(n_83), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_8), .A2(n_260), .B1(n_372), .B2(n_376), .Y(n_371) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_9), .A2(n_113), .B1(n_452), .B2(n_453), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_10), .A2(n_218), .B1(n_854), .B2(n_857), .Y(n_853) );
XOR2x2_ASAP7_75t_SL g1064 ( .A(n_11), .B(n_1065), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_11), .A2(n_1090), .B1(n_1092), .B2(n_1095), .Y(n_1089) );
INVx1_ASAP7_75t_L g1075 ( .A(n_12), .Y(n_1075) );
INVx1_ASAP7_75t_L g1078 ( .A(n_13), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_14), .A2(n_182), .B1(n_449), .B2(n_450), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_15), .A2(n_62), .B1(n_393), .B2(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_16), .A2(n_148), .B1(n_576), .B2(n_581), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_17), .A2(n_101), .B1(n_667), .B2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_18), .A2(n_270), .B1(n_438), .B2(n_439), .Y(n_437) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_19), .A2(n_408), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g777 ( .A(n_20), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_21), .A2(n_160), .B1(n_655), .B2(n_658), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g831 ( .A1(n_22), .A2(n_244), .B1(n_458), .B2(n_459), .Y(n_831) );
AOI21xp33_ASAP7_75t_SL g348 ( .A1(n_23), .A2(n_349), .B(n_355), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_24), .A2(n_255), .B1(n_435), .B2(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g1074 ( .A(n_25), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_26), .A2(n_34), .B1(n_471), .B2(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g819 ( .A(n_27), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_27), .A2(n_139), .B1(n_874), .B2(n_885), .Y(n_884) );
AO22x1_ASAP7_75t_L g457 ( .A1(n_28), .A2(n_163), .B1(n_458), .B2(n_459), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_30), .A2(n_63), .B1(n_484), .B2(n_553), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_31), .A2(n_175), .B1(n_479), .B2(n_480), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_32), .A2(n_267), .B1(n_539), .B2(n_634), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_33), .A2(n_75), .B1(n_436), .B2(n_438), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_35), .A2(n_112), .B1(n_433), .B2(n_441), .Y(n_597) );
INVx1_ASAP7_75t_L g1081 ( .A(n_36), .Y(n_1081) );
INVx1_ASAP7_75t_L g721 ( .A(n_37), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_38), .A2(n_441), .B(n_442), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_39), .B(n_225), .Y(n_306) );
INVx1_ASAP7_75t_L g345 ( .A(n_39), .Y(n_345) );
INVxp67_ASAP7_75t_L g424 ( .A(n_39), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_40), .A2(n_1065), .B1(n_1093), .B2(n_1094), .Y(n_1092) );
CKINVDCx20_ASAP7_75t_R g1093 ( .A(n_40), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_41), .A2(n_126), .B1(n_629), .B2(n_697), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_42), .A2(n_208), .B1(n_414), .B2(n_416), .Y(n_413) );
AOI21xp33_ASAP7_75t_SL g525 ( .A1(n_43), .A2(n_526), .B(n_527), .Y(n_525) );
INVx1_ASAP7_75t_L g751 ( .A(n_44), .Y(n_751) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_45), .A2(n_79), .B1(n_433), .B2(n_441), .C(n_502), .Y(n_501) );
AO22x1_ASAP7_75t_L g451 ( .A1(n_46), .A2(n_156), .B1(n_452), .B2(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_47), .B(n_562), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_48), .B(n_486), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_49), .A2(n_121), .B1(n_449), .B2(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_50), .B(n_330), .Y(n_341) );
INVx1_ASAP7_75t_L g679 ( .A(n_51), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_52), .A2(n_278), .B1(n_534), .B2(n_536), .Y(n_810) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_53), .A2(n_287), .B1(n_397), .B2(n_543), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_54), .A2(n_136), .B1(n_393), .B2(n_397), .Y(n_392) );
OAI21x1_ASAP7_75t_L g493 ( .A1(n_55), .A2(n_494), .B(n_511), .Y(n_493) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_55), .B(n_495), .C(n_500), .D(n_507), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_56), .A2(n_199), .B1(n_474), .B2(n_476), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_57), .A2(n_205), .B1(n_476), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_58), .A2(n_96), .B1(n_438), .B2(n_439), .Y(n_598) );
INVxp67_ASAP7_75t_R g318 ( .A(n_59), .Y(n_318) );
INVx1_ASAP7_75t_L g427 ( .A(n_59), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_60), .A2(n_226), .B1(n_414), .B2(n_484), .Y(n_626) );
OAI22x1_ASAP7_75t_L g547 ( .A1(n_61), .A2(n_548), .B1(n_584), .B2(n_585), .Y(n_547) );
INVx1_ASAP7_75t_L g585 ( .A(n_61), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g866 ( .A1(n_61), .A2(n_190), .B1(n_847), .B2(n_851), .Y(n_866) );
XOR2x2_ASAP7_75t_L g671 ( .A(n_64), .B(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_65), .A2(n_272), .B1(n_552), .B2(n_554), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_66), .A2(n_168), .B1(n_581), .B2(n_583), .Y(n_580) );
NAND2xp33_ASAP7_75t_L g822 ( .A(n_67), .B(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_68), .A2(n_211), .B1(n_655), .B2(n_697), .Y(n_1067) );
INVx2_ASAP7_75t_L g303 ( .A(n_69), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_70), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g719 ( .A(n_71), .Y(n_719) );
AOI21xp33_ASAP7_75t_L g488 ( .A1(n_72), .A2(n_489), .B(n_490), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_73), .A2(n_234), .B1(n_531), .B2(n_532), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_74), .A2(n_196), .B1(n_576), .B2(n_582), .Y(n_630) );
INVx1_ASAP7_75t_L g849 ( .A(n_76), .Y(n_849) );
AND2x4_ASAP7_75t_L g852 ( .A(n_76), .B(n_303), .Y(n_852) );
INVx1_ASAP7_75t_SL g883 ( .A(n_76), .Y(n_883) );
INVx1_ASAP7_75t_L g782 ( .A(n_77), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_78), .A2(n_232), .B1(n_458), .B2(n_459), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_80), .A2(n_207), .B1(n_861), .B2(n_905), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_81), .B(n_323), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_82), .A2(n_169), .B1(n_393), .B2(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_84), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_86), .A2(n_166), .B1(n_435), .B2(n_436), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_87), .A2(n_206), .B1(n_438), .B2(n_439), .Y(n_506) );
INVx1_ASAP7_75t_L g835 ( .A(n_88), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_89), .A2(n_217), .B1(n_435), .B2(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_90), .A2(n_102), .B1(n_572), .B2(n_573), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_91), .A2(n_129), .B1(n_400), .B2(n_402), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_92), .A2(n_198), .B1(n_435), .B2(n_436), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_93), .A2(n_233), .B1(n_693), .B2(n_793), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_94), .A2(n_141), .B1(n_384), .B2(n_545), .Y(n_691) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_95), .A2(n_280), .B1(n_449), .B2(n_499), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_97), .A2(n_246), .B1(n_509), .B2(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_98), .B(n_436), .Y(n_784) );
INVx1_ASAP7_75t_L g802 ( .A(n_99), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g871 ( .A1(n_100), .A2(n_180), .B1(n_854), .B2(n_872), .Y(n_871) );
OAI22x1_ASAP7_75t_L g789 ( .A1(n_103), .A2(n_790), .B1(n_804), .B2(n_815), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_103), .B(n_791), .C(n_795), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_103), .A2(n_215), .B1(n_847), .B2(n_851), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_104), .A2(n_192), .B1(n_851), .B2(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_105), .A2(n_241), .B1(n_509), .B2(n_629), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_106), .A2(n_675), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g331 ( .A(n_107), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_107), .B(n_224), .Y(n_421) );
INVx1_ASAP7_75t_L g503 ( .A(n_108), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_109), .A2(n_115), .B1(n_400), .B2(n_402), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_110), .A2(n_247), .B1(n_384), .B2(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g491 ( .A(n_111), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_114), .A2(n_171), .B1(n_393), .B2(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_116), .A2(n_186), .B1(n_854), .B2(n_902), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_117), .A2(n_273), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_118), .A2(n_128), .B1(n_854), .B2(n_857), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_119), .A2(n_214), .B1(n_376), .B2(n_634), .Y(n_1069) );
INVx1_ASAP7_75t_L g443 ( .A(n_120), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_122), .B(n_661), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_123), .A2(n_203), .B1(n_455), .B2(n_456), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_124), .A2(n_200), .B1(n_376), .B2(n_634), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_125), .A2(n_285), .B1(n_449), .B2(n_452), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_127), .A2(n_251), .B1(n_379), .B2(n_384), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_130), .A2(n_132), .B1(n_379), .B2(n_384), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_131), .A2(n_235), .B1(n_482), .B2(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g623 ( .A(n_133), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_134), .B(n_682), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_135), .A2(n_145), .B1(n_902), .B2(n_931), .Y(n_930) );
AO22x2_ASAP7_75t_L g734 ( .A1(n_137), .A2(n_735), .B1(n_740), .B2(n_757), .Y(n_734) );
INVxp33_ASAP7_75t_SL g756 ( .A(n_137), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_138), .A2(n_219), .B1(n_400), .B2(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_140), .A2(n_201), .B1(n_476), .B2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_142), .A2(n_173), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_143), .A2(n_279), .B1(n_854), .B2(n_857), .Y(n_867) );
INVx1_ASAP7_75t_L g749 ( .A(n_144), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_146), .A2(n_154), .B1(n_372), .B2(n_539), .Y(n_538) );
AO22x1_ASAP7_75t_L g454 ( .A1(n_147), .A2(n_284), .B1(n_455), .B2(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g1079 ( .A(n_149), .Y(n_1079) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_150), .A2(n_236), .B1(n_450), .B2(n_456), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_151), .A2(n_256), .B1(n_453), .B2(n_455), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_152), .A2(n_204), .B1(n_452), .B2(n_453), .Y(n_829) );
INVx1_ASAP7_75t_L g753 ( .A(n_153), .Y(n_753) );
INVx1_ASAP7_75t_L g779 ( .A(n_155), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_157), .A2(n_164), .B1(n_534), .B2(n_536), .Y(n_533) );
INVx1_ASAP7_75t_L g669 ( .A(n_158), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_159), .A2(n_239), .B1(n_452), .B2(n_453), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_161), .A2(n_183), .B1(n_543), .B2(n_700), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_162), .A2(n_176), .B1(n_582), .B2(n_629), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g881 ( .A1(n_165), .A2(n_276), .B1(n_857), .B2(n_882), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_167), .A2(n_189), .B1(n_449), .B2(n_450), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_170), .B(n_524), .Y(n_523) );
CKINVDCx14_ASAP7_75t_R g593 ( .A(n_172), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_174), .A2(n_238), .B1(n_807), .B2(n_809), .Y(n_806) );
AOI22xp5_ASAP7_75t_L g692 ( .A1(n_177), .A2(n_253), .B1(n_372), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_178), .A2(n_188), .B1(n_372), .B2(n_376), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_179), .A2(n_228), .B1(n_400), .B2(n_700), .Y(n_710) );
XNOR2x2_ASAP7_75t_L g429 ( .A(n_181), .B(n_430), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g873 ( .A1(n_184), .A2(n_240), .B1(n_847), .B2(n_874), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_185), .B(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_187), .A2(n_216), .B1(n_543), .B2(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g775 ( .A(n_191), .Y(n_775) );
AO221x2_ASAP7_75t_L g875 ( .A1(n_193), .A2(n_250), .B1(n_854), .B2(n_872), .C(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_194), .A2(n_258), .B1(n_480), .B2(n_668), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_195), .A2(n_265), .B1(n_452), .B2(n_453), .Y(n_768) );
OA22x2_ASAP7_75t_L g335 ( .A1(n_197), .A2(n_225), .B1(n_330), .B2(n_334), .Y(n_335) );
INVx1_ASAP7_75t_L g368 ( .A(n_197), .Y(n_368) );
AOI21xp5_ASAP7_75t_SL g773 ( .A1(n_202), .A2(n_441), .B(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_209), .A2(n_227), .B1(n_414), .B2(n_661), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_210), .A2(n_229), .B1(n_458), .B2(n_459), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_212), .A2(n_277), .B1(n_576), .B2(n_578), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_213), .A2(n_282), .B1(n_847), .B2(n_905), .Y(n_904) );
INVx1_ASAP7_75t_L g528 ( .A(n_220), .Y(n_528) );
INVx1_ASAP7_75t_L g746 ( .A(n_221), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_222), .A2(n_252), .B1(n_384), .B2(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_223), .A2(n_796), .B(n_799), .Y(n_795) );
INVx1_ASAP7_75t_L g347 ( .A(n_224), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_224), .B(n_365), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g387 ( .A1(n_225), .A2(n_248), .B(n_388), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g765 ( .A1(n_230), .A2(n_266), .B1(n_449), .B2(n_450), .Y(n_765) );
INVx1_ASAP7_75t_L g771 ( .A(n_231), .Y(n_771) );
INVx1_ASAP7_75t_L g724 ( .A(n_237), .Y(n_724) );
INVx1_ASAP7_75t_L g520 ( .A(n_240), .Y(n_520) );
INVx1_ASAP7_75t_L g716 ( .A(n_242), .Y(n_716) );
INVx1_ASAP7_75t_L g800 ( .A(n_243), .Y(n_800) );
INVx1_ASAP7_75t_SL g727 ( .A(n_245), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_248), .B(n_281), .Y(n_307) );
INVx1_ASAP7_75t_L g333 ( .A(n_248), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_249), .A2(n_292), .B1(n_455), .B2(n_456), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_254), .A2(n_291), .B1(n_560), .B2(n_561), .C(n_563), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_257), .A2(n_264), .B1(n_697), .B2(n_814), .Y(n_813) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_259), .Y(n_356) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_261), .A2(n_269), .B1(n_480), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g464 ( .A(n_262), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_263), .A2(n_283), .B1(n_400), .B2(n_658), .Y(n_657) );
AOI21xp33_ASAP7_75t_SL g833 ( .A1(n_268), .A2(n_441), .B(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_271), .A2(n_294), .B1(n_408), .B2(n_410), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_274), .A2(n_296), .B1(n_699), .B2(n_700), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_275), .A2(n_687), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_281), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_286), .B(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_288), .A2(n_290), .B1(n_400), .B2(n_707), .Y(n_738) );
INVx1_ASAP7_75t_L g856 ( .A(n_289), .Y(n_856) );
INVx1_ASAP7_75t_L g564 ( .A(n_293), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_295), .B(n_323), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_309), .B(n_839), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
BUFx4_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
NAND3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_304), .C(n_308), .Y(n_300) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_301), .B(n_1087), .Y(n_1086) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_301), .B(n_1088), .Y(n_1091) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OA21x2_ASAP7_75t_L g1096 ( .A1(n_302), .A2(n_883), .B(n_1097), .Y(n_1096) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g848 ( .A(n_303), .B(n_849), .Y(n_848) );
AND3x4_ASAP7_75t_L g882 ( .A(n_303), .B(n_855), .C(n_883), .Y(n_882) );
NOR2xp33_ASAP7_75t_L g1087 ( .A(n_304), .B(n_1088), .Y(n_1087) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AO21x2_ASAP7_75t_L g360 ( .A1(n_305), .A2(n_361), .B(n_363), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g1088 ( .A(n_308), .Y(n_1088) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_644), .Y(n_309) );
XNOR2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_514), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_460), .B2(n_513), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OA22x2_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_317), .B1(n_428), .B2(n_429), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B(n_425), .Y(n_317) );
NOR4xp75_ASAP7_75t_L g319 ( .A(n_320), .B(n_369), .C(n_390), .D(n_405), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND4xp75_ASAP7_75t_L g425 ( .A(n_321), .B(n_370), .C(n_391), .D(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_348), .Y(n_321) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g524 ( .A(n_324), .Y(n_524) );
INVx1_ASAP7_75t_L g562 ( .A(n_324), .Y(n_562) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g677 ( .A(n_325), .Y(n_677) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g487 ( .A(n_326), .Y(n_487) );
BUFx3_ASAP7_75t_L g667 ( .A(n_326), .Y(n_667) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_336), .Y(n_326) );
AND2x4_ASAP7_75t_L g380 ( .A(n_327), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g401 ( .A(n_327), .B(n_395), .Y(n_401) );
AND2x2_ASAP7_75t_L g415 ( .A(n_327), .B(n_354), .Y(n_415) );
AND2x2_ASAP7_75t_L g433 ( .A(n_327), .B(n_336), .Y(n_433) );
AND2x4_ASAP7_75t_L g435 ( .A(n_327), .B(n_354), .Y(n_435) );
AND2x4_ASAP7_75t_L g449 ( .A(n_327), .B(n_389), .Y(n_449) );
AND2x4_ASAP7_75t_L g452 ( .A(n_327), .B(n_395), .Y(n_452) );
AND2x2_ASAP7_75t_L g577 ( .A(n_327), .B(n_395), .Y(n_577) );
AND2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_335), .Y(n_327) );
INVx1_ASAP7_75t_L g353 ( .A(n_328), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
NAND2xp33_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g334 ( .A(n_330), .Y(n_334) );
INVx3_ASAP7_75t_L g340 ( .A(n_330), .Y(n_340) );
NAND2xp33_ASAP7_75t_L g346 ( .A(n_330), .B(n_347), .Y(n_346) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
INVx1_ASAP7_75t_L g388 ( .A(n_330), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_331), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_333), .A2(n_388), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g352 ( .A(n_335), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
AND2x2_ASAP7_75t_L g422 ( .A(n_335), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g377 ( .A(n_336), .B(n_374), .Y(n_377) );
AND2x4_ASAP7_75t_L g409 ( .A(n_336), .B(n_352), .Y(n_409) );
AND2x4_ASAP7_75t_L g412 ( .A(n_336), .B(n_386), .Y(n_412) );
AND2x4_ASAP7_75t_L g439 ( .A(n_336), .B(n_386), .Y(n_439) );
AND2x2_ASAP7_75t_L g441 ( .A(n_336), .B(n_352), .Y(n_441) );
AND2x4_ASAP7_75t_L g459 ( .A(n_336), .B(n_374), .Y(n_459) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_342), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g354 ( .A(n_338), .B(n_342), .Y(n_354) );
OR2x2_ASAP7_75t_L g382 ( .A(n_338), .B(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g395 ( .A(n_338), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g419 ( .A(n_338), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .Y(n_344) );
INVxp67_ASAP7_75t_L g365 ( .A(n_340), .Y(n_365) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_341), .B(n_364), .C(n_366), .Y(n_363) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g383 ( .A(n_343), .Y(n_383) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g526 ( .A(n_350), .Y(n_526) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g479 ( .A(n_351), .Y(n_479) );
BUFx3_ASAP7_75t_L g553 ( .A(n_351), .Y(n_553) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_351), .Y(n_687) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
AND2x4_ASAP7_75t_L g438 ( .A(n_352), .B(n_354), .Y(n_438) );
AND2x4_ASAP7_75t_L g374 ( .A(n_353), .B(n_375), .Y(n_374) );
AND2x4_ASAP7_75t_L g373 ( .A(n_354), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g458 ( .A(n_354), .B(n_374), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_357), .B(n_528), .Y(n_527) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_SL g601 ( .A(n_359), .Y(n_601) );
BUFx6f_ASAP7_75t_L g624 ( .A(n_359), .Y(n_624) );
INVx1_ASAP7_75t_L g682 ( .A(n_359), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_359), .B(n_775), .Y(n_774) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx3_ASAP7_75t_L g445 ( .A(n_360), .Y(n_445) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_362), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_365), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g386 ( .A(n_366), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_378), .Y(n_370) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx3_ASAP7_75t_L g475 ( .A(n_373), .Y(n_475) );
BUFx12f_ASAP7_75t_L g634 ( .A(n_373), .Y(n_634) );
AND2x4_ASAP7_75t_L g394 ( .A(n_374), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g398 ( .A(n_374), .B(n_389), .Y(n_398) );
AND2x4_ASAP7_75t_L g455 ( .A(n_374), .B(n_395), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_374), .B(n_381), .Y(n_456) );
BUFx2_ASAP7_75t_SL g573 ( .A(n_376), .Y(n_573) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g476 ( .A(n_377), .Y(n_476) );
BUFx5_ASAP7_75t_L g539 ( .A(n_377), .Y(n_539) );
INVx1_ASAP7_75t_L g695 ( .A(n_377), .Y(n_695) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_380), .Y(n_545) );
BUFx12f_ASAP7_75t_L g582 ( .A(n_380), .Y(n_582) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_380), .Y(n_707) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g389 ( .A(n_382), .Y(n_389) );
INVx1_ASAP7_75t_L g396 ( .A(n_383), .Y(n_396) );
BUFx3_ASAP7_75t_L g583 ( .A(n_384), .Y(n_583) );
BUFx12f_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx6_ASAP7_75t_L g469 ( .A(n_385), .Y(n_469) );
AND2x4_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
AND2x4_ASAP7_75t_L g404 ( .A(n_386), .B(n_395), .Y(n_404) );
AND2x4_ASAP7_75t_L g450 ( .A(n_386), .B(n_389), .Y(n_450) );
AND2x4_ASAP7_75t_L g453 ( .A(n_386), .B(n_395), .Y(n_453) );
INVx2_ASAP7_75t_SL g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_399), .Y(n_391) );
BUFx6f_ASAP7_75t_L g568 ( .A(n_393), .Y(n_568) );
BUFx12f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_394), .Y(n_543) );
BUFx6f_ASAP7_75t_L g655 ( .A(n_394), .Y(n_655) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_398), .Y(n_471) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_398), .Y(n_509) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_398), .Y(n_697) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx8_ASAP7_75t_L g699 ( .A(n_401), .Y(n_699) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g579 ( .A(n_403), .Y(n_579) );
INVx1_ASAP7_75t_L g632 ( .A(n_403), .Y(n_632) );
INVx4_ASAP7_75t_L g658 ( .A(n_403), .Y(n_658) );
INVx4_ASAP7_75t_L g700 ( .A(n_403), .Y(n_700) );
INVx4_ASAP7_75t_L g1071 ( .A(n_403), .Y(n_1071) );
INVx8_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g426 ( .A(n_406), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_413), .Y(n_406) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_409), .Y(n_489) );
INVx2_ASAP7_75t_L g535 ( .A(n_409), .Y(n_535) );
INVx2_ASAP7_75t_L g665 ( .A(n_409), .Y(n_665) );
BUFx3_ASAP7_75t_L g745 ( .A(n_409), .Y(n_745) );
INVx3_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g558 ( .A(n_411), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_411), .A2(n_744), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
INVx3_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_412), .Y(n_484) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_412), .Y(n_536) );
BUFx3_ASAP7_75t_L g554 ( .A(n_414), .Y(n_554) );
INVx3_ASAP7_75t_L g725 ( .A(n_414), .Y(n_725) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g483 ( .A(n_415), .Y(n_483) );
BUFx3_ASAP7_75t_L g531 ( .A(n_415), .Y(n_531) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g532 ( .A(n_417), .Y(n_532) );
INVx3_ASAP7_75t_L g560 ( .A(n_417), .Y(n_560) );
INVx4_ASAP7_75t_L g661 ( .A(n_417), .Y(n_661) );
INVx5_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
BUFx4f_ASAP7_75t_L g480 ( .A(n_418), .Y(n_480) );
BUFx2_ASAP7_75t_L g620 ( .A(n_418), .Y(n_620) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_422), .Y(n_418) );
AND2x4_ASAP7_75t_L g436 ( .A(n_419), .B(n_422), .Y(n_436) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_446), .Y(n_430) );
AND4x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .C(n_437), .D(n_440), .Y(n_431) );
INVx2_ASAP7_75t_L g772 ( .A(n_433), .Y(n_772) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_433), .Y(n_823) );
INVx1_ASAP7_75t_L g783 ( .A(n_435), .Y(n_783) );
INVx2_ASAP7_75t_L g778 ( .A(n_438), .Y(n_778) );
INVx2_ASAP7_75t_L g780 ( .A(n_439), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx4_ASAP7_75t_L g668 ( .A(n_444), .Y(n_668) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g492 ( .A(n_445), .Y(n_492) );
NOR4xp25_ASAP7_75t_L g446 ( .A(n_447), .B(n_451), .C(n_454), .D(n_457), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_461), .Y(n_513) );
AO22x2_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_463), .B1(n_493), .B2(n_512), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
XNOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_466), .B(n_477), .Y(n_465) );
NAND4xp25_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .C(n_472), .D(n_473), .Y(n_466) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_L g499 ( .A(n_469), .Y(n_499) );
INVx5_ASAP7_75t_L g629 ( .A(n_469), .Y(n_629) );
INVx1_ASAP7_75t_L g814 ( .A(n_469), .Y(n_814) );
INVx1_ASAP7_75t_L g570 ( .A(n_471), .Y(n_570) );
BUFx4f_ASAP7_75t_L g793 ( .A(n_474), .Y(n_793) );
INVx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g497 ( .A(n_475), .Y(n_497) );
INVx1_ASAP7_75t_L g572 ( .A(n_475), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_481), .C(n_485), .D(n_488), .Y(n_477) );
INVx2_ASAP7_75t_L g808 ( .A(n_479), .Y(n_808) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g689 ( .A(n_483), .Y(n_689) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g798 ( .A(n_487), .Y(n_798) );
INVx2_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_492), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_492), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g512 ( .A(n_493), .Y(n_512) );
AND3x1_ASAP7_75t_L g494 ( .A(n_495), .B(n_500), .C(n_507), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_504), .Y(n_500) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_510), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_589), .B1(n_642), .B2(n_643), .Y(n_514) );
INVx1_ASAP7_75t_L g642 ( .A(n_515), .Y(n_642) );
AO22x2_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_546), .B1(n_586), .B2(n_587), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_SL g588 ( .A(n_519), .Y(n_588) );
XNOR2x1_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
NOR4xp75_ASAP7_75t_L g521 ( .A(n_522), .B(n_529), .C(n_537), .D(n_541), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_525), .Y(n_522) );
INVx2_ASAP7_75t_L g750 ( .A(n_526), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_533), .Y(n_529) );
INVx2_ASAP7_75t_L g1076 ( .A(n_531), .Y(n_1076) );
INVx2_ASAP7_75t_L g720 ( .A(n_534), .Y(n_720) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
BUFx3_ASAP7_75t_L g685 ( .A(n_536), .Y(n_685) );
INVx4_ASAP7_75t_L g722 ( .A(n_536), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_538), .B(n_540), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_542), .B(n_544), .Y(n_541) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g586 ( .A(n_547), .Y(n_586) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_565), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_549), .B(n_565), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_559), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g747 ( .A(n_558), .Y(n_747) );
INVx1_ASAP7_75t_L g801 ( .A(n_560), .Y(n_801) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_566), .B(n_574), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_571), .Y(n_566) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_580), .Y(n_574) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
BUFx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g643 ( .A(n_589), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_610), .B2(n_641), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI21x1_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_607), .Y(n_592) );
NAND3xp33_ASAP7_75t_SL g607 ( .A(n_593), .B(n_608), .C(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_602), .Y(n_595) );
INVx1_ASAP7_75t_L g609 ( .A(n_596), .Y(n_609) );
NAND4xp25_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .C(n_599), .D(n_600), .Y(n_596) );
INVxp67_ASAP7_75t_L g608 ( .A(n_602), .Y(n_608) );
NAND4xp25_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .C(n_605), .D(n_606), .Y(n_602) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g641 ( .A(n_611), .Y(n_641) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI21x1_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_616), .B(n_635), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_614), .B(n_626), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_615), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g616 ( .A(n_617), .B(n_627), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g617 ( .A(n_618), .B(n_625), .C(n_626), .Y(n_617) );
INVx1_ASAP7_75t_L g639 ( .A(n_618), .Y(n_639) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_621), .Y(n_618) );
INVxp67_ASAP7_75t_L g680 ( .A(n_620), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g755 ( .A(n_624), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_624), .B(n_835), .Y(n_834) );
INVxp67_ASAP7_75t_L g637 ( .A(n_625), .Y(n_637) );
INVx1_ASAP7_75t_L g640 ( .A(n_627), .Y(n_640) );
NAND4xp25_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .C(n_631), .D(n_633), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_640), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .C(n_639), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_730), .B1(n_837), .B2(n_838), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
HB1xp67_ASAP7_75t_L g837 ( .A(n_646), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_701), .B1(n_728), .B2(n_729), .Y(n_646) );
INVx1_ASAP7_75t_L g728 ( .A(n_647), .Y(n_728) );
AO22x2_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_649), .B1(n_670), .B2(n_671), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_669), .Y(n_650) );
NOR2x1_ASAP7_75t_L g651 ( .A(n_652), .B(n_659), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .C(n_656), .D(n_657), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_662), .C(n_663), .D(n_666), .Y(n_659) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g684 ( .A(n_665), .Y(n_684) );
INVx2_ASAP7_75t_L g803 ( .A(n_668), .Y(n_803) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NOR2x1_ASAP7_75t_L g672 ( .A(n_673), .B(n_690), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_683), .C(n_686), .Y(n_673) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_676), .A2(n_753), .B(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g717 ( .A(n_682), .Y(n_717) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g809 ( .A(n_689), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g690 ( .A(n_691), .B(n_692), .C(n_696), .D(n_698), .Y(n_690) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g729 ( .A(n_703), .Y(n_729) );
XOR2x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_727), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_705), .B(n_711), .Y(n_704) );
AND4x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .C(n_709), .D(n_710), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_712), .B(n_718), .C(n_723), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_721), .B2(n_722), .Y(n_718) );
OAI21xp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_725), .B(n_726), .Y(n_723) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_725), .A2(n_749), .B1(n_750), .B2(n_751), .Y(n_748) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g838 ( .A(n_731), .Y(n_838) );
OAI22x1_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B1(n_787), .B2(n_788), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AO22x2_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_758), .B1(n_785), .B2(n_786), .Y(n_733) );
INVx2_ASAP7_75t_L g786 ( .A(n_734), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_735), .B(n_741), .Y(n_757) );
AND4x1_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .C(n_738), .D(n_739), .Y(n_735) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_756), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g741 ( .A(n_742), .B(n_748), .C(n_752), .Y(n_741) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_746), .B2(n_747), .Y(n_742) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_750), .A2(n_1074), .B1(n_1075), .B2(n_1076), .Y(n_1073) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
XNOR2x1_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
XNOR2xp5_ASAP7_75t_L g785 ( .A(n_760), .B(n_761), .Y(n_785) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_769), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_768), .Y(n_766) );
NOR3xp33_ASAP7_75t_L g769 ( .A(n_770), .B(n_776), .C(n_781), .Y(n_769) );
OAI21xp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_772), .B(n_773), .Y(n_770) );
OAI22xp33_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_776) );
INVxp67_ASAP7_75t_L g825 ( .A(n_780), .Y(n_825) );
OAI21xp5_ASAP7_75t_SL g781 ( .A1(n_782), .A2(n_783), .B(n_784), .Y(n_781) );
INVx2_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
OA22x2_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_816), .B1(n_817), .B2(n_836), .Y(n_788) );
INVx2_ASAP7_75t_L g836 ( .A(n_789), .Y(n_836) );
AND4x1_ASAP7_75t_L g815 ( .A(n_791), .B(n_795), .C(n_805), .D(n_811), .Y(n_815) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_794), .Y(n_791) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1082 ( .A(n_798), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_811), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_810), .Y(n_805) );
INVx2_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
INVx2_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
INVx3_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
XNOR2x1_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NOR2x1_ASAP7_75t_L g820 ( .A(n_821), .B(n_827), .Y(n_820) );
NAND3xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .C(n_826), .Y(n_821) );
NAND4xp25_ASAP7_75t_SL g827 ( .A(n_828), .B(n_829), .C(n_830), .D(n_833), .Y(n_827) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_832), .Y(n_830) );
OAI221xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_1060), .B1(n_1062), .B2(n_1084), .C(n_1089), .Y(n_839) );
NOR3xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_1018), .C(n_1042), .Y(n_840) );
AOI33xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_906), .A3(n_934), .B1(n_971), .B2(n_996), .B3(n_1009), .Y(n_841) );
A2O1A1Ixp33_ASAP7_75t_SL g842 ( .A1(n_843), .A2(n_863), .B(n_877), .C(n_899), .Y(n_842) );
AND2x2_ASAP7_75t_L g952 ( .A(n_843), .B(n_898), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_843), .B(n_897), .Y(n_1059) );
INVx1_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_844), .A2(n_886), .B1(n_919), .B2(n_924), .C(n_928), .Y(n_918) );
NOR2xp33_ASAP7_75t_L g989 ( .A(n_844), .B(n_942), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_844), .B(n_1005), .Y(n_1004) );
OR2x2_ASAP7_75t_L g844 ( .A(n_845), .B(n_858), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_845), .B(n_864), .Y(n_891) );
INVx4_ASAP7_75t_L g914 ( .A(n_845), .Y(n_914) );
OR2x2_ASAP7_75t_L g917 ( .A(n_845), .B(n_859), .Y(n_917) );
AND2x2_ASAP7_75t_L g959 ( .A(n_845), .B(n_858), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_845), .B(n_864), .Y(n_986) );
NOR2xp33_ASAP7_75t_L g1051 ( .A(n_845), .B(n_865), .Y(n_1051) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_853), .Y(n_845) );
AND2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
AND2x4_ASAP7_75t_L g854 ( .A(n_848), .B(n_855), .Y(n_854) );
AND2x4_ASAP7_75t_L g861 ( .A(n_848), .B(n_850), .Y(n_861) );
AND2x2_ASAP7_75t_L g885 ( .A(n_848), .B(n_850), .Y(n_885) );
AND2x2_ASAP7_75t_L g851 ( .A(n_850), .B(n_852), .Y(n_851) );
AND2x2_ASAP7_75t_L g874 ( .A(n_850), .B(n_852), .Y(n_874) );
AND2x4_ASAP7_75t_L g905 ( .A(n_850), .B(n_852), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g1097 ( .A(n_850), .Y(n_1097) );
AND2x4_ASAP7_75t_L g857 ( .A(n_852), .B(n_855), .Y(n_857) );
AND2x4_ASAP7_75t_L g872 ( .A(n_852), .B(n_855), .Y(n_872) );
INVx3_ASAP7_75t_L g932 ( .A(n_854), .Y(n_932) );
INVx2_ASAP7_75t_SL g903 ( .A(n_857), .Y(n_903) );
INVx2_ASAP7_75t_L g886 ( .A(n_858), .Y(n_886) );
OR2x2_ASAP7_75t_L g950 ( .A(n_858), .B(n_914), .Y(n_950) );
INVxp67_ASAP7_75t_L g981 ( .A(n_858), .Y(n_981) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_858), .B(n_974), .Y(n_1034) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_859), .B(n_900), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_860), .B(n_862), .Y(n_859) );
AND2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_868), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_864), .B(n_869), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_864), .B(n_956), .Y(n_955) );
A2O1A1Ixp33_ASAP7_75t_L g966 ( .A1(n_864), .A2(n_888), .B(n_967), .C(n_969), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_864), .B(n_912), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_864), .B(n_915), .Y(n_1040) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx3_ASAP7_75t_L g898 ( .A(n_865), .Y(n_898) );
INVx2_ASAP7_75t_L g922 ( .A(n_865), .Y(n_922) );
AND2x2_ASAP7_75t_L g927 ( .A(n_865), .B(n_869), .Y(n_927) );
NOR2xp33_ASAP7_75t_L g979 ( .A(n_865), .B(n_961), .Y(n_979) );
AOI321xp33_ASAP7_75t_L g1009 ( .A1(n_865), .A2(n_886), .A3(n_893), .B1(n_1010), .B2(n_1013), .C(n_1014), .Y(n_1009) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_875), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_869), .B(n_889), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_869), .B(n_945), .Y(n_944) );
AND2x2_ASAP7_75t_L g992 ( .A(n_869), .B(n_894), .Y(n_992) );
AND2x2_ASAP7_75t_L g999 ( .A(n_869), .B(n_926), .Y(n_999) );
AND2x2_ASAP7_75t_L g1012 ( .A(n_869), .B(n_879), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_869), .B(n_907), .Y(n_1026) );
A2O1A1Ixp33_ASAP7_75t_SL g1035 ( .A1(n_869), .A2(n_1036), .B(n_1040), .C(n_1041), .Y(n_1035) );
CKINVDCx6p67_ASAP7_75t_R g869 ( .A(n_870), .Y(n_869) );
AND2x2_ASAP7_75t_L g888 ( .A(n_870), .B(n_889), .Y(n_888) );
AND2x2_ASAP7_75t_L g896 ( .A(n_870), .B(n_897), .Y(n_896) );
AND2x2_ASAP7_75t_L g915 ( .A(n_870), .B(n_894), .Y(n_915) );
AND2x2_ASAP7_75t_L g935 ( .A(n_870), .B(n_936), .Y(n_935) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_870), .B(n_889), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g961 ( .A(n_870), .B(n_875), .Y(n_961) );
AND2x2_ASAP7_75t_L g963 ( .A(n_870), .B(n_879), .Y(n_963) );
AND2x2_ASAP7_75t_L g976 ( .A(n_870), .B(n_945), .Y(n_976) );
AND2x2_ASAP7_75t_L g987 ( .A(n_870), .B(n_926), .Y(n_987) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_870), .B(n_880), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_870), .B(n_946), .Y(n_1029) );
AND2x2_ASAP7_75t_L g870 ( .A(n_871), .B(n_873), .Y(n_870) );
AND2x2_ASAP7_75t_L g879 ( .A(n_875), .B(n_880), .Y(n_879) );
OR2x2_ASAP7_75t_L g895 ( .A(n_875), .B(n_880), .Y(n_895) );
AND2x2_ASAP7_75t_L g926 ( .A(n_875), .B(n_889), .Y(n_926) );
INVx1_ASAP7_75t_L g946 ( .A(n_875), .Y(n_946) );
OAI321xp33_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .A3(n_886), .B1(n_887), .B2(n_890), .C(n_892), .Y(n_877) );
AND2x2_ASAP7_75t_L g936 ( .A(n_879), .B(n_898), .Y(n_936) );
INVx1_ASAP7_75t_L g993 ( .A(n_879), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_879), .B(n_896), .Y(n_1058) );
INVx1_ASAP7_75t_L g889 ( .A(n_880), .Y(n_889) );
AND2x2_ASAP7_75t_L g945 ( .A(n_880), .B(n_946), .Y(n_945) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_884), .Y(n_880) );
INVx3_ASAP7_75t_SL g958 ( .A(n_886), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_886), .B(n_974), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g1014 ( .A(n_886), .B(n_1015), .Y(n_1014) );
AOI221xp5_ASAP7_75t_L g1027 ( .A1(n_886), .A2(n_1013), .B1(n_1028), .B2(n_1030), .C(n_1032), .Y(n_1027) );
NAND2xp5_ASAP7_75t_SL g1010 ( .A(n_887), .B(n_1011), .Y(n_1010) );
INVx1_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g951 ( .A(n_888), .B(n_952), .Y(n_951) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_888), .A2(n_928), .B1(n_979), .B2(n_980), .C(n_982), .Y(n_978) );
INVxp67_ASAP7_75t_SL g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_893), .B(n_937), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_893), .B(n_1047), .Y(n_1046) );
AND2x2_ASAP7_75t_L g893 ( .A(n_894), .B(n_896), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
NOR2x1_ASAP7_75t_L g907 ( .A(n_895), .B(n_897), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_897), .B(n_945), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_897), .B(n_983), .Y(n_982) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_897), .B(n_943), .Y(n_1044) );
INVx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g998 ( .A(n_898), .B(n_999), .Y(n_998) );
OAI221xp5_ASAP7_75t_L g953 ( .A1(n_899), .A2(n_954), .B1(n_962), .B2(n_964), .C(n_966), .Y(n_953) );
OAI211xp5_ASAP7_75t_L g1018 ( .A1(n_899), .A2(n_1019), .B(n_1027), .C(n_1035), .Y(n_1018) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
AND2x2_ASAP7_75t_L g948 ( .A(n_900), .B(n_949), .Y(n_948) );
AND2x2_ASAP7_75t_L g965 ( .A(n_900), .B(n_920), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_900), .B(n_938), .Y(n_970) );
INVx4_ASAP7_75t_L g974 ( .A(n_900), .Y(n_974) );
NOR2xp33_ASAP7_75t_L g1008 ( .A(n_900), .B(n_950), .Y(n_1008) );
AND2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_904), .Y(n_900) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
BUFx2_ASAP7_75t_L g1061 ( .A(n_905), .Y(n_1061) );
AOI221xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_908), .B1(n_915), .B2(n_916), .C(n_918), .Y(n_906) );
HB1xp67_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_910), .Y(n_909) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_910), .Y(n_1025) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_912), .Y(n_1047) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
INVx1_ASAP7_75t_L g938 ( .A(n_913), .Y(n_938) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx2_ASAP7_75t_L g920 ( .A(n_914), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_915), .B(n_948), .Y(n_1001) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g995 ( .A(n_917), .B(n_922), .Y(n_995) );
NOR2xp33_ASAP7_75t_L g1041 ( .A(n_917), .B(n_974), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_922), .B(n_941), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_922), .B(n_976), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_922), .B(n_1016), .Y(n_1023) );
INVx1_ASAP7_75t_L g941 ( .A(n_923), .Y(n_941) );
INVxp67_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g1039 ( .A(n_926), .Y(n_1039) );
NOR2xp33_ASAP7_75t_L g988 ( .A(n_928), .B(n_974), .Y(n_988) );
CKINVDCx5p33_ASAP7_75t_R g928 ( .A(n_929), .Y(n_928) );
AND2x2_ASAP7_75t_L g929 ( .A(n_930), .B(n_933), .Y(n_929) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
AOI211xp5_ASAP7_75t_L g934 ( .A1(n_935), .A2(n_937), .B(n_939), .C(n_953), .Y(n_934) );
INVx1_ASAP7_75t_L g1003 ( .A(n_936), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1028 ( .A(n_937), .B(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_942), .B(n_947), .C(n_951), .Y(n_939) );
INVx1_ASAP7_75t_L g1006 ( .A(n_941), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_942), .A2(n_1055), .B1(n_1058), .B2(n_1059), .Y(n_1054) );
INVx2_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g1038 ( .A(n_945), .Y(n_1038) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
O2A1O1Ixp33_ASAP7_75t_L g1048 ( .A1(n_952), .A2(n_1049), .B(n_1052), .C(n_1054), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_958), .B1(n_959), .B2(n_960), .Y(n_954) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx1_ASAP7_75t_L g983 ( .A(n_959), .Y(n_983) );
O2A1O1Ixp33_ASAP7_75t_SL g1019 ( .A1(n_959), .A2(n_992), .B(n_1020), .C(n_1024), .Y(n_1019) );
INVxp67_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
AOI21xp33_ASAP7_75t_L g1032 ( .A1(n_962), .A2(n_1015), .B(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g967 ( .A(n_968), .Y(n_967) );
AOI211xp5_ASAP7_75t_L g996 ( .A1(n_969), .A2(n_997), .B(n_1000), .C(n_1002), .Y(n_996) );
INVx1_ASAP7_75t_L g969 ( .A(n_970), .Y(n_969) );
NOR4xp25_ASAP7_75t_L g971 ( .A(n_972), .B(n_977), .C(n_989), .D(n_990), .Y(n_971) );
NOR2xp33_ASAP7_75t_L g972 ( .A(n_973), .B(n_975), .Y(n_972) );
INVx1_ASAP7_75t_L g1013 ( .A(n_973), .Y(n_1013) );
INVx2_ASAP7_75t_L g1005 ( .A(n_974), .Y(n_1005) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_974), .B(n_981), .Y(n_1045) );
NOR2xp33_ASAP7_75t_L g1053 ( .A(n_976), .B(n_992), .Y(n_1053) );
AOI21xp33_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_984), .B(n_988), .Y(n_977) );
NOR2xp33_ASAP7_75t_L g1021 ( .A(n_979), .B(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_985), .B(n_987), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
AOI21xp33_ASAP7_75t_L g990 ( .A1(n_991), .A2(n_993), .B(n_994), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVxp67_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVxp67_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1004), .B1(n_1006), .B2(n_1007), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1042 ( .A1(n_1005), .A2(n_1043), .B1(n_1045), .B2(n_1046), .C(n_1048), .Y(n_1042) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_1005), .B(n_1050), .Y(n_1049) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .Y(n_1015) );
INVxp67_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
NOR2xp33_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1026), .Y(n_1024) );
INVxp67_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1039), .Y(n_1037) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1047), .B(n_1057), .Y(n_1056) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVxp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
CKINVDCx5p33_ASAP7_75t_R g1060 ( .A(n_1061), .Y(n_1060) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1065), .Y(n_1094) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1072), .Y(n_1065) );
AND4x1_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1068), .C(n_1069), .D(n_1070), .Y(n_1066) );
NOR3xp33_ASAP7_75t_L g1072 ( .A(n_1073), .B(n_1077), .C(n_1080), .Y(n_1072) );
OAI21xp33_ASAP7_75t_L g1080 ( .A1(n_1081), .A2(n_1082), .B(n_1083), .Y(n_1080) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
HB1xp67_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
BUFx2_ASAP7_75t_SL g1090 ( .A(n_1091), .Y(n_1090) );
HB1xp67_ASAP7_75t_L g1095 ( .A(n_1096), .Y(n_1095) );
endmodule