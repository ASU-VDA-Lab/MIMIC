module fake_jpeg_23522_n_136 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_27),
.B(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_39),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

NOR2x1p5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_1),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_48),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_28),
.B1(n_21),
.B2(n_29),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_28),
.B1(n_29),
.B2(n_19),
.Y(n_68)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_17),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_49),
.B(n_56),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_32),
.Y(n_66)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_18),
.Y(n_55)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_26),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_44),
.B(n_42),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_66),
.B(n_71),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_49),
.Y(n_85)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_63),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_33),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_73),
.B1(n_20),
.B2(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_53),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_36),
.B1(n_28),
.B2(n_31),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_43),
.B1(n_51),
.B2(n_46),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_33),
.C(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_20),
.B1(n_25),
.B2(n_22),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_48),
.B1(n_54),
.B2(n_43),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_79),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_81),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_60),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_49),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_66),
.B1(n_58),
.B2(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_84),
.B1(n_85),
.B2(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_59),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_97),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_59),
.B(n_68),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_98),
.B(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_71),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_86),
.A2(n_61),
.B(n_73),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_70),
.B(n_24),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_26),
.B(n_22),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_74),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_89),
.C(n_88),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_108),
.B(n_109),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_110),
.B(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_88),
.Y(n_109)
);

FAx1_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_82),
.CI(n_76),
.CON(n_110),
.SN(n_110)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_106),
.A2(n_97),
.A3(n_93),
.B1(n_101),
.B2(n_95),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_7),
.B1(n_11),
.B2(n_10),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_91),
.C(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_116),
.C(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_74),
.C(n_23),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_15),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_119)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_103),
.B(n_112),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_5),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_1),
.B(n_2),
.C(n_4),
.Y(n_122)
);

OAI21x1_ASAP7_75t_SL g124 ( 
.A1(n_118),
.A2(n_2),
.B(n_4),
.Y(n_124)
);

OA21x2_ASAP7_75t_SL g127 ( 
.A1(n_124),
.A2(n_9),
.B(n_12),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_125),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_127),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_123),
.B(n_122),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_128),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_120),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_129),
.B(n_131),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule