module real_jpeg_18764_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_0),
.A2(n_15),
.B(n_451),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_0),
.B(n_452),
.Y(n_451)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_1),
.A2(n_68),
.A3(n_71),
.B1(n_74),
.B2(n_80),
.Y(n_67)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_1),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_1),
.B(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_1),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_1),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_1),
.A2(n_43),
.B1(n_225),
.B2(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_2),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_2),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_3),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_133),
.B1(n_161),
.B2(n_164),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_3),
.A2(n_133),
.B1(n_174),
.B2(n_176),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_3),
.A2(n_22),
.B1(n_133),
.B2(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_4),
.Y(n_159)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_4),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_4),
.Y(n_199)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_5),
.A2(n_46),
.B1(n_174),
.B2(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_6),
.A2(n_53),
.B1(n_301),
.B2(n_303),
.Y(n_300)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_6),
.A2(n_53),
.B1(n_321),
.B2(n_324),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_6),
.A2(n_53),
.B1(n_424),
.B2(n_425),
.Y(n_423)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_7),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_7),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_7),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_8),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_8),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_8),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_8),
.Y(n_323)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_9),
.Y(n_452)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_12),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_12),
.Y(n_94)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_12),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g266 ( 
.A(n_13),
.Y(n_266)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_13),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_58),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_57),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_54),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_18),
.B(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_18),
.B(n_444),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B1(n_40),
.B2(n_50),
.Y(n_18)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_19),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_20),
.B(n_31),
.Y(n_56)
);

OA22x2_ASAP7_75t_L g262 ( 
.A1(n_20),
.A2(n_31),
.B1(n_263),
.B2(n_267),
.Y(n_262)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_20),
.A2(n_31),
.B1(n_263),
.B2(n_267),
.Y(n_294)
);

OAI21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_27),
.B(n_31),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_21),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_24),
.Y(n_21)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_31),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_31),
.A2(n_40),
.B(n_439),
.Y(n_438)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_31)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_32),
.Y(n_406)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_32),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_33),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_33),
.Y(n_284)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_46),
.A2(n_75),
.B1(n_315),
.B2(n_317),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_46),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_47),
.B(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_50),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_56),
.B(n_336),
.Y(n_335)
);

OA21x2_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_390),
.B(n_445),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AO221x1_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_289),
.B1(n_291),
.B2(n_383),
.C(n_389),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_251),
.B(n_288),
.Y(n_61)
);

AOI21x1_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_234),
.B(n_250),
.Y(n_62)
);

OAI21x1_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_182),
.B(n_233),
.Y(n_63)
);

NOR2xp67_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_168),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_65),
.B(n_168),
.Y(n_233)
);

XOR2x2_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_107),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_66),
.B(n_137),
.C(n_166),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_86),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_67),
.B(n_86),
.Y(n_237)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_77),
.Y(n_325)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_79),
.B(n_143),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_79),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_84),
.Y(n_80)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_95),
.Y(n_86)
);

OA22x2_ASAP7_75t_L g171 ( 
.A1(n_87),
.A2(n_172),
.B1(n_173),
.B2(n_178),
.Y(n_171)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_88),
.B(n_96),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_89),
.A2(n_139),
.B(n_142),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g155 ( 
.A1(n_91),
.A2(n_151),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_91),
.Y(n_175)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_91),
.Y(n_214)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_91),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_94),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g333 ( 
.A(n_95),
.B(n_300),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_96),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_99),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_100),
.Y(n_191)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_103),
.A2(n_173),
.B(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_106),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_137),
.B1(n_166),
.B2(n_167),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_108),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_108),
.A2(n_166),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_108),
.B(n_294),
.C(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_108),
.A2(n_166),
.B1(n_294),
.B2(n_341),
.Y(n_340)
);

OA22x2_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_116),
.B1(n_122),
.B2(n_129),
.Y(n_108)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_109),
.A2(n_116),
.B1(n_122),
.B2(n_129),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_109),
.A2(n_116),
.B(n_122),
.Y(n_354)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_109),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_109),
.B(n_116),
.Y(n_437)
);

NAND2x1p5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_116),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_122),
.Y(n_401)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_126),
.Y(n_426)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx2_ASAP7_75t_SL g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_136),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_137),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_137),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_137),
.A2(n_167),
.B1(n_185),
.B2(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_137),
.B(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_137),
.A2(n_167),
.B1(n_347),
.B2(n_375),
.Y(n_374)
);

AO22x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_145),
.B1(n_155),
.B2(n_160),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_145),
.B1(n_155),
.B2(n_160),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_138),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_138),
.B(n_312),
.Y(n_330)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_186),
.A3(n_190),
.B1(n_192),
.B2(n_197),
.Y(n_185)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_145),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_145),
.Y(n_312)
);

NOR2x1p5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_149),
.Y(n_319)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_155),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_155),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_155),
.A2(n_312),
.B1(n_313),
.B2(n_320),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_157),
.Y(n_305)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_166),
.B(n_257),
.C(n_378),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_180),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_169),
.A2(n_170),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_169),
.B(n_237),
.C(n_239),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_169),
.A2(n_170),
.B1(n_296),
.B2(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_180),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_170),
.B(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_223),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_171),
.A2(n_204),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_172),
.A2(n_297),
.B1(n_300),
.B2(n_306),
.Y(n_296)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_181),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_181),
.A2(n_402),
.B1(n_403),
.B2(n_423),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_207),
.B(n_232),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_203),
.Y(n_183)
);

NOR2xp67_ASAP7_75t_SL g232 ( 
.A(n_184),
.B(n_203),
.Y(n_232)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_204),
.B(n_275),
.Y(n_365)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_227),
.B(n_231),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_222),
.B(n_226),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_220),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_228),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_220),
.B(n_241),
.C(n_245),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_221),
.A2(n_297),
.B(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_249),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_249),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_248),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_236),
.Y(n_248)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_243),
.B2(n_247),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_241),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_241),
.A2(n_311),
.B(n_326),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_241),
.B(n_311),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_241),
.B(n_294),
.C(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_241),
.A2(n_247),
.B1(n_294),
.B2(n_341),
.Y(n_371)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_253),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_271),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_254),
.B(n_272),
.C(n_273),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_258),
.B(n_259),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_259),
.A2(n_314),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_261),
.A2(n_262),
.B1(n_353),
.B2(n_354),
.Y(n_360)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_262),
.Y(n_378)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_263),
.Y(n_336)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_366),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_355),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_338),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_292),
.B(n_338),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_309),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_293),
.B(n_310),
.C(n_327),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_294),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_294),
.A2(n_341),
.B1(n_419),
.B2(n_420),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_294),
.B(n_398),
.C(n_442),
.Y(n_441)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_295),
.B(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_327),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_315),
.A2(n_316),
.B1(n_404),
.B2(n_407),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_320),
.B(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_326),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_326),
.A2(n_394),
.B1(n_410),
.B2(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_334),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g412 ( 
.A(n_328),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.Y(n_328)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_329),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_331),
.A2(n_332),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_333),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_332),
.A2(n_337),
.B(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_336),
.B(n_440),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.C(n_345),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_339),
.B(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_345),
.B(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.C(n_353),
.Y(n_345)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_346),
.B(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_347),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_352),
.B(n_400),
.C(n_415),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_352),
.A2(n_395),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_355),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_356),
.B(n_358),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.C(n_364),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_362),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

XNOR2x1_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_365),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_379),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_369),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_370),
.B(n_374),
.C(n_376),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_376),
.B2(n_377),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_378),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_378),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_378),
.B(n_414),
.C(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_386),
.Y(n_385)
);

NAND2x1_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_382),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_382),
.Y(n_384)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_385),
.B(n_387),
.C(n_388),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_432),
.C(n_443),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_427),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_392),
.A2(n_447),
.B(n_448),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_413),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_393),
.B(n_413),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_410),
.C(n_411),
.Y(n_393)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_398),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_398),
.A2(n_415),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_407),
.Y(n_424)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_430),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVxp33_ASAP7_75t_L g434 ( 
.A(n_418),
.Y(n_434)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_429),
.Y(n_447)
);

A2O1A1O1Ixp25_ASAP7_75t_L g445 ( 
.A1(n_432),
.A2(n_443),
.B(n_446),
.C(n_449),
.D(n_450),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_435),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_435),
.Y(n_449)
);

BUFx24_ASAP7_75t_SL g454 ( 
.A(n_435),
.Y(n_454)
);

FAx1_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_438),
.CI(n_441),
.CON(n_435),
.SN(n_435)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_438),
.C(n_441),
.Y(n_444)
);


endmodule