module fake_jpeg_30050_n_517 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_517);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_517;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx10_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_16),
.B(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_53),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_54),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_55),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_64),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_68),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_98),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_9),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_84),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_76),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_27),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_77),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_82),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_83),
.B(n_86),
.Y(n_164)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_94),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_9),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_39),
.B(n_6),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_38),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_100),
.B(n_103),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_72),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_111),
.B(n_112),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_57),
.A2(n_32),
.B(n_48),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_115),
.B(n_133),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_139),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_54),
.A2(n_36),
.B1(n_37),
.B2(n_47),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_127),
.A2(n_140),
.B1(n_142),
.B2(n_18),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_54),
.A2(n_32),
.B(n_48),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_82),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_40),
.B1(n_39),
.B2(n_44),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_55),
.B(n_40),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_144),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_85),
.A2(n_15),
.B1(n_43),
.B2(n_46),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_55),
.B(n_44),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_53),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_149),
.B(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_83),
.B(n_42),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_49),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_99),
.B(n_42),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_86),
.A2(n_45),
.B(n_35),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_49),
.Y(n_187)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_119),
.A2(n_92),
.B1(n_97),
.B2(n_96),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_167),
.A2(n_177),
.B1(n_78),
.B2(n_58),
.Y(n_237)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_169),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_124),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_179),
.Y(n_216)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_172),
.Y(n_247)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_174),
.Y(n_221)
);

BUFx16f_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_175),
.Y(n_243)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_176),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_119),
.A2(n_101),
.B1(n_90),
.B2(n_81),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_196),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_156),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_182),
.A2(n_184),
.B1(n_185),
.B2(n_191),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_36),
.B1(n_34),
.B2(n_45),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_148),
.A2(n_52),
.B1(n_47),
.B2(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_192),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_105),
.Y(n_188)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_116),
.A2(n_47),
.B1(n_37),
.B2(n_61),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_122),
.B(n_0),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_135),
.C(n_22),
.Y(n_227)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_197),
.Y(n_230)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_113),
.B(n_47),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_159),
.Y(n_197)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_208),
.Y(n_226)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_202),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_107),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_201),
.A2(n_209),
.B1(n_210),
.B2(n_212),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_106),
.B(n_47),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_134),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_206),
.Y(n_241)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

NAND2xp33_ASAP7_75t_R g239 ( 
.A(n_207),
.B(n_142),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_116),
.A2(n_61),
.B1(n_63),
.B2(n_43),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_155),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_213),
.B(n_180),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_170),
.B(n_106),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_229),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_183),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_170),
.B(n_208),
.C(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_228),
.B(n_203),
.C(n_200),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_145),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_235),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_168),
.B(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_194),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_175),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_153),
.B1(n_143),
.B2(n_118),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_SL g238 ( 
.A(n_178),
.B(n_114),
.C(n_127),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_155),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_239),
.A2(n_242),
.B1(n_165),
.B2(n_129),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_181),
.A2(n_143),
.B1(n_153),
.B2(n_145),
.Y(n_242)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_169),
.A2(n_136),
.B1(n_120),
.B2(n_128),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_199),
.B(n_146),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx13_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_253),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_255),
.B(n_257),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g256 ( 
.A(n_215),
.B(n_186),
.CI(n_171),
.CON(n_256),
.SN(n_256)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_256),
.B(n_260),
.Y(n_309)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_217),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_229),
.B(n_179),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_263),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_281),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_215),
.B(n_197),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_217),
.B(n_213),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_264),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_204),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_266),
.B(n_267),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_234),
.B(n_166),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_176),
.Y(n_268)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_245),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_270),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_271),
.A2(n_246),
.B1(n_198),
.B2(n_209),
.Y(n_289)
);

INVx11_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_272),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_279),
.C(n_240),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_211),
.Y(n_274)
);

O2A1O1Ixp33_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_241),
.B(n_223),
.C(n_243),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_215),
.B(n_206),
.Y(n_275)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_275),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_276),
.A2(n_242),
.B1(n_244),
.B2(n_226),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_214),
.A2(n_205),
.B(n_175),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_262),
.B(n_232),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_180),
.B(n_104),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_228),
.B(n_22),
.C(n_18),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_219),
.B(n_189),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_230),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_282),
.A2(n_285),
.B1(n_291),
.B2(n_307),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_244),
.B(n_219),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_284),
.B(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_230),
.B1(n_249),
.B2(n_250),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_302),
.B(n_277),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_289),
.A2(n_270),
.B1(n_266),
.B2(n_245),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_261),
.A2(n_230),
.B1(n_249),
.B2(n_241),
.Y(n_291)
);

AOI211xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_216),
.B(n_227),
.C(n_223),
.Y(n_292)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_292),
.A2(n_257),
.B(n_256),
.C(n_279),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_252),
.A2(n_274),
.B1(n_281),
.B2(n_275),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_295),
.A2(n_312),
.B1(n_278),
.B2(n_280),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_254),
.Y(n_297)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_232),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_268),
.B(n_233),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_305),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_269),
.A2(n_220),
.B1(n_137),
.B2(n_132),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_273),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_267),
.B(n_265),
.Y(n_330)
);

OAI22x1_ASAP7_75t_SL g312 ( 
.A1(n_278),
.A2(n_221),
.B1(n_218),
.B2(n_147),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_313),
.Y(n_350)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_309),
.B(n_264),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_315),
.B(n_321),
.Y(n_365)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_317),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_318),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_287),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_319),
.B(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_263),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_324),
.B(n_340),
.C(n_285),
.Y(n_375)
);

AND2x6_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_254),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_326),
.B(n_327),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_287),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_256),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_335),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_329),
.A2(n_289),
.B1(n_306),
.B2(n_288),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_331),
.B(n_293),
.Y(n_345)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_304),
.Y(n_332)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_283),
.Y(n_334)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_334),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_258),
.B1(n_270),
.B2(n_272),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_290),
.B(n_255),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_337),
.Y(n_352)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_305),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_338),
.Y(n_368)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_339),
.B(n_343),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_279),
.C(n_233),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_296),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_309),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_303),
.A2(n_247),
.B1(n_235),
.B2(n_253),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_290),
.B(n_298),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_284),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_345),
.B(n_351),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_324),
.B(n_295),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_348),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_340),
.B(n_294),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_336),
.B(n_293),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_355),
.A2(n_342),
.B1(n_311),
.B2(n_307),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_358),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_320),
.B(n_298),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_363),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_320),
.B(n_310),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_331),
.B(n_310),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_366),
.B(n_18),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_344),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_323),
.A2(n_306),
.B1(n_303),
.B2(n_292),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_369),
.A2(n_374),
.B1(n_221),
.B2(n_210),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_291),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_372),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_325),
.A2(n_303),
.B1(n_284),
.B2(n_282),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_375),
.B(n_338),
.C(n_343),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_376),
.Y(n_391)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_357),
.Y(n_377)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_377),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_375),
.B(n_322),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_385),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_379),
.B(n_383),
.C(n_384),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_381),
.A2(n_404),
.B1(n_362),
.B2(n_350),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_349),
.A2(n_326),
.B1(n_328),
.B2(n_342),
.Y(n_382)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_382),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_347),
.B(n_334),
.C(n_333),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_366),
.C(n_369),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_330),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_317),
.C(n_316),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_396),
.C(n_373),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_316),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_388),
.B(n_399),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_349),
.A2(n_339),
.B1(n_332),
.B2(n_318),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_389),
.A2(n_362),
.B1(n_350),
.B2(n_221),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_353),
.A2(n_300),
.B1(n_299),
.B2(n_301),
.Y(n_390)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_376),
.A2(n_300),
.B(n_299),
.Y(n_392)
);

AO21x1_ASAP7_75t_L g422 ( 
.A1(n_392),
.A2(n_259),
.B(n_251),
.Y(n_422)
);

MAJx2_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_247),
.C(n_251),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_393),
.B(n_402),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_356),
.B(n_248),
.C(n_236),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_354),
.A2(n_355),
.B1(n_346),
.B2(n_352),
.Y(n_397)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_351),
.B(n_248),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_371),
.A2(n_188),
.B1(n_190),
.B2(n_201),
.Y(n_403)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_403),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_413),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_377),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_410),
.B(n_417),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_371),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_407),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_401),
.A2(n_368),
.B1(n_361),
.B2(n_370),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_412),
.A2(n_125),
.B1(n_146),
.B2(n_158),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_367),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_364),
.C(n_359),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_428),
.C(n_402),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_416),
.A2(n_389),
.B1(n_394),
.B2(n_396),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_391),
.A2(n_394),
.B(n_392),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_398),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_422),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_421),
.A2(n_120),
.B1(n_137),
.B2(n_132),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_379),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_386),
.Y(n_431)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_393),
.Y(n_426)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_426),
.Y(n_429)
);

AO21x1_ASAP7_75t_L g427 ( 
.A1(n_380),
.A2(n_259),
.B(n_180),
.Y(n_427)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_427),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_240),
.C(n_174),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_431),
.B(n_439),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_409),
.Y(n_432)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

NOR2xp67_ASAP7_75t_SL g433 ( 
.A(n_408),
.B(n_387),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_433),
.B(n_446),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_434),
.B(n_437),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_385),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_404),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_387),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_441),
.A2(n_445),
.B1(n_415),
.B2(n_56),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_428),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_395),
.C(n_195),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_449),
.C(n_406),
.Y(n_452)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_444),
.B(n_147),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_424),
.A2(n_118),
.B1(n_165),
.B2(n_129),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_447),
.A2(n_425),
.B1(n_422),
.B2(n_162),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_405),
.B(n_172),
.C(n_128),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_451),
.B(n_456),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_452),
.B(n_461),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_414),
.C(n_413),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_464),
.C(n_447),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_443),
.B(n_420),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_416),
.C(n_419),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_460),
.Y(n_469)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_459),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_448),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_415),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_440),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_158),
.C(n_138),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_465),
.B(n_466),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_125),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_147),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_467),
.B(n_24),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_483),
.C(n_474),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_463),
.A2(n_436),
.B(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_455),
.A2(n_435),
.B(n_438),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_472),
.A2(n_11),
.B(n_14),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_474),
.B(n_475),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_454),
.A2(n_432),
.B(n_138),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g476 ( 
.A1(n_452),
.A2(n_162),
.B(n_151),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_477),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_464),
.A2(n_77),
.B(n_75),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_479),
.A2(n_46),
.B1(n_12),
.B2(n_14),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_453),
.A2(n_74),
.B1(n_67),
.B2(n_66),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_481),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_462),
.B(n_11),
.CI(n_12),
.CON(n_481),
.SN(n_481)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_46),
.C(n_15),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_473),
.A2(n_450),
.B(n_458),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_485),
.B(n_490),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_478),
.A2(n_458),
.B1(n_15),
.B2(n_12),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_487),
.Y(n_497)
);

AOI31xp67_ASAP7_75t_L g489 ( 
.A1(n_472),
.A2(n_11),
.A3(n_14),
.B(n_3),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_489),
.A2(n_482),
.B(n_10),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_46),
.C(n_23),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_493),
.B(n_494),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_469),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_495),
.B(n_477),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_484),
.B(n_481),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_499),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_470),
.C(n_476),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_502),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_488),
.B(n_483),
.C(n_24),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g506 ( 
.A1(n_503),
.A2(n_491),
.B(n_492),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_SL g505 ( 
.A(n_496),
.B(n_489),
.Y(n_505)
);

AOI322xp5_ASAP7_75t_L g509 ( 
.A1(n_505),
.A2(n_496),
.A3(n_500),
.B1(n_493),
.B2(n_6),
.C1(n_10),
.C2(n_0),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_506),
.B(n_508),
.C(n_24),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_486),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_509),
.A2(n_510),
.B(n_1),
.Y(n_513)
);

AOI322xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_23),
.C1(n_24),
.C2(n_504),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_1),
.B(n_2),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g514 ( 
.A1(n_512),
.A2(n_513),
.B1(n_1),
.B2(n_23),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_23),
.C(n_24),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_515),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_23),
.Y(n_517)
);


endmodule