module fake_netlist_1_12425_n_35 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
HB1xp67_ASAP7_75t_L g14 ( .A(n_7), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_0), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_13), .B(n_3), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_4), .B(n_8), .Y(n_17) );
AOI22xp5_ASAP7_75t_L g18 ( .A1(n_0), .A2(n_3), .B1(n_9), .B2(n_11), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_10), .B(n_2), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_1), .Y(n_20) );
INVx4_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_14), .Y(n_22) );
BUFx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_23), .B(n_15), .Y(n_26) );
INVx4_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_27), .B(n_25), .Y(n_28) );
NOR3xp33_ASAP7_75t_L g29 ( .A(n_28), .B(n_21), .C(n_18), .Y(n_29) );
AOI22xp5_ASAP7_75t_SL g30 ( .A1(n_28), .A2(n_16), .B1(n_19), .B2(n_20), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
NAND3xp33_ASAP7_75t_L g32 ( .A(n_29), .B(n_17), .C(n_6), .Y(n_32) );
BUFx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
OAI22xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_32), .B1(n_5), .B2(n_12), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
endmodule