module fake_jpeg_165_n_90 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_4),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

CKINVDCx6p67_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_35),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_9),
.C(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_25),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_47),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_51),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_35),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_31),
.B(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_37),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_34),
.B1(n_26),
.B2(n_24),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_54),
.B(n_29),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g54 ( 
.A(n_46),
.B(n_36),
.C(n_30),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_31),
.B(n_32),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_55),
.A2(n_44),
.B(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_41),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_37),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_48),
.C(n_45),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_63),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_62),
.B(n_43),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_44),
.B(n_37),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_27),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_26),
.B1(n_24),
.B2(n_43),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_73),
.B(n_75),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_62),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_64),
.Y(n_72)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_66),
.A2(n_22),
.B(n_20),
.C(n_19),
.D(n_18),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_17),
.C(n_16),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_77),
.C(n_80),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_11),
.C(n_2),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_1),
.C(n_2),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_74),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_71),
.C(n_5),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_3),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_4),
.B(n_5),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_85),
.B(n_83),
.Y(n_86)
);

NOR2xp67_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_6),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_88),
.A2(n_6),
.B(n_7),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_7),
.C(n_8),
.Y(n_90)
);


endmodule