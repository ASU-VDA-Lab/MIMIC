module fake_netlist_6_3995_n_1766 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1766);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1766;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_83),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_35),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_32),
.Y(n_166)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_31),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_16),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_16),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_63),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_91),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_15),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_35),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_67),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_33),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_116),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_70),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_8),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_109),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_25),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_57),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_74),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_138),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_84),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_66),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_22),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_69),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_118),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_86),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_99),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_163),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_79),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_8),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_43),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_68),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_101),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_142),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_42),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_85),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_161),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_55),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_75),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_34),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_71),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_4),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_139),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_100),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_155),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_157),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_33),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_15),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_41),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_53),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_156),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_128),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_104),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_48),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_132),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_13),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_60),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_22),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_111),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_105),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_58),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_94),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_117),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_17),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_131),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_125),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_73),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_152),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_119),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_24),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_52),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_65),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_48),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_81),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_96),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_122),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_141),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_31),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_59),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_54),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_129),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_0),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_44),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_21),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_124),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_150),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_0),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_87),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_112),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_82),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_29),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_10),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_115),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_29),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_52),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_93),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_1),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_90),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_103),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_2),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_123),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_26),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_154),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_18),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_114),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_97),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_78),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_36),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_34),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_23),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_92),
.Y(n_298)
);

INVxp33_ASAP7_75t_L g299 ( 
.A(n_25),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_27),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_50),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_158),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_14),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_49),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_153),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_108),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_46),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_121),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_20),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_135),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_77),
.Y(n_315)
);

INVxp67_ASAP7_75t_SL g316 ( 
.A(n_41),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_6),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_45),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_148),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_38),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_19),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_10),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_146),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_107),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

INVx2_ASAP7_75t_SL g327 ( 
.A(n_51),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_151),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_18),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_160),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_61),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_32),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_170),
.B(n_2),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_164),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_170),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_302),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_171),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_172),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_200),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_211),
.B(n_3),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_224),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_178),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_224),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_176),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_165),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_193),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_241),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_165),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_180),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_183),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_223),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_277),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_210),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_277),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_169),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_241),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_187),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_188),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_169),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_4),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_174),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_174),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_235),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_211),
.B(n_5),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_189),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_255),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_175),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_190),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_175),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_236),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_247),
.Y(n_378)
);

NOR2xp67_ASAP7_75t_L g379 ( 
.A(n_327),
.B(n_5),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_181),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_195),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_196),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_245),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_307),
.B(n_6),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_181),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_307),
.B(n_7),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_201),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_202),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_203),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_255),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_204),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_223),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_205),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_231),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_271),
.Y(n_395)
);

NOR2xp67_ASAP7_75t_L g396 ( 
.A(n_231),
.B(n_9),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_244),
.B(n_9),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_244),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_206),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_248),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_209),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_248),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_256),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_256),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_272),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_212),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_287),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_271),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_272),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_245),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_295),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_235),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_220),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_221),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_225),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_334),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_337),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_362),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_366),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_179),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_345),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_341),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_335),
.B(n_299),
.Y(n_429)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_348),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_354),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_363),
.B(n_227),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_R g436 ( 
.A(n_382),
.B(n_228),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_410),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_410),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_369),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_355),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_369),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_360),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_336),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_338),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_338),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_339),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_353),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_376),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_376),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_364),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_339),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_340),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_365),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_344),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_344),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_351),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_380),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_350),
.B(n_287),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_346),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_394),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_372),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_346),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_375),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_381),
.B(n_173),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_347),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_R g475 ( 
.A(n_387),
.B(n_168),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_392),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_400),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_359),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_347),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_395),
.B(n_229),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_388),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_391),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

CKINVDCx16_ASAP7_75t_R g484 ( 
.A(n_357),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_349),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_393),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_402),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_349),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_357),
.B(n_199),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_399),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_401),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_402),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_395),
.B(n_232),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_426),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_426),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_434),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_436),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_430),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_484),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_429),
.A2(n_333),
.B1(n_343),
.B2(n_384),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_SL g501 ( 
.A1(n_434),
.A2(n_386),
.B1(n_342),
.B2(n_371),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_245),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_425),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_417),
.B(n_352),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_425),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_471),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_418),
.A2(n_416),
.B1(n_389),
.B2(n_414),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_426),
.Y(n_509)
);

NAND2xp33_ASAP7_75t_L g510 ( 
.A(n_480),
.B(n_245),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_493),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_475),
.A2(n_406),
.B1(n_413),
.B2(n_407),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_428),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_430),
.B(n_179),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_428),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_437),
.Y(n_519)
);

CKINVDCx8_ASAP7_75t_R g520 ( 
.A(n_484),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_493),
.B(n_182),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_476),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_419),
.B(n_373),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_420),
.B(n_390),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_420),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_432),
.B(n_408),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_447),
.B(n_395),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_421),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

NAND2xp33_ASAP7_75t_L g535 ( 
.A(n_428),
.B(n_245),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_433),
.B(n_182),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_424),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_424),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_438),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_489),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_447),
.B(n_425),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_428),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_448),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_447),
.B(n_186),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_463),
.B(n_367),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_440),
.B(n_186),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_465),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_431),
.B(n_370),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_447),
.B(n_197),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_448),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_431),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_435),
.B(n_412),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_435),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_423),
.Y(n_556)
);

BUFx4f_ASAP7_75t_L g557 ( 
.A(n_448),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_465),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_442),
.B(n_197),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_465),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_439),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_452),
.B(n_370),
.C(n_379),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_439),
.A2(n_397),
.B1(n_396),
.B2(n_301),
.Y(n_563)
);

BUFx8_ASAP7_75t_SL g564 ( 
.A(n_460),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_448),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_456),
.B(n_356),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_422),
.B(n_218),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_441),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_467),
.B(n_356),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_441),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_443),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_444),
.B(n_358),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_448),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_444),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_450),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_450),
.B(n_358),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_465),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_469),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_470),
.B(n_286),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_451),
.B(n_361),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_451),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_481),
.A2(n_313),
.B1(n_316),
.B2(n_213),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_478),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_422),
.B(n_284),
.Y(n_586)
);

INVx1_ASAP7_75t_SL g587 ( 
.A(n_482),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_492),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_453),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_445),
.B(n_361),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_486),
.B(n_377),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_453),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_461),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_469),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_492),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_469),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_462),
.A2(n_311),
.B1(n_297),
.B2(n_301),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_445),
.B(n_233),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_490),
.A2(n_378),
.B1(n_166),
.B2(n_278),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_469),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_491),
.B(n_286),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_462),
.B(n_177),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_473),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_464),
.Y(n_605)
);

OAI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_464),
.A2(n_264),
.B1(n_298),
.B2(n_258),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_473),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_446),
.B(n_454),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_466),
.Y(n_609)
);

AND2x6_ASAP7_75t_L g610 ( 
.A(n_446),
.B(n_289),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_466),
.B(n_403),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_468),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_472),
.A2(n_297),
.B1(n_311),
.B2(n_326),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_472),
.B(n_184),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_474),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_474),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_492),
.B(n_289),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_446),
.B(n_222),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_477),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_473),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_477),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_483),
.B(n_191),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_483),
.B(n_192),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_454),
.Y(n_626)
);

OAI21xp33_ASAP7_75t_SL g627 ( 
.A1(n_487),
.A2(n_194),
.B(n_192),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_487),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_458),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_454),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_455),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_458),
.B(n_208),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_455),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_455),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_457),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_457),
.A2(n_269),
.B1(n_268),
.B2(n_267),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_457),
.A2(n_250),
.B1(n_265),
.B2(n_331),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_458),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_459),
.B(n_234),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_459),
.Y(n_640)
);

OAI21xp33_ASAP7_75t_SL g641 ( 
.A1(n_459),
.A2(n_274),
.B(n_194),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_550),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_496),
.B(n_198),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_554),
.B(n_167),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_496),
.B(n_198),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_512),
.B(n_207),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_512),
.B(n_567),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_501),
.B(n_222),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_621),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_640),
.B(n_553),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_594),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_640),
.B(n_207),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_611),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_611),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_516),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_621),
.B(n_403),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_572),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_553),
.B(n_214),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_561),
.B(n_629),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_580),
.B(n_222),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_561),
.B(n_214),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_524),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_505),
.B(n_216),
.Y(n_664)
);

INVx8_ASAP7_75t_L g665 ( 
.A(n_547),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_500),
.B(n_245),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g667 ( 
.A1(n_504),
.A2(n_528),
.B1(n_554),
.B2(n_570),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_525),
.B(n_217),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_504),
.A2(n_270),
.B1(n_239),
.B2(n_240),
.Y(n_669)
);

O2A1O1Ixp5_ASAP7_75t_L g670 ( 
.A1(n_517),
.A2(n_522),
.B(n_597),
.C(n_580),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_606),
.A2(n_613),
.B(n_522),
.C(n_510),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_588),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_594),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_528),
.B(n_230),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_541),
.A2(n_292),
.B(n_258),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_623),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_516),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_564),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_494),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_513),
.B(n_237),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_580),
.B(n_222),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_623),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_578),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_556),
.B(n_524),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_634),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_529),
.B(n_237),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_578),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_532),
.B(n_264),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_625),
.A2(n_510),
.B1(n_502),
.B2(n_544),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_497),
.B(n_215),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_533),
.B(n_273),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_544),
.B(n_245),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_537),
.B(n_273),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_516),
.Y(n_694)
);

INVx4_ASAP7_75t_L g695 ( 
.A(n_516),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_507),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_597),
.B(n_222),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_597),
.B(n_245),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_582),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_582),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_514),
.B(n_242),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_503),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_494),
.Y(n_703)
);

INVxp67_ASAP7_75t_L g704 ( 
.A(n_530),
.Y(n_704)
);

INVx8_ASAP7_75t_L g705 ( 
.A(n_547),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_506),
.B(n_219),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_538),
.B(n_274),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_555),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_574),
.Y(n_709)
);

AOI221xp5_ASAP7_75t_L g710 ( 
.A1(n_584),
.A2(n_246),
.B1(n_226),
.B2(n_326),
.C(n_332),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_506),
.B(n_238),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_506),
.B(n_253),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_634),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_544),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_569),
.B(n_283),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_571),
.B(n_283),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_625),
.A2(n_332),
.B1(n_292),
.B2(n_315),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_536),
.B(n_254),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_547),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_573),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_495),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_576),
.B(n_298),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_577),
.Y(n_723)
);

AND2x6_ASAP7_75t_SL g724 ( 
.A(n_591),
.B(n_404),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_625),
.A2(n_320),
.B1(n_315),
.B2(n_324),
.Y(n_725)
);

NOR2x1p5_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_259),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_L g727 ( 
.A1(n_517),
.A2(n_324),
.B(n_320),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_583),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_498),
.B(n_245),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_589),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_508),
.B(n_243),
.Y(n_731)
);

INVx5_ASAP7_75t_L g732 ( 
.A(n_544),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_605),
.B(n_167),
.Y(n_733)
);

NOR2xp67_ASAP7_75t_L g734 ( 
.A(n_600),
.B(n_249),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_544),
.B(n_251),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_592),
.B(n_479),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_498),
.B(n_252),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_605),
.B(n_257),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_509),
.Y(n_739)
);

INVx2_ASAP7_75t_SL g740 ( 
.A(n_605),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_536),
.B(n_262),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_595),
.B(n_260),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_499),
.B(n_404),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_593),
.B(n_479),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_609),
.B(n_485),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_502),
.A2(n_167),
.B1(n_415),
.B2(n_411),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_595),
.B(n_261),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_551),
.A2(n_167),
.B1(n_415),
.B2(n_411),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_601),
.B(n_263),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_548),
.B(n_266),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_612),
.B(n_485),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_616),
.B(n_485),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_617),
.B(n_488),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_551),
.A2(n_405),
.B1(n_409),
.B2(n_306),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_SL g755 ( 
.A1(n_548),
.A2(n_305),
.B1(n_276),
.B2(n_279),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_601),
.B(n_275),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_604),
.B(n_281),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_628),
.B(n_488),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_604),
.B(n_288),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_626),
.B(n_488),
.Y(n_760)
);

AND2x6_ASAP7_75t_SL g761 ( 
.A(n_547),
.B(n_405),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_551),
.B(n_293),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_607),
.B(n_294),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_551),
.A2(n_409),
.B1(n_310),
.B2(n_329),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_607),
.B(n_330),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_626),
.B(n_328),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_559),
.B(n_280),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_626),
.Y(n_768)
);

INVxp67_ASAP7_75t_L g769 ( 
.A(n_540),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_618),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_568),
.B(n_325),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_599),
.B(n_308),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_559),
.B(n_323),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_304),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_618),
.Y(n_775)
);

NOR2x1p5_ASAP7_75t_L g776 ( 
.A(n_585),
.B(n_322),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_581),
.B(n_321),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_632),
.B(n_312),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_622),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_581),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_622),
.B(n_314),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_602),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_586),
.B(n_319),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_531),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_602),
.Y(n_785)
);

NOR3xp33_ASAP7_75t_L g786 ( 
.A(n_523),
.B(n_318),
.C(n_309),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_588),
.B(n_303),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_596),
.B(n_300),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_596),
.B(n_296),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_511),
.Y(n_790)
);

INVxp33_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_587),
.B(n_290),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_585),
.B(n_291),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_596),
.B(n_285),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_563),
.B(n_162),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_603),
.B(n_282),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_627),
.A2(n_598),
.B(n_614),
.C(n_615),
.Y(n_797)
);

INVx4_ASAP7_75t_L g798 ( 
.A(n_534),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_L g799 ( 
.A(n_796),
.B(n_668),
.C(n_710),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_647),
.B(n_526),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_L g801 ( 
.A1(n_796),
.A2(n_624),
.B(n_636),
.Y(n_801)
);

OAI21x1_ASAP7_75t_L g802 ( 
.A1(n_670),
.A2(n_558),
.B(n_545),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_714),
.Y(n_803)
);

OAI22xp5_ASAP7_75t_L g804 ( 
.A1(n_647),
.A2(n_667),
.B1(n_768),
.B2(n_651),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_663),
.B(n_526),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_704),
.B(n_596),
.Y(n_806)
);

NOR2x1_ASAP7_75t_L g807 ( 
.A(n_776),
.B(n_590),
.Y(n_807)
);

AO22x1_ASAP7_75t_L g808 ( 
.A1(n_668),
.A2(n_551),
.B1(n_520),
.B2(n_610),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_SL g809 ( 
.A(n_678),
.B(n_526),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_666),
.A2(n_637),
.B(n_641),
.C(n_638),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_768),
.A2(n_521),
.B(n_557),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_795),
.B(n_520),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_689),
.A2(n_557),
.B1(n_521),
.B2(n_549),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_672),
.A2(n_557),
.B(n_521),
.Y(n_814)
);

O2A1O1Ixp33_ASAP7_75t_SL g815 ( 
.A1(n_797),
.A2(n_620),
.B(n_619),
.C(n_608),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_689),
.A2(n_545),
.B1(n_558),
.B2(n_560),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_684),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_760),
.A2(n_729),
.B(n_798),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_798),
.A2(n_565),
.B(n_552),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_650),
.B(n_518),
.Y(n_820)
);

OAI21xp33_ASAP7_75t_L g821 ( 
.A1(n_718),
.A2(n_619),
.B(n_620),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_656),
.A2(n_552),
.B(n_565),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_702),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_795),
.B(n_542),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_780),
.B(n_542),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_644),
.B(n_631),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_650),
.B(n_546),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_656),
.A2(n_546),
.B(n_518),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_743),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_L g830 ( 
.A1(n_784),
.A2(n_511),
.B(n_515),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_792),
.B(n_633),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_660),
.B(n_575),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_677),
.A2(n_575),
.B(n_534),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_677),
.A2(n_534),
.B(n_542),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_694),
.A2(n_534),
.B(n_542),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_694),
.A2(n_579),
.B(n_543),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_718),
.B(n_535),
.C(n_635),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_695),
.A2(n_766),
.B(n_732),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_782),
.B(n_549),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_642),
.B(n_631),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_L g841 ( 
.A(n_649),
.B(n_551),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_654),
.B(n_515),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_684),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_695),
.A2(n_579),
.B(n_543),
.Y(n_844)
);

OAI21x1_ASAP7_75t_L g845 ( 
.A1(n_702),
.A2(n_566),
.B(n_560),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_679),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_714),
.Y(n_847)
);

AOI21x1_ASAP7_75t_L g848 ( 
.A1(n_661),
.A2(n_566),
.B(n_630),
.Y(n_848)
);

O2A1O1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_797),
.A2(n_535),
.B(n_633),
.C(n_539),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_658),
.B(n_519),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_655),
.B(n_539),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_770),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_732),
.A2(n_543),
.B(n_527),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_684),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_681),
.A2(n_610),
.B(n_159),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_683),
.B(n_610),
.Y(n_856)
);

AOI21xp33_ASAP7_75t_L g857 ( 
.A1(n_741),
.A2(n_11),
.B(n_12),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_785),
.B(n_11),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_687),
.B(n_610),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_699),
.B(n_700),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_643),
.A2(n_610),
.B(n_20),
.C(n_21),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_645),
.A2(n_17),
.B(n_26),
.C(n_27),
.Y(n_862)
);

CKINVDCx10_ASAP7_75t_R g863 ( 
.A(n_791),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_741),
.A2(n_28),
.B(n_30),
.C(n_36),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_775),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_708),
.B(n_37),
.Y(n_866)
);

AOI21x1_ASAP7_75t_L g867 ( 
.A1(n_697),
.A2(n_72),
.B(n_143),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_649),
.B(n_62),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_679),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_720),
.B(n_723),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_725),
.A2(n_56),
.B1(n_140),
.B2(n_137),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_706),
.B(n_37),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_737),
.A2(n_102),
.B(n_98),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_649),
.B(n_95),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_728),
.B(n_730),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_772),
.A2(n_89),
.B(n_80),
.Y(n_876)
);

INVx6_ASAP7_75t_L g877 ( 
.A(n_657),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_R g878 ( 
.A(n_690),
.B(n_38),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_774),
.A2(n_698),
.B(n_794),
.Y(n_879)
);

A2O1A1Ixp33_ASAP7_75t_L g880 ( 
.A1(n_750),
.A2(n_51),
.B(n_42),
.C(n_43),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_706),
.B(n_40),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_657),
.B(n_674),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_646),
.B(n_40),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_698),
.A2(n_789),
.B(n_787),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_671),
.A2(n_44),
.B(n_45),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_725),
.A2(n_754),
.B1(n_676),
.B2(n_682),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_754),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_783),
.B(n_778),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_703),
.Y(n_890)
);

OAI21xp33_ASAP7_75t_L g891 ( 
.A1(n_750),
.A2(n_777),
.B(n_773),
.Y(n_891)
);

NOR2x1_ASAP7_75t_L g892 ( 
.A(n_731),
.B(n_738),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_767),
.B(n_773),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_767),
.B(n_777),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_649),
.B(n_764),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_709),
.B(n_659),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_721),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_662),
.B(n_664),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_711),
.B(n_712),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_733),
.B(n_648),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_648),
.B(n_675),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_740),
.B(n_717),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_680),
.A2(n_715),
.B(n_722),
.C(n_707),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_696),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_649),
.B(n_764),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_711),
.B(n_712),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_721),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_717),
.B(n_771),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_739),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_736),
.A2(n_745),
.B(n_753),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_686),
.B(n_693),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_744),
.A2(n_752),
.B(n_751),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_748),
.A2(n_714),
.B1(n_746),
.B2(n_727),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_688),
.B(n_716),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_793),
.B(n_734),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_649),
.B(n_714),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_691),
.B(n_758),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_739),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_790),
.A2(n_652),
.B(n_713),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_788),
.A2(n_738),
.B(n_669),
.C(n_781),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_788),
.B(n_746),
.Y(n_921)
);

AOI21x1_ASAP7_75t_L g922 ( 
.A1(n_742),
.A2(n_763),
.B(n_757),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_742),
.A2(n_757),
.B(n_781),
.C(n_765),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_755),
.B(n_748),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_735),
.A2(n_762),
.B(n_765),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_747),
.A2(n_763),
.B(n_749),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_761),
.B(n_665),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_769),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_673),
.B(n_685),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_747),
.A2(n_749),
.B(n_756),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_724),
.Y(n_931)
);

AO21x1_ASAP7_75t_L g932 ( 
.A1(n_756),
.A2(n_759),
.B(n_692),
.Y(n_932)
);

INVx4_ASAP7_75t_L g933 ( 
.A(n_665),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_759),
.B(n_701),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_665),
.A2(n_705),
.B(n_719),
.Y(n_935)
);

NOR2x1_ASAP7_75t_R g936 ( 
.A(n_705),
.B(n_719),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_SL g937 ( 
.A(n_705),
.B(n_719),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_726),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_786),
.A2(n_768),
.B(n_498),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_663),
.B(n_647),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_684),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_666),
.A2(n_797),
.B(n_653),
.C(n_501),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_647),
.B(n_496),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_647),
.B(n_496),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_946)
);

OAI22xp5_ASAP7_75t_L g947 ( 
.A1(n_647),
.A2(n_667),
.B1(n_768),
.B2(n_651),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_663),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_L g950 ( 
.A(n_769),
.B(n_508),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_647),
.B(n_496),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_670),
.A2(n_666),
.B(n_784),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_647),
.B(n_704),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_647),
.B(n_496),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_768),
.B(n_795),
.Y(n_956)
);

CKINVDCx8_ASAP7_75t_R g957 ( 
.A(n_724),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_663),
.B(n_647),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_768),
.B(n_795),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_647),
.B(n_704),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_702),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_770),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_729),
.A2(n_681),
.B(n_661),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_647),
.B(n_496),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_966)
);

NAND2x1p5_ASAP7_75t_L g967 ( 
.A(n_732),
.B(n_768),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_768),
.A2(n_498),
.B(n_521),
.Y(n_968)
);

AOI21x1_ASAP7_75t_L g969 ( 
.A1(n_729),
.A2(n_681),
.B(n_661),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_768),
.B(n_795),
.Y(n_970)
);

AO31x2_ASAP7_75t_L g971 ( 
.A1(n_932),
.A2(n_813),
.A3(n_947),
.B(n_804),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_942),
.Y(n_972)
);

NOR2x1_ASAP7_75t_L g973 ( 
.A(n_805),
.B(n_944),
.Y(n_973)
);

AND3x4_ASAP7_75t_L g974 ( 
.A(n_950),
.B(n_938),
.C(n_807),
.Y(n_974)
);

OAI22x1_ASAP7_75t_L g975 ( 
.A1(n_799),
.A2(n_906),
.B1(n_899),
.B2(n_881),
.Y(n_975)
);

OA21x2_ASAP7_75t_L g976 ( 
.A1(n_953),
.A2(n_886),
.B(n_901),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_891),
.A2(n_894),
.B(n_893),
.C(n_906),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_954),
.B(n_960),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_954),
.B(n_960),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_899),
.A2(n_801),
.B(n_872),
.C(n_881),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_872),
.A2(n_943),
.B(n_920),
.C(n_900),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_811),
.A2(n_841),
.B(n_925),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_800),
.A2(n_878),
.B1(n_915),
.B2(n_940),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_941),
.A2(n_949),
.B(n_946),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_890),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_951),
.A2(n_966),
.B(n_961),
.Y(n_986)
);

AOI21x1_ASAP7_75t_SL g987 ( 
.A1(n_934),
.A2(n_921),
.B(n_908),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_945),
.B(n_952),
.Y(n_988)
);

BUFx10_ASAP7_75t_L g989 ( 
.A(n_800),
.Y(n_989)
);

BUFx8_ASAP7_75t_SL g990 ( 
.A(n_928),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_818),
.A2(n_849),
.B(n_885),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_816),
.A2(n_838),
.B(n_968),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_895),
.A2(n_905),
.B(n_879),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_889),
.A2(n_930),
.B(n_923),
.C(n_902),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_858),
.A2(n_882),
.B(n_821),
.C(n_924),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_948),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_955),
.B(n_965),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_933),
.B(n_935),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_958),
.B(n_829),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_895),
.A2(n_905),
.B(n_970),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_956),
.A2(n_970),
.B(n_959),
.Y(n_1001)
);

AOI221xp5_ASAP7_75t_L g1002 ( 
.A1(n_857),
.A2(n_888),
.B1(n_878),
.B2(n_858),
.C(n_812),
.Y(n_1002)
);

NAND2x1_ASAP7_75t_SL g1003 ( 
.A(n_892),
.B(n_933),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_840),
.B(n_831),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_817),
.B(n_860),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_948),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_870),
.B(n_875),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_812),
.B(n_824),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_956),
.A2(n_959),
.B(n_917),
.Y(n_1009)
);

INVx4_ASAP7_75t_L g1010 ( 
.A(n_803),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_904),
.B(n_896),
.Y(n_1011)
);

OAI22x1_ASAP7_75t_L g1012 ( 
.A1(n_854),
.A2(n_927),
.B1(n_931),
.B2(n_924),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_918),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_910),
.A2(n_912),
.B(n_967),
.Y(n_1014)
);

AOI21x1_ASAP7_75t_L g1015 ( 
.A1(n_964),
.A2(n_969),
.B(n_825),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_916),
.A2(n_898),
.B(n_911),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_842),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_815),
.A2(n_913),
.B(n_810),
.Y(n_1018)
);

INVx5_ASAP7_75t_L g1019 ( 
.A(n_803),
.Y(n_1019)
);

AND2x4_ASAP7_75t_L g1020 ( 
.A(n_904),
.B(n_826),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_914),
.A2(n_820),
.B(n_827),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_819),
.A2(n_822),
.B(n_919),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_L g1023 ( 
.A(n_884),
.B(n_864),
.C(n_880),
.Y(n_1023)
);

AOI21x1_ASAP7_75t_SL g1024 ( 
.A1(n_866),
.A2(n_856),
.B(n_859),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_815),
.A2(n_887),
.B(n_824),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_806),
.B(n_843),
.Y(n_1026)
);

OAI21x1_ASAP7_75t_L g1027 ( 
.A1(n_814),
.A2(n_828),
.B(n_830),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_834),
.A2(n_835),
.B(n_833),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_939),
.A2(n_903),
.B(n_837),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_851),
.Y(n_1030)
);

INVx5_ASAP7_75t_L g1031 ( 
.A(n_803),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_869),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_832),
.A2(n_868),
.B(n_874),
.Y(n_1033)
);

A2O1A1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_850),
.A2(n_873),
.B(n_963),
.C(n_852),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_868),
.A2(n_874),
.B(n_825),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_823),
.B(n_962),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_927),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_922),
.A2(n_926),
.B(n_839),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_847),
.Y(n_1039)
);

AO31x2_ASAP7_75t_L g1040 ( 
.A1(n_871),
.A2(n_850),
.A3(n_876),
.B(n_865),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_962),
.B(n_823),
.Y(n_1041)
);

AO31x2_ASAP7_75t_L g1042 ( 
.A1(n_883),
.A2(n_897),
.A3(n_907),
.B(n_909),
.Y(n_1042)
);

O2A1O1Ixp5_ASAP7_75t_L g1043 ( 
.A1(n_808),
.A2(n_929),
.B(n_867),
.C(n_855),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_836),
.A2(n_844),
.B(n_853),
.Y(n_1044)
);

INVx1_ASAP7_75t_SL g1045 ( 
.A(n_877),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_877),
.A2(n_847),
.B1(n_843),
.B2(n_862),
.Y(n_1046)
);

AOI21x1_ASAP7_75t_L g1047 ( 
.A1(n_861),
.A2(n_877),
.B(n_937),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_957),
.Y(n_1048)
);

INVx2_ASAP7_75t_SL g1049 ( 
.A(n_863),
.Y(n_1049)
);

AOI21x1_ASAP7_75t_L g1050 ( 
.A1(n_936),
.A2(n_905),
.B(n_895),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_809),
.B(n_944),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_944),
.B(n_945),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_803),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_895),
.A2(n_905),
.B(n_885),
.Y(n_1054)
);

AOI221xp5_ASAP7_75t_L g1055 ( 
.A1(n_799),
.A2(n_710),
.B1(n_335),
.B2(n_906),
.C(n_899),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_799),
.A2(n_891),
.B(n_894),
.C(n_893),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_890),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_893),
.B(n_894),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_893),
.B(n_894),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_799),
.A2(n_943),
.B(n_905),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_893),
.B(n_894),
.Y(n_1061)
);

AOI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_799),
.A2(n_891),
.B1(n_906),
.B2(n_899),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_799),
.B(n_891),
.C(n_899),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_845),
.A2(n_802),
.B(n_848),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_893),
.B(n_894),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_890),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_935),
.B(n_684),
.Y(n_1067)
);

O2A1O1Ixp5_ASAP7_75t_L g1068 ( 
.A1(n_893),
.A2(n_894),
.B(n_906),
.C(n_899),
.Y(n_1068)
);

O2A1O1Ixp5_ASAP7_75t_L g1069 ( 
.A1(n_893),
.A2(n_894),
.B(n_906),
.C(n_899),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_890),
.Y(n_1070)
);

AO31x2_ASAP7_75t_L g1071 ( 
.A1(n_932),
.A2(n_813),
.A3(n_947),
.B(n_804),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_846),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_811),
.A2(n_768),
.B(n_841),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_845),
.A2(n_802),
.B(n_848),
.Y(n_1074)
);

OA22x2_ASAP7_75t_L g1075 ( 
.A1(n_886),
.A2(n_489),
.B1(n_891),
.B2(n_514),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_863),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_890),
.Y(n_1077)
);

AOI221x1_ASAP7_75t_L g1078 ( 
.A1(n_891),
.A2(n_893),
.B1(n_894),
.B2(n_881),
.C(n_872),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_846),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_846),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_956),
.A2(n_970),
.B(n_959),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_846),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_944),
.B(n_945),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_803),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_846),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_845),
.A2(n_802),
.B(n_848),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_SL g1087 ( 
.A1(n_956),
.A2(n_970),
.B(n_959),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_954),
.B(n_960),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_948),
.Y(n_1089)
);

NAND2xp33_ASAP7_75t_SL g1090 ( 
.A(n_893),
.B(n_894),
.Y(n_1090)
);

INVx5_ASAP7_75t_L g1091 ( 
.A(n_803),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_811),
.A2(n_768),
.B(n_841),
.Y(n_1092)
);

AOI21x1_ASAP7_75t_L g1093 ( 
.A1(n_895),
.A2(n_905),
.B(n_885),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_846),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_811),
.A2(n_768),
.B(n_841),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_845),
.A2(n_802),
.B(n_848),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_845),
.A2(n_802),
.B(n_848),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_799),
.A2(n_894),
.B1(n_893),
.B2(n_891),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_811),
.A2(n_768),
.B(n_841),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_799),
.A2(n_891),
.B(n_894),
.C(n_893),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_944),
.B(n_945),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_799),
.A2(n_891),
.B1(n_906),
.B2(n_899),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_944),
.B(n_945),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_890),
.Y(n_1104)
);

INVx6_ASAP7_75t_L g1105 ( 
.A(n_942),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_845),
.A2(n_802),
.B(n_848),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_899),
.B(n_906),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_890),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_899),
.B(n_906),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_899),
.B(n_906),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_811),
.A2(n_768),
.B(n_841),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_893),
.B(n_894),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_811),
.A2(n_768),
.B(n_841),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_893),
.B(n_894),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_1042),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_990),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_978),
.B(n_979),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_1105),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_985),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_978),
.B(n_979),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_1055),
.B(n_1004),
.Y(n_1122)
);

OA21x2_ASAP7_75t_L g1123 ( 
.A1(n_1018),
.A2(n_1025),
.B(n_1060),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1013),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_980),
.A2(n_1069),
.B(n_1068),
.C(n_1062),
.Y(n_1125)
);

OA21x2_ASAP7_75t_L g1126 ( 
.A1(n_1018),
.A2(n_1025),
.B(n_1060),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1105),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_999),
.B(n_1004),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1061),
.B(n_1065),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_972),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1102),
.A2(n_1114),
.B1(n_1112),
.B2(n_977),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1112),
.B(n_1114),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1088),
.B(n_988),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1089),
.Y(n_1136)
);

AND2x6_ASAP7_75t_L g1137 ( 
.A(n_1008),
.B(n_1039),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1057),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1010),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1020),
.B(n_983),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_996),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_988),
.B(n_997),
.Y(n_1142)
);

BUFx12f_ASAP7_75t_L g1143 ( 
.A(n_1076),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_997),
.B(n_1107),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1006),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1109),
.B(n_1110),
.Y(n_1146)
);

OA21x2_ASAP7_75t_L g1147 ( 
.A1(n_1064),
.A2(n_1106),
.B(n_1074),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1052),
.B(n_1083),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1020),
.B(n_1005),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_1051),
.B(n_1101),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1048),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_1039),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1075),
.A2(n_975),
.B1(n_1063),
.B2(n_1002),
.Y(n_1153)
);

O2A1O1Ixp5_ASAP7_75t_L g1154 ( 
.A1(n_1098),
.A2(n_1029),
.B(n_1090),
.C(n_981),
.Y(n_1154)
);

CKINVDCx16_ASAP7_75t_R g1155 ( 
.A(n_1049),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1005),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1103),
.B(n_1007),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_1003),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_1039),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_1019),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1007),
.B(n_973),
.Y(n_1161)
);

BUFx4_ASAP7_75t_SL g1162 ( 
.A(n_1067),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1063),
.B(n_1098),
.Y(n_1163)
);

CKINVDCx11_ASAP7_75t_R g1164 ( 
.A(n_989),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_989),
.B(n_1011),
.Y(n_1165)
);

BUFx12f_ASAP7_75t_L g1166 ( 
.A(n_1067),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1056),
.B(n_1100),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1072),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1086),
.A2(n_1097),
.B(n_1096),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1017),
.B(n_1030),
.Y(n_1170)
);

NAND2x1_ASAP7_75t_L g1171 ( 
.A(n_1010),
.B(n_998),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1026),
.B(n_1045),
.Y(n_1172)
);

OAI21xp33_ASAP7_75t_L g1173 ( 
.A1(n_1023),
.A2(n_995),
.B(n_994),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1023),
.A2(n_976),
.B1(n_1016),
.B2(n_974),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1079),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1066),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_1012),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1037),
.B(n_1045),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1080),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1070),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1078),
.B(n_1009),
.Y(n_1181)
);

INVx3_ASAP7_75t_SL g1182 ( 
.A(n_1067),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1082),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1077),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1034),
.B(n_1001),
.C(n_1000),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1085),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1104),
.B(n_1108),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1094),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_976),
.B(n_1087),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1046),
.A2(n_998),
.B1(n_1032),
.B2(n_1036),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1036),
.Y(n_1191)
);

INVx3_ASAP7_75t_SL g1192 ( 
.A(n_1019),
.Y(n_1192)
);

OR2x6_ASAP7_75t_L g1193 ( 
.A(n_1081),
.B(n_1046),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1041),
.B(n_1053),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1041),
.B(n_1050),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1031),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1014),
.A2(n_982),
.B(n_1113),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1021),
.B(n_971),
.Y(n_1198)
);

OR2x6_ASAP7_75t_SL g1199 ( 
.A(n_987),
.B(n_1024),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_971),
.B(n_1071),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_1084),
.Y(n_1201)
);

NOR2xp67_ASAP7_75t_L g1202 ( 
.A(n_1031),
.B(n_1091),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1073),
.A2(n_1111),
.B(n_1092),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_1033),
.A2(n_1035),
.B(n_993),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1071),
.B(n_1040),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1091),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1040),
.Y(n_1207)
);

CKINVDCx8_ASAP7_75t_R g1208 ( 
.A(n_1047),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_991),
.B(n_1028),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1015),
.B(n_1044),
.Y(n_1210)
);

AND2x6_ASAP7_75t_L g1211 ( 
.A(n_1043),
.B(n_1093),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1099),
.B(n_1095),
.Y(n_1212)
);

OA21x2_ASAP7_75t_L g1213 ( 
.A1(n_992),
.A2(n_1027),
.B(n_1054),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_984),
.A2(n_986),
.B(n_1022),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1038),
.B(n_1058),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1039),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1107),
.B(n_1109),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_999),
.B(n_958),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_990),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1220)
);

INVx1_ASAP7_75t_SL g1221 ( 
.A(n_999),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1004),
.B(n_1020),
.Y(n_1222)
);

BUFx6f_ASAP7_75t_L g1223 ( 
.A(n_1039),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_985),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_985),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1014),
.A2(n_768),
.B(n_994),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1055),
.A2(n_799),
.B1(n_906),
.B2(n_899),
.Y(n_1227)
);

AO31x2_ASAP7_75t_L g1228 ( 
.A1(n_980),
.A2(n_981),
.A3(n_1078),
.B(n_994),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_985),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1067),
.B(n_935),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_990),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1039),
.Y(n_1234)
);

BUFx2_ASAP7_75t_L g1235 ( 
.A(n_990),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_990),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_990),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1004),
.B(n_1020),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1004),
.B(n_1020),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_985),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_999),
.B(n_958),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1014),
.A2(n_768),
.B(n_994),
.Y(n_1243)
);

AND2x2_ASAP7_75t_SL g1244 ( 
.A(n_1002),
.B(n_899),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_996),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_978),
.B(n_979),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_980),
.A2(n_799),
.B(n_977),
.C(n_894),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1010),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1088),
.A2(n_931),
.B1(n_799),
.B2(n_906),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1250)
);

BUFx6f_ASAP7_75t_L g1251 ( 
.A(n_1039),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_980),
.A2(n_891),
.B(n_799),
.C(n_899),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_990),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1058),
.B(n_1059),
.Y(n_1255)
);

INVx5_ASAP7_75t_L g1256 ( 
.A(n_1039),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1115),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1187),
.Y(n_1258)
);

CKINVDCx20_ASAP7_75t_R g1259 ( 
.A(n_1155),
.Y(n_1259)
);

CKINVDCx8_ASAP7_75t_R g1260 ( 
.A(n_1116),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1227),
.A2(n_1253),
.B(n_1244),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1142),
.B(n_1157),
.Y(n_1262)
);

BUFx8_ASAP7_75t_L g1263 ( 
.A(n_1233),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1249),
.A2(n_1255),
.B1(n_1229),
.B2(n_1127),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1245),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1150),
.B(n_1135),
.Y(n_1266)
);

BUFx10_ASAP7_75t_L g1267 ( 
.A(n_1254),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1187),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1153),
.A2(n_1122),
.B1(n_1193),
.B2(n_1173),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1203),
.A2(n_1212),
.B(n_1154),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1119),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1208),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1245),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1124),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1203),
.A2(n_1197),
.B(n_1226),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1215),
.Y(n_1276)
);

AO21x1_ASAP7_75t_L g1277 ( 
.A1(n_1247),
.A2(n_1174),
.B(n_1133),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1193),
.A2(n_1217),
.B1(n_1163),
.B2(n_1140),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1191),
.Y(n_1279)
);

OAI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1135),
.A2(n_1148),
.B1(n_1134),
.B2(n_1255),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_SL g1281 ( 
.A(n_1219),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1193),
.A2(n_1177),
.B1(n_1133),
.B2(n_1161),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1145),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1166),
.Y(n_1284)
);

AND2x2_ASAP7_75t_L g1285 ( 
.A(n_1142),
.B(n_1121),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1199),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1138),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1146),
.A2(n_1218),
.B1(n_1242),
.B2(n_1130),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1146),
.A2(n_1221),
.B1(n_1167),
.B2(n_1172),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1176),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1121),
.A2(n_1230),
.B1(n_1220),
.B2(n_1229),
.Y(n_1291)
);

BUFx2_ASAP7_75t_R g1292 ( 
.A(n_1238),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1180),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1184),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1197),
.A2(n_1214),
.B(n_1243),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1127),
.A2(n_1131),
.B1(n_1250),
.B2(n_1236),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1171),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1123),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1129),
.A2(n_1131),
.B1(n_1250),
.B2(n_1236),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1129),
.B(n_1220),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1224),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1123),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1126),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1230),
.A2(n_1252),
.B1(n_1117),
.B2(n_1120),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1212),
.A2(n_1154),
.B(n_1125),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1225),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1231),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1252),
.A2(n_1246),
.B1(n_1221),
.B2(n_1144),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1144),
.B(n_1194),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1167),
.A2(n_1156),
.B1(n_1165),
.B2(n_1182),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1241),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1178),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1170),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1118),
.Y(n_1314)
);

AO21x1_ASAP7_75t_SL g1315 ( 
.A1(n_1200),
.A2(n_1189),
.B(n_1181),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1170),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1126),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1132),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1149),
.A2(n_1207),
.B1(n_1174),
.B2(n_1222),
.Y(n_1319)
);

CKINVDCx9p33_ASAP7_75t_R g1320 ( 
.A(n_1235),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1222),
.B(n_1239),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_SL g1322 ( 
.A1(n_1247),
.A2(n_1204),
.B(n_1190),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1141),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1239),
.A2(n_1240),
.B1(n_1195),
.B2(n_1185),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1151),
.Y(n_1325)
);

INVx4_ASAP7_75t_SL g1326 ( 
.A(n_1137),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1240),
.A2(n_1185),
.B1(n_1205),
.B2(n_1232),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1232),
.A2(n_1164),
.B1(n_1211),
.B2(n_1189),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1198),
.A2(n_1200),
.B(n_1209),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1228),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1211),
.A2(n_1210),
.B(n_1232),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1143),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1136),
.B(n_1175),
.Y(n_1333)
);

OAI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1158),
.A2(n_1237),
.B1(n_1192),
.B2(n_1128),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1168),
.Y(n_1335)
);

INVxp67_ASAP7_75t_L g1336 ( 
.A(n_1201),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1179),
.A2(n_1188),
.B1(n_1186),
.B2(n_1183),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1211),
.A2(n_1213),
.B(n_1228),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1228),
.Y(n_1339)
);

INVx3_ASAP7_75t_L g1340 ( 
.A(n_1137),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1160),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1137),
.B(n_1139),
.Y(n_1342)
);

OA21x2_ASAP7_75t_L g1343 ( 
.A1(n_1213),
.A2(n_1147),
.B(n_1169),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1196),
.A2(n_1248),
.B1(n_1251),
.B2(n_1152),
.Y(n_1344)
);

BUFx4f_ASAP7_75t_SL g1345 ( 
.A(n_1206),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1248),
.A2(n_1202),
.B(n_1162),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1152),
.B(n_1223),
.Y(n_1347)
);

AO21x2_ASAP7_75t_L g1348 ( 
.A1(n_1162),
.A2(n_1159),
.B(n_1256),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1216),
.B(n_1234),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_1234),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1115),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1244),
.A2(n_799),
.B1(n_1075),
.B2(n_891),
.Y(n_1352)
);

NAND2x1p5_ASAP7_75t_L g1353 ( 
.A(n_1190),
.B(n_1123),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1187),
.Y(n_1354)
);

NAND2x1p5_ASAP7_75t_L g1355 ( 
.A(n_1190),
.B(n_1123),
.Y(n_1355)
);

BUFx8_ASAP7_75t_SL g1356 ( 
.A(n_1143),
.Y(n_1356)
);

AO21x2_ASAP7_75t_L g1357 ( 
.A1(n_1197),
.A2(n_1214),
.B(n_1203),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1187),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1187),
.Y(n_1359)
);

AO21x2_ASAP7_75t_L g1360 ( 
.A1(n_1197),
.A2(n_1214),
.B(n_1203),
.Y(n_1360)
);

AOI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1227),
.A2(n_899),
.B1(n_906),
.B2(n_799),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1221),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1145),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_SL g1364 ( 
.A1(n_1244),
.A2(n_906),
.B1(n_899),
.B2(n_799),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1244),
.B(n_1142),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1257),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1265),
.Y(n_1367)
);

INVx5_ASAP7_75t_SL g1368 ( 
.A(n_1320),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1265),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1273),
.Y(n_1370)
);

NAND3xp33_ASAP7_75t_L g1371 ( 
.A(n_1364),
.B(n_1361),
.C(n_1352),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1365),
.B(n_1309),
.Y(n_1372)
);

HB1xp67_ASAP7_75t_L g1373 ( 
.A(n_1273),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1340),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1365),
.B(n_1309),
.Y(n_1375)
);

AO21x1_ASAP7_75t_SL g1376 ( 
.A1(n_1330),
.A2(n_1261),
.B(n_1328),
.Y(n_1376)
);

CKINVDCx14_ASAP7_75t_R g1377 ( 
.A(n_1259),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1340),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1322),
.A2(n_1275),
.B(n_1277),
.Y(n_1379)
);

INVx3_ASAP7_75t_L g1380 ( 
.A(n_1329),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1262),
.B(n_1266),
.Y(n_1381)
);

NAND2x1p5_ASAP7_75t_L g1382 ( 
.A(n_1305),
.B(n_1329),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1270),
.A2(n_1360),
.B(n_1357),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1298),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1283),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1283),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1331),
.B(n_1351),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1322),
.A2(n_1277),
.B(n_1295),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1262),
.B(n_1285),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1302),
.Y(n_1390)
);

INVxp67_ASAP7_75t_L g1391 ( 
.A(n_1363),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1303),
.Y(n_1392)
);

OAI21xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1269),
.A2(n_1300),
.B(n_1299),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1285),
.B(n_1304),
.Y(n_1394)
);

AND2x6_ASAP7_75t_L g1395 ( 
.A(n_1340),
.B(n_1297),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1362),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1317),
.Y(n_1397)
);

OR2x6_ASAP7_75t_L g1398 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1348),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1276),
.B(n_1329),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1346),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1276),
.B(n_1315),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1341),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1315),
.B(n_1278),
.Y(n_1404)
);

INVx3_ASAP7_75t_L g1405 ( 
.A(n_1338),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1312),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1339),
.B(n_1353),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1343),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1294),
.Y(n_1410)
);

OR2x6_ASAP7_75t_L g1411 ( 
.A(n_1353),
.B(n_1355),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1279),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1264),
.A2(n_1280),
.B(n_1324),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1301),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1305),
.B(n_1338),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1271),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1274),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1290),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1306),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1307),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1311),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1313),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1316),
.B(n_1291),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_1258),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1268),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_SL g1426 ( 
.A1(n_1282),
.A2(n_1327),
.B(n_1296),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1354),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1319),
.A2(n_1359),
.B(n_1358),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1409),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1402),
.B(n_1382),
.Y(n_1430)
);

INVxp67_ASAP7_75t_L g1431 ( 
.A(n_1367),
.Y(n_1431)
);

BUFx2_ASAP7_75t_SL g1432 ( 
.A(n_1399),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1400),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1400),
.B(n_1286),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1402),
.B(n_1286),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1401),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1382),
.B(n_1384),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1390),
.B(n_1335),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1392),
.B(n_1288),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1394),
.B(n_1308),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1397),
.B(n_1289),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1371),
.A2(n_1413),
.B(n_1310),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1380),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1398),
.B(n_1326),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1388),
.B(n_1349),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1380),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1395),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1405),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1383),
.A2(n_1348),
.B(n_1272),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1370),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1415),
.B(n_1272),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1388),
.B(n_1347),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1388),
.B(n_1379),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1398),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1423),
.B(n_1272),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1379),
.B(n_1347),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1366),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1415),
.B(n_1398),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1379),
.B(n_1349),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1373),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1395),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1398),
.B(n_1326),
.Y(n_1462)
);

NAND3xp33_ASAP7_75t_L g1463 ( 
.A(n_1442),
.B(n_1371),
.C(n_1393),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1442),
.A2(n_1440),
.B(n_1377),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1430),
.B(n_1445),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1440),
.B(n_1393),
.C(n_1404),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1455),
.A2(n_1391),
.B1(n_1426),
.B2(n_1334),
.C(n_1385),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1455),
.A2(n_1426),
.B1(n_1386),
.B2(n_1406),
.C(n_1381),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1431),
.B(n_1372),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1431),
.B(n_1372),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1450),
.A2(n_1396),
.B1(n_1375),
.B2(n_1336),
.C(n_1389),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1450),
.B(n_1369),
.Y(n_1472)
);

NAND2xp33_ASAP7_75t_L g1473 ( 
.A(n_1454),
.B(n_1395),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1460),
.B(n_1403),
.Y(n_1474)
);

NAND3xp33_ASAP7_75t_L g1475 ( 
.A(n_1449),
.B(n_1424),
.C(n_1428),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1445),
.B(n_1398),
.Y(n_1476)
);

NOR3xp33_ASAP7_75t_L g1477 ( 
.A(n_1449),
.B(n_1342),
.C(n_1284),
.Y(n_1477)
);

NAND3xp33_ASAP7_75t_L g1478 ( 
.A(n_1453),
.B(n_1428),
.C(n_1427),
.Y(n_1478)
);

AOI21xp33_ASAP7_75t_L g1479 ( 
.A1(n_1451),
.A2(n_1441),
.B(n_1434),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1445),
.B(n_1452),
.Y(n_1480)
);

OAI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1460),
.A2(n_1284),
.B1(n_1321),
.B2(n_1318),
.C(n_1344),
.Y(n_1481)
);

NAND3xp33_ASAP7_75t_L g1482 ( 
.A(n_1453),
.B(n_1428),
.C(n_1422),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1439),
.B(n_1417),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1439),
.B(n_1417),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1435),
.B(n_1325),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1439),
.A2(n_1376),
.B1(n_1462),
.B2(n_1444),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1444),
.A2(n_1401),
.B(n_1387),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1441),
.B(n_1418),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_SL g1489 ( 
.A(n_1447),
.B(n_1401),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1441),
.B(n_1418),
.Y(n_1490)
);

AND2x2_ASAP7_75t_SL g1491 ( 
.A(n_1454),
.B(n_1428),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1447),
.A2(n_1368),
.B1(n_1259),
.B2(n_1350),
.Y(n_1492)
);

NAND4xp25_ASAP7_75t_L g1493 ( 
.A(n_1451),
.B(n_1333),
.C(n_1420),
.D(n_1419),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1447),
.A2(n_1368),
.B1(n_1350),
.B2(n_1425),
.Y(n_1494)
);

OAI21xp33_ASAP7_75t_L g1495 ( 
.A1(n_1453),
.A2(n_1387),
.B(n_1427),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1435),
.B(n_1421),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1456),
.B(n_1411),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1435),
.B(n_1421),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1434),
.B(n_1416),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1447),
.A2(n_1368),
.B1(n_1425),
.B2(n_1422),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1447),
.A2(n_1368),
.B1(n_1374),
.B2(n_1378),
.Y(n_1501)
);

NAND3xp33_ASAP7_75t_L g1502 ( 
.A(n_1451),
.B(n_1412),
.C(n_1323),
.Y(n_1502)
);

OAI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1434),
.A2(n_1416),
.B(n_1420),
.Y(n_1503)
);

OAI221xp5_ASAP7_75t_SL g1504 ( 
.A1(n_1458),
.A2(n_1411),
.B1(n_1407),
.B2(n_1399),
.C(n_1419),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1456),
.B(n_1411),
.Y(n_1505)
);

AOI221xp5_ASAP7_75t_L g1506 ( 
.A1(n_1437),
.A2(n_1337),
.B1(n_1387),
.B2(n_1410),
.C(n_1414),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1438),
.B(n_1408),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1456),
.B(n_1407),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1438),
.B(n_1408),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1446),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1499),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1480),
.B(n_1433),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1491),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1488),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1490),
.Y(n_1516)
);

AND2x4_ASAP7_75t_L g1517 ( 
.A(n_1489),
.B(n_1454),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1483),
.Y(n_1518)
);

NAND2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1491),
.B(n_1461),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1484),
.B(n_1433),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1465),
.B(n_1446),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1496),
.B(n_1458),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1507),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1498),
.B(n_1458),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1508),
.B(n_1437),
.Y(n_1525)
);

INVx3_ASAP7_75t_L g1526 ( 
.A(n_1497),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1474),
.B(n_1437),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1497),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1503),
.B(n_1459),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1509),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1476),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1472),
.B(n_1459),
.Y(n_1533)
);

INVx3_ASAP7_75t_L g1534 ( 
.A(n_1505),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1469),
.B(n_1459),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1470),
.B(n_1457),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1505),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1479),
.B(n_1443),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1495),
.B(n_1443),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1487),
.B(n_1443),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.B(n_1448),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1478),
.B(n_1429),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1482),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1517),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1539),
.B(n_1468),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1543),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1539),
.B(n_1506),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1543),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1512),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1531),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1512),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1517),
.B(n_1454),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1510),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1510),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1510),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1544),
.B(n_1529),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1526),
.B(n_1454),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1513),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1544),
.B(n_1475),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1466),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1519),
.Y(n_1566)
);

OAI22xp5_ASAP7_75t_L g1567 ( 
.A1(n_1519),
.A2(n_1463),
.B1(n_1464),
.B2(n_1486),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1534),
.B(n_1477),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.B(n_1493),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1513),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1533),
.B(n_1504),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1536),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1517),
.B(n_1444),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1513),
.Y(n_1574)
);

NOR2xp67_ASAP7_75t_L g1575 ( 
.A(n_1514),
.B(n_1485),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1521),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1527),
.B(n_1281),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1511),
.B(n_1467),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1536),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1534),
.B(n_1436),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1533),
.B(n_1429),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1535),
.B(n_1429),
.Y(n_1582)
);

INVx1_ASAP7_75t_SL g1583 ( 
.A(n_1527),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1551),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1546),
.A2(n_1514),
.B(n_1471),
.C(n_1540),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1569),
.B(n_1522),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1562),
.B(n_1515),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1569),
.B(n_1522),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1548),
.B(n_1281),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1562),
.B(n_1515),
.Y(n_1591)
);

NAND2x2_ASAP7_75t_L g1592 ( 
.A(n_1578),
.B(n_1528),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1584),
.B(n_1517),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1565),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1516),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1547),
.B(n_1516),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1549),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1549),
.Y(n_1598)
);

NOR2x1_ASAP7_75t_L g1599 ( 
.A(n_1564),
.B(n_1492),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1537),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1554),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1566),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1555),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1577),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1545),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1573),
.B(n_1537),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1564),
.Y(n_1608)
);

AOI221xp5_ASAP7_75t_L g1609 ( 
.A1(n_1567),
.A2(n_1481),
.B1(n_1518),
.B2(n_1530),
.C(n_1523),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1517),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1559),
.B(n_1524),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1559),
.B(n_1524),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1555),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1558),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1545),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1558),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1550),
.B(n_1518),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_L g1618 ( 
.A(n_1571),
.B(n_1519),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1550),
.B(n_1523),
.Y(n_1619)
);

AND2x4_ASAP7_75t_SL g1620 ( 
.A(n_1556),
.B(n_1267),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1563),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1571),
.A2(n_1473),
.B(n_1494),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1545),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1563),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1570),
.Y(n_1625)
);

NAND2x1p5_ASAP7_75t_L g1626 ( 
.A(n_1566),
.B(n_1461),
.Y(n_1626)
);

AOI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1575),
.A2(n_1538),
.B(n_1520),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1593),
.B(n_1553),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1593),
.Y(n_1629)
);

AND3x1_ASAP7_75t_L g1630 ( 
.A(n_1599),
.B(n_1568),
.C(n_1557),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1608),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1627),
.B(n_1553),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1608),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1601),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1586),
.A2(n_1519),
.B1(n_1583),
.B2(n_1553),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1552),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1603),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1610),
.B(n_1568),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1556),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1618),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1587),
.B(n_1552),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1602),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1557),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1615),
.B(n_1560),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1585),
.Y(n_1645)
);

AO21x2_ASAP7_75t_L g1646 ( 
.A1(n_1585),
.A2(n_1579),
.B(n_1572),
.Y(n_1646)
);

OAI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1592),
.A2(n_1622),
.B1(n_1609),
.B2(n_1605),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1597),
.B(n_1572),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1623),
.B(n_1560),
.Y(n_1649)
);

AOI222xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1598),
.A2(n_1579),
.B1(n_1570),
.B2(n_1576),
.C1(n_1574),
.C2(n_1530),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1589),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1588),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1609),
.B(n_1574),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1561),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1626),
.B(n_1561),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1611),
.B(n_1576),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1590),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1588),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1591),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1600),
.B(n_1580),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1604),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1591),
.Y(n_1662)
);

CKINVDCx16_ASAP7_75t_R g1663 ( 
.A(n_1607),
.Y(n_1663)
);

AOI21xp33_ASAP7_75t_SL g1664 ( 
.A1(n_1647),
.A2(n_1332),
.B(n_1612),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1663),
.B(n_1620),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1631),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1637),
.B(n_1622),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_SL g1668 ( 
.A1(n_1635),
.A2(n_1595),
.B1(n_1596),
.B2(n_1614),
.Y(n_1668)
);

AOI222xp33_ASAP7_75t_L g1669 ( 
.A1(n_1653),
.A2(n_1595),
.B1(n_1596),
.B2(n_1624),
.C1(n_1625),
.C2(n_1621),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1657),
.B(n_1356),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1630),
.A2(n_1619),
.B1(n_1617),
.B2(n_1616),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1651),
.B(n_1619),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1631),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1630),
.A2(n_1617),
.B1(n_1613),
.B2(n_1501),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1631),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1638),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1635),
.A2(n_1538),
.B(n_1540),
.C(n_1541),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1645),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1637),
.B(n_1645),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1651),
.B(n_1532),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1653),
.B(n_1535),
.Y(n_1681)
);

OAI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1640),
.A2(n_1542),
.A3(n_1541),
.B1(n_1580),
.B2(n_1534),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1657),
.A2(n_1376),
.B1(n_1432),
.B2(n_1500),
.Y(n_1683)
);

OAI322xp33_ASAP7_75t_L g1684 ( 
.A1(n_1633),
.A2(n_1581),
.A3(n_1582),
.B1(n_1520),
.B2(n_1525),
.C1(n_1528),
.C2(n_1542),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1633),
.Y(n_1685)
);

OAI31xp33_ASAP7_75t_L g1686 ( 
.A1(n_1640),
.A2(n_1541),
.A3(n_1538),
.B(n_1542),
.Y(n_1686)
);

AOI21xp33_ASAP7_75t_L g1687 ( 
.A1(n_1629),
.A2(n_1540),
.B(n_1263),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1629),
.B(n_1532),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

NOR3xp33_ASAP7_75t_SL g1690 ( 
.A(n_1679),
.B(n_1670),
.C(n_1678),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1685),
.B(n_1638),
.Y(n_1692)
);

NAND2x1p5_ASAP7_75t_L g1693 ( 
.A(n_1666),
.B(n_1673),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1676),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.B(n_1641),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1675),
.B(n_1689),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1665),
.B(n_1638),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1689),
.Y(n_1698)
);

NOR2x1_ASAP7_75t_L g1699 ( 
.A(n_1672),
.B(n_1646),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1659),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1674),
.B(n_1659),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1681),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1664),
.B(n_1660),
.Y(n_1703)
);

NOR2xp67_ASAP7_75t_L g1704 ( 
.A(n_1671),
.B(n_1632),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1680),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1687),
.B(n_1639),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1688),
.B(n_1639),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1684),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1682),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1690),
.A2(n_1686),
.B(n_1677),
.C(n_1632),
.Y(n_1710)
);

OAI21xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1704),
.A2(n_1699),
.B(n_1691),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1690),
.A2(n_1668),
.B1(n_1632),
.B2(n_1662),
.C(n_1652),
.Y(n_1712)
);

NOR3xp33_ASAP7_75t_L g1713 ( 
.A(n_1691),
.B(n_1636),
.C(n_1652),
.Y(n_1713)
);

NOR3xp33_ASAP7_75t_L g1714 ( 
.A(n_1700),
.B(n_1636),
.C(n_1658),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1708),
.A2(n_1683),
.B(n_1639),
.Y(n_1715)
);

AOI21xp33_ASAP7_75t_L g1716 ( 
.A1(n_1702),
.A2(n_1662),
.B(n_1658),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1701),
.A2(n_1683),
.B1(n_1646),
.B2(n_1642),
.C(n_1634),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1703),
.A2(n_1646),
.B(n_1648),
.Y(n_1718)
);

NAND4xp75_ASAP7_75t_L g1719 ( 
.A(n_1698),
.B(n_1628),
.C(n_1654),
.D(n_1655),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1709),
.A2(n_1646),
.B1(n_1634),
.B2(n_1642),
.C(n_1661),
.Y(n_1720)
);

OA21x2_ASAP7_75t_L g1721 ( 
.A1(n_1696),
.A2(n_1642),
.B(n_1634),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1715),
.B(n_1692),
.Y(n_1722)
);

OA22x2_ASAP7_75t_L g1723 ( 
.A1(n_1711),
.A2(n_1697),
.B1(n_1694),
.B2(n_1705),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1713),
.B(n_1693),
.Y(n_1724)
);

AND3x1_ASAP7_75t_L g1725 ( 
.A(n_1714),
.B(n_1694),
.C(n_1706),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_L g1726 ( 
.A(n_1720),
.B(n_1706),
.C(n_1695),
.Y(n_1726)
);

NAND3xp33_ASAP7_75t_L g1727 ( 
.A(n_1717),
.B(n_1650),
.C(n_1707),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1719),
.B(n_1693),
.Y(n_1728)
);

OAI211xp5_ASAP7_75t_SL g1729 ( 
.A1(n_1710),
.A2(n_1641),
.B(n_1661),
.C(n_1260),
.Y(n_1729)
);

NAND2xp33_ASAP7_75t_SL g1730 ( 
.A(n_1712),
.B(n_1332),
.Y(n_1730)
);

NOR2x1_ASAP7_75t_L g1731 ( 
.A(n_1721),
.B(n_1707),
.Y(n_1731)
);

NAND2x1p5_ASAP7_75t_L g1732 ( 
.A(n_1721),
.B(n_1318),
.Y(n_1732)
);

NOR2x1_ASAP7_75t_L g1733 ( 
.A(n_1718),
.B(n_1661),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1731),
.Y(n_1734)
);

OAI21xp5_ASAP7_75t_L g1735 ( 
.A1(n_1727),
.A2(n_1716),
.B(n_1628),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1725),
.A2(n_1628),
.B1(n_1648),
.B2(n_1649),
.C(n_1643),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1726),
.B(n_1660),
.Y(n_1737)
);

NOR4xp25_ASAP7_75t_L g1738 ( 
.A(n_1724),
.B(n_1641),
.C(n_1649),
.D(n_1644),
.Y(n_1738)
);

XNOR2xp5_ASAP7_75t_L g1739 ( 
.A(n_1723),
.B(n_1356),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1729),
.B(n_1314),
.C(n_1654),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1734),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1737),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1739),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_1735),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1738),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1736),
.Y(n_1746)
);

AO22x2_ASAP7_75t_L g1747 ( 
.A1(n_1745),
.A2(n_1728),
.B1(n_1722),
.B2(n_1740),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_1743),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1741),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1744),
.B(n_1730),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1744),
.A2(n_1733),
.B(n_1260),
.C(n_1732),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1749),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1748),
.B(n_1746),
.C(n_1742),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1747),
.B(n_1750),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1752),
.Y(n_1755)
);

OAI222xp33_ASAP7_75t_L g1756 ( 
.A1(n_1755),
.A2(n_1754),
.B1(n_1751),
.B2(n_1753),
.C1(n_1345),
.C2(n_1655),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_R g1757 ( 
.A(n_1756),
.B(n_1325),
.Y(n_1757)
);

AOI221x1_ASAP7_75t_L g1758 ( 
.A1(n_1756),
.A2(n_1654),
.B1(n_1655),
.B2(n_1643),
.C(n_1649),
.Y(n_1758)
);

BUFx2_ASAP7_75t_L g1759 ( 
.A(n_1757),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1758),
.B(n_1267),
.Y(n_1760)
);

XNOR2xp5_ASAP7_75t_L g1761 ( 
.A(n_1759),
.B(n_1314),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1760),
.Y(n_1762)
);

OR2x6_ASAP7_75t_L g1763 ( 
.A(n_1762),
.B(n_1267),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1763),
.A2(n_1761),
.B1(n_1281),
.B2(n_1263),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1644),
.B1(n_1643),
.B2(n_1660),
.C(n_1656),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1263),
.B(n_1292),
.C(n_1644),
.Y(n_1766)
);


endmodule