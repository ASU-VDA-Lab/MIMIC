module real_jpeg_32270_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_546, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_546;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_534;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_15;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_468;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_0),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_0),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_1),
.A2(n_277),
.B1(n_280),
.B2(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_1),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_1),
.A2(n_280),
.B1(n_336),
.B2(n_339),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_1),
.A2(n_280),
.B1(n_436),
.B2(n_438),
.Y(n_435)
);

OAI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_1),
.A2(n_280),
.B1(n_468),
.B2(n_470),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_3),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_5),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_5),
.Y(n_127)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_6),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_7),
.A2(n_108),
.B1(n_113),
.B2(n_114),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_7),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_7),
.A2(n_113),
.B1(n_186),
.B2(n_190),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_7),
.A2(n_113),
.B1(n_229),
.B2(n_232),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_7),
.A2(n_113),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_8),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_43),
.B1(n_98),
.B2(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_8),
.A2(n_43),
.B1(n_132),
.B2(n_135),
.Y(n_131)
);

AO22x1_ASAP7_75t_L g219 ( 
.A1(n_8),
.A2(n_43),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_8),
.B(n_25),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_SL g427 ( 
.A(n_8),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_8),
.B(n_119),
.Y(n_463)
);

OAI32xp33_ASAP7_75t_L g479 ( 
.A1(n_8),
.A2(n_480),
.A3(n_482),
.B1(n_483),
.B2(n_489),
.Y(n_479)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_9),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_9),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_11),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_12),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_13),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_13),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g139 ( 
.A1(n_13),
.A2(n_54),
.B1(n_140),
.B2(n_144),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_13),
.A2(n_54),
.B1(n_229),
.B2(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_13),
.A2(n_54),
.B1(n_215),
.B2(n_267),
.Y(n_266)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21x1_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_532),
.B(n_543),
.Y(n_17)
);

NOR2x1_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_292),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_199),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_170),
.Y(n_20)
);

AOI32xp33_ASAP7_75t_L g542 ( 
.A1(n_21),
.A2(n_170),
.A3(n_536),
.B1(n_537),
.B2(n_546),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_66),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_23),
.Y(n_533)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_23),
.B(n_66),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_49),
.Y(n_23)
);

NAND2x1_ASAP7_75t_SL g274 ( 
.A(n_24),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_39),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_51),
.Y(n_166)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_26),
.A2(n_49),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_26),
.B(n_164),
.Y(n_244)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2x1p5_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_27),
.B(n_276),
.Y(n_319)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_29),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_29),
.Y(n_360)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_31),
.Y(n_338)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_32),
.Y(n_136)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_33),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_34),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_34),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_39),
.B(n_58),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_39),
.B(n_244),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_43),
.B(n_44),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_42),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_42),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_45),
.Y(n_44)
);

AOI32xp33_ASAP7_75t_L g422 ( 
.A1(n_43),
.A2(n_423),
.A3(n_425),
.B1(n_426),
.B2(n_427),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_43),
.B(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_43),
.B(n_511),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_43),
.B(n_519),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_44),
.Y(n_365)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_50),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_57),
.Y(n_355)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_58),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_58),
.B(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_163),
.C(n_167),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_67),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_R g67 ( 
.A(n_68),
.B(n_105),
.C(n_115),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_68),
.A2(n_116),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_68),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_68),
.B(n_182),
.C(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_68),
.A2(n_176),
.B1(n_184),
.B2(n_205),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_68),
.B(n_376),
.C(n_378),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_68),
.A2(n_176),
.B1(n_376),
.B2(n_388),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_83),
.B(n_97),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_69),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_69),
.B(n_97),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_69),
.B(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_69),
.B(n_435),
.Y(n_448)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_84),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_70),
.Y(n_511)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_76),
.Y(n_469)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_76),
.Y(n_472)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_79),
.Y(n_313)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_83),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_83),
.B(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_83),
.B(n_97),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_83),
.B(n_435),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_122),
.B1(n_125),
.B2(n_128),
.Y(n_121)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_94),
.Y(n_437)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_101),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_101),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_101),
.Y(n_440)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_104),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_105),
.A2(n_106),
.B1(n_174),
.B2(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21x1_ASAP7_75t_SL g163 ( 
.A1(n_107),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_137),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_118),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_130),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_139),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_119),
.A2(n_137),
.B(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_119),
.B(n_335),
.Y(n_377)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_120),
.A2(n_131),
.B(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_150),
.B(n_157),
.Y(n_149)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_129),
.Y(n_231)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_131),
.B(n_149),
.Y(n_273)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_138),
.B(n_377),
.Y(n_376)
);

NAND2x1_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_148),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_141),
.Y(n_348)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_148),
.B(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_154),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_151),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_151),
.Y(n_425)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_153),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_157),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_167),
.B1(n_168),
.B2(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_163),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_179),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_166),
.B(n_275),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_167),
.B(n_306),
.C(n_318),
.Y(n_305)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2x1_ASAP7_75t_L g325 ( 
.A(n_169),
.B(n_318),
.Y(n_325)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_196),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_172),
.B(n_196),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.C(n_180),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_173),
.A2(n_178),
.B1(n_182),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_173),
.Y(n_255)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_178),
.A2(n_182),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_179),
.B(n_319),
.Y(n_378)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_254),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_193),
.B(n_194),
.Y(n_184)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_185),
.Y(n_248)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_194),
.B(n_334),
.Y(n_392)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2x1_ASAP7_75t_L g272 ( 
.A(n_195),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_252),
.B1(n_256),
.B2(n_288),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_201),
.B(n_253),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_201),
.B(n_253),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.C(n_245),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_202),
.A2(n_245),
.B1(n_246),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_206),
.B(n_290),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_225),
.B(n_242),
.Y(n_206)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_207),
.B(n_243),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_207),
.A2(n_226),
.B1(n_241),
.B2(n_304),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_207),
.B(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_207),
.A2(n_241),
.B1(n_422),
.B2(n_454),
.Y(n_453)
);

AO21x2_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_211),
.B(n_218),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_208),
.A2(n_265),
.B(n_311),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_210),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_211),
.A2(n_311),
.B(n_314),
.Y(n_310)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_212),
.B(n_219),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_212),
.B(n_467),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g506 ( 
.A(n_214),
.Y(n_506)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_215),
.Y(n_481)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_217),
.Y(n_269)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_217),
.Y(n_312)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g286 ( 
.A(n_225),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_241),
.Y(n_225)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_234),
.B(n_235),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_231),
.Y(n_233)
);

INVx5_ASAP7_75t_L g482 ( 
.A(n_231),
.Y(n_482)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_235),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_235),
.B(n_434),
.Y(n_461)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_242),
.A2(n_533),
.B(n_534),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_242),
.B(n_533),
.Y(n_543)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_249),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g284 ( 
.A(n_247),
.B(n_249),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_250),
.B(n_434),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_251),
.B(n_260),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_251),
.B(n_448),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_257),
.B(n_289),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_284),
.C(n_285),
.Y(n_257)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_258),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_270),
.C(n_274),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g300 ( 
.A(n_259),
.B(n_301),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_261),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

AND2x2_ASAP7_75t_SL g465 ( 
.A(n_262),
.B(n_466),
.Y(n_465)
);

BUFx4f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_265),
.B(n_504),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_266),
.B(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_271),
.A2(n_272),
.B1(n_274),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_273),
.Y(n_451)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx4_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_284),
.B(n_286),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2x1p5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_413),
.Y(n_293)
);

OAI21x1_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_366),
.B(n_407),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_321),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_305),
.B2(n_320),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_298),
.B(n_305),
.Y(n_406)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_299),
.B(n_320),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_300),
.B(n_303),
.C(n_305),
.Y(n_409)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22x1_ASAP7_75t_L g323 ( 
.A1(n_307),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_307),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_309),
.B(n_448),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_314),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_314),
.B(n_466),
.Y(n_512)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g404 ( 
.A1(n_321),
.A2(n_405),
.B(n_406),
.Y(n_404)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.C(n_330),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_323),
.B(n_328),
.Y(n_370)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_341),
.B(n_343),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_332),
.A2(n_342),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_333),
.A2(n_341),
.B1(n_342),
.B2(n_374),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_338),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_345),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

HAxp5_ASAP7_75t_SL g400 ( 
.A(n_346),
.B(n_347),
.CON(n_400),
.SN(n_400)
);

OAI31xp33_ASAP7_75t_L g347 ( 
.A1(n_348),
.A2(n_349),
.A3(n_352),
.B(n_356),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_361),
.B(n_365),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_382),
.B(n_404),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

NAND2x1p5_ASAP7_75t_L g383 ( 
.A(n_368),
.B(n_371),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.C(n_379),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_376),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_377),
.B(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_378),
.B(n_387),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_383),
.B(n_530),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_402),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_385),
.B(n_402),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_389),
.B(n_401),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_386),
.B(n_442),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_399),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_390),
.B(n_399),
.Y(n_401)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_391),
.B(n_400),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_393),
.C(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_392),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.Y(n_419)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

NOR2x1_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_397),
.Y(n_515)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_400),
.Y(n_545)
);

NOR3xp33_ASAP7_75t_L g528 ( 
.A(n_404),
.B(n_408),
.C(n_529),
.Y(n_528)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_408),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_409),
.B(n_410),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g413 ( 
.A1(n_414),
.A2(n_528),
.B(n_531),
.Y(n_413)
);

AO21x1_ASAP7_75t_L g414 ( 
.A1(n_415),
.A2(n_443),
.B(n_527),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_441),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_416),
.B(n_441),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_420),
.C(n_433),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_456),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_421),
.B(n_433),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_422),
.Y(n_454)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_457),
.B(n_526),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_455),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_445),
.B(n_455),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.C(n_452),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_446),
.A2(n_447),
.B1(n_449),
.B2(n_450),
.Y(n_474)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_474),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_475),
.B(n_525),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_473),
.Y(n_458)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_459),
.B(n_473),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.C(n_464),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_461),
.A2(n_462),
.B1(n_463),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_461),
.Y(n_500)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_465),
.B(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_467),
.B(n_505),
.Y(n_504)
);

INVx6_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx12f_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_501),
.B(n_524),
.Y(n_475)
);

NOR2x1_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_498),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_477),
.B(n_498),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_496),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_478),
.A2(n_479),
.B1(n_496),
.B2(n_497),
.Y(n_507)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_480),
.Y(n_517)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_508),
.B(n_523),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_507),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_SL g523 ( 
.A(n_503),
.B(n_507),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_504),
.B(n_515),
.Y(n_514)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_513),
.B(n_522),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_512),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_512),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_516),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_535),
.A2(n_538),
.B(n_542),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_536),
.B(n_537),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_SL g538 ( 
.A1(n_539),
.A2(n_540),
.B(n_541),
.Y(n_538)
);


endmodule