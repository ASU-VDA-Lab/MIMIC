module fake_jpeg_21197_n_147 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_147);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_147;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx8_ASAP7_75t_SL g65 ( 
.A(n_23),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_0),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_79),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_22),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_74),
.A2(n_62),
.B1(n_65),
.B2(n_59),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_81),
.A2(n_91),
.B1(n_75),
.B2(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_61),
.B1(n_52),
.B2(n_76),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_79),
.B1(n_78),
.B2(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_95),
.B1(n_90),
.B2(n_68),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_60),
.B1(n_53),
.B2(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_104),
.B1(n_57),
.B2(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_85),
.A2(n_78),
.B1(n_50),
.B2(n_72),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_68),
.B(n_66),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_102),
.A2(n_48),
.B(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_88),
.A2(n_63),
.B1(n_71),
.B2(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_102),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_106),
.B(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_119),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_70),
.B1(n_69),
.B2(n_49),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_111),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_110),
.A2(n_2),
.B(n_3),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_50),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_112),
.B(n_113),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_69),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_118),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_1),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_120),
.A2(n_3),
.B(n_4),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_115),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_125),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_126),
.B(n_129),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_116),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_118),
.B1(n_108),
.B2(n_119),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_5),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_133),
.B1(n_127),
.B2(n_8),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_113),
.C(n_114),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_110),
.B(n_117),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_129),
.B(n_122),
.C(n_128),
.D(n_121),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_136),
.A2(n_137),
.B1(n_135),
.B2(n_131),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_135),
.B1(n_32),
.B2(n_33),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_29),
.C(n_45),
.Y(n_140)
);

NAND4xp25_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_27),
.C(n_43),
.D(n_41),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_141),
.A2(n_26),
.B(n_36),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_21),
.C(n_35),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_17),
.B(n_34),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_14),
.C(n_30),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_46),
.B(n_8),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_6),
.Y(n_147)
);


endmodule