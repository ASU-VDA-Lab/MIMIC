module fake_netlist_6_1376_n_1806 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1806);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1806;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_37),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_87),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_55),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_9),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_30),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_23),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_10),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_15),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_134),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_31),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_89),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_84),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_95),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_50),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_7),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_49),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_109),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_67),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_13),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_44),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_51),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_86),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_61),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_25),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_46),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_76),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_72),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_55),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_40),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_122),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_8),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_121),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_119),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_130),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_18),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_38),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_44),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_80),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_14),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_118),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_60),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_58),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_40),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_69),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_1),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_5),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_79),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_36),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_97),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_107),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_8),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_73),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_45),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_141),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_131),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_91),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_1),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_25),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_57),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_6),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_2),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_46),
.Y(n_245)
);

BUFx2_ASAP7_75t_SL g246 ( 
.A(n_42),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_64),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_62),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_45),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_120),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_103),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_16),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_47),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_126),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_146),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_132),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_6),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_114),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_83),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_104),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_96),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_75),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_3),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_150),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_56),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_12),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_52),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_29),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_4),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_77),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_82),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_90),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_94),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_139),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_20),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_125),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_115),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_28),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_24),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_47),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_24),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_128),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_19),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_124),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_20),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_116),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_106),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_53),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_23),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_10),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_100),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_54),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_34),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_102),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_21),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_52),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_149),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_14),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_26),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_22),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_138),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_11),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_37),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_22),
.Y(n_311)
);

INVxp33_ASAP7_75t_SL g312 ( 
.A(n_306),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_162),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_168),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_163),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_168),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_168),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_202),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_195),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_166),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_168),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_205),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_208),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_168),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_212),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_242),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_169),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_169),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_216),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_259),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_211),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_221),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_229),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_169),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_219),
.B(n_0),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_213),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_230),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_237),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_238),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_169),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_169),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_252),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_217),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_206),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_217),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_207),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_194),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_276),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_217),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_217),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_166),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_159),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_159),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_199),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_278),
.B(n_0),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_222),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_160),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_227),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_213),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_231),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_240),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_217),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_241),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_213),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_244),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_251),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_253),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_215),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_215),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_235),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_160),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_173),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_173),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_174),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_174),
.Y(n_378)
);

INVxp33_ASAP7_75t_SL g379 ( 
.A(n_161),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_235),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_176),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_199),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_176),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_256),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_179),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_179),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_180),
.Y(n_387)
);

NAND2x1_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_278),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_158),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

BUFx8_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_267),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_267),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_314),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_316),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_317),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

NAND2x1_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_291),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_291),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_324),
.B(n_158),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_327),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_332),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_328),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_328),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_334),
.B(n_198),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_343),
.B(n_198),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_347),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g418 ( 
.A1(n_358),
.A2(n_257),
.B(n_164),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_351),
.B(n_257),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_351),
.B(n_157),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_365),
.B(n_295),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

CKINVDCx8_ASAP7_75t_R g427 ( 
.A(n_320),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_371),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_372),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_380),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_384),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_384),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_331),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_346),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_313),
.B(n_311),
.Y(n_440)
);

AND2x6_ASAP7_75t_L g441 ( 
.A(n_335),
.B(n_194),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_318),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_322),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_323),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_350),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_325),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_329),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_315),
.B(n_196),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_348),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_375),
.B(n_171),
.Y(n_451)
);

OA21x2_ASAP7_75t_L g452 ( 
.A1(n_336),
.A2(n_256),
.B(n_178),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_320),
.B(n_166),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_338),
.B(n_172),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_340),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_353),
.B(n_239),
.Y(n_456)
);

INVx4_ASAP7_75t_SL g457 ( 
.A(n_441),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_442),
.B(n_353),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_362),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_312),
.B1(n_379),
.B2(n_249),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_246),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_396),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_435),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_442),
.B(n_376),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_423),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_341),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_399),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_392),
.B(n_393),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_344),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g473 ( 
.A1(n_441),
.A2(n_266),
.B1(n_191),
.B2(n_192),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_441),
.A2(n_186),
.B1(n_274),
.B2(n_175),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_442),
.B(n_383),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_441),
.A2(n_271),
.B1(n_285),
.B2(n_200),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_194),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_392),
.Y(n_478)
);

BUFx10_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_452),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_435),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_435),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_194),
.Y(n_483)
);

INVxp33_ASAP7_75t_L g484 ( 
.A(n_440),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_392),
.B(n_393),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_392),
.B(n_387),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_393),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_393),
.B(n_357),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_451),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_399),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_394),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_397),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_397),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_395),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_395),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_444),
.B(n_359),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_440),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_388),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_446),
.B(n_361),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_425),
.B(n_363),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_395),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_444),
.B(n_177),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_449),
.B(n_364),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_449),
.B(n_366),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_449),
.B(n_368),
.Y(n_514)
);

INVx4_ASAP7_75t_SL g515 ( 
.A(n_441),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_451),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_391),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_446),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_L g519 ( 
.A1(n_438),
.A2(n_167),
.B1(n_367),
.B2(n_232),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_399),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_449),
.B(n_369),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_451),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_455),
.B(n_370),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_455),
.B(n_333),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_416),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_416),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_455),
.B(n_226),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_389),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_447),
.B(n_354),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_416),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_405),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_391),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_455),
.B(n_182),
.Y(n_538)
);

AND2x2_ASAP7_75t_SL g539 ( 
.A(n_452),
.B(n_194),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_452),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_405),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_447),
.B(n_355),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_407),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_399),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_399),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_388),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_391),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_391),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_447),
.B(n_360),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_399),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_440),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_422),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_407),
.Y(n_554)
);

INVx8_ASAP7_75t_L g555 ( 
.A(n_441),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_407),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_450),
.B(n_374),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_441),
.A2(n_296),
.B1(n_203),
.B2(n_204),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_R g559 ( 
.A(n_406),
.B(n_319),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_408),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_422),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_438),
.B(n_377),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_422),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_426),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_451),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_438),
.B(n_445),
.Y(n_566)
);

NAND2xp33_ASAP7_75t_L g567 ( 
.A(n_441),
.B(n_201),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_426),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_445),
.B(n_378),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_408),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_381),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_425),
.B(n_214),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_426),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_408),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_452),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_441),
.B(n_452),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_441),
.A2(n_243),
.B1(n_225),
.B2(n_272),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_450),
.B(n_201),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_411),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_441),
.B(n_264),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_450),
.B(n_385),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_425),
.B(n_220),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_391),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_450),
.B(n_386),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_390),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_411),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_450),
.B(n_239),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_441),
.A2(n_418),
.B1(n_425),
.B2(n_450),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_427),
.B(n_239),
.Y(n_590)
);

NAND3xp33_ASAP7_75t_L g591 ( 
.A(n_421),
.B(n_401),
.C(n_403),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_417),
.B(n_188),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_411),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_399),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_414),
.Y(n_595)
);

BUFx4f_ASAP7_75t_L g596 ( 
.A(n_389),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_414),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_414),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_399),
.Y(n_599)
);

AO21x2_ASAP7_75t_L g600 ( 
.A1(n_418),
.A2(n_218),
.B(n_268),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_453),
.A2(n_299),
.B1(n_310),
.B2(n_305),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_424),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_424),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_418),
.A2(n_456),
.B1(n_453),
.B2(n_273),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_427),
.B(n_180),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_424),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_470),
.B(n_439),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_485),
.A2(n_388),
.B(n_400),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_489),
.B(n_443),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_489),
.B(n_443),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g611 ( 
.A(n_459),
.B(n_439),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_586),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_478),
.B(n_443),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_481),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_470),
.B(n_443),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_586),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_467),
.B(n_471),
.Y(n_617)
);

NAND2x1_ASAP7_75t_L g618 ( 
.A(n_505),
.B(n_398),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_540),
.B(n_427),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_586),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

BUFx8_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_566),
.B(n_417),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_492),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_596),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_540),
.B(n_427),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_530),
.B(n_417),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_481),
.B(n_417),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_487),
.B(n_456),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_482),
.B(n_417),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_494),
.B(n_181),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_482),
.B(n_417),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_540),
.B(n_201),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_486),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_L g635 ( 
.A(n_562),
.B(n_406),
.C(n_286),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_494),
.B(n_400),
.Y(n_636)
);

INVx2_ASAP7_75t_SL g637 ( 
.A(n_466),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_577),
.A2(n_400),
.B(n_403),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_508),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_516),
.B(n_430),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_516),
.B(n_430),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_493),
.B(n_326),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_524),
.B(n_430),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_486),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_R g645 ( 
.A(n_472),
.B(n_330),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_508),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_596),
.Y(n_647)
);

OR2x6_ASAP7_75t_L g648 ( 
.A(n_524),
.B(n_418),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_565),
.B(n_181),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_565),
.B(n_430),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_591),
.B(n_430),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_430),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_604),
.B(n_539),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_539),
.B(n_201),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_463),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_503),
.B(n_421),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_539),
.B(n_201),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_512),
.B(n_421),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_573),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_468),
.A2(n_528),
.B1(n_576),
.B2(n_480),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_L g661 ( 
.A1(n_581),
.A2(n_401),
.B(n_420),
.C(n_403),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_570),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_461),
.B(n_187),
.C(n_184),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g664 ( 
.A(n_460),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_463),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_596),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_488),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_555),
.A2(n_413),
.B(n_409),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_521),
.B(n_401),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_460),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_398),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_506),
.B(n_184),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_490),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_572),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g675 ( 
.A(n_559),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_496),
.B(n_501),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_468),
.A2(n_528),
.B1(n_576),
.B2(n_480),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_496),
.B(n_398),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_459),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_468),
.A2(n_287),
.B1(n_284),
.B2(n_289),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_501),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_502),
.B(n_398),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_502),
.B(n_398),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_458),
.B(n_187),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_509),
.B(n_398),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_491),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_509),
.B(n_410),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_491),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_497),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_510),
.B(n_410),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_510),
.B(n_410),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_513),
.B(n_514),
.Y(n_692)
);

NAND3x1_ASAP7_75t_L g693 ( 
.A(n_601),
.B(n_292),
.C(n_297),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_533),
.B(n_428),
.Y(n_694)
);

NAND2x1_ASAP7_75t_L g695 ( 
.A(n_505),
.B(n_410),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_522),
.B(n_410),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_589),
.B(n_210),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_497),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_522),
.B(n_410),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_542),
.B(n_448),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_480),
.A2(n_303),
.B1(n_302),
.B2(n_300),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_573),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_557),
.A2(n_283),
.B1(n_228),
.B2(n_233),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_498),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_525),
.B(n_190),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_528),
.B(n_223),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_523),
.B(n_412),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_523),
.B(n_412),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_576),
.B(n_236),
.Y(n_709)
);

BUFx5_ASAP7_75t_L g710 ( 
.A(n_579),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_531),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_465),
.B(n_190),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_531),
.B(n_412),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_526),
.B(n_247),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_536),
.B(n_412),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_536),
.Y(n_716)
);

AO22x2_ASAP7_75t_L g717 ( 
.A1(n_590),
.A2(n_308),
.B1(n_262),
.B2(n_265),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_475),
.B(n_258),
.Y(n_718)
);

NAND2xp33_ASAP7_75t_L g719 ( 
.A(n_555),
.B(n_258),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_479),
.B(n_250),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_479),
.B(n_280),
.Y(n_721)
);

NOR2x1p5_ASAP7_75t_L g722 ( 
.A(n_583),
.B(n_161),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_479),
.B(n_288),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_541),
.B(n_412),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_498),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_460),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_541),
.B(n_412),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_462),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_543),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_543),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_554),
.B(n_556),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_554),
.B(n_415),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_549),
.B(n_293),
.C(n_261),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_556),
.B(n_415),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_555),
.B(n_261),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_583),
.A2(n_437),
.B(n_429),
.C(n_428),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_560),
.B(n_415),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_460),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_499),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_479),
.B(n_301),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_518),
.B(n_434),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_588),
.B(n_263),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_518),
.B(n_605),
.Y(n_743)
);

NAND3xp33_ASAP7_75t_L g744 ( 
.A(n_582),
.B(n_293),
.C(n_263),
.Y(n_744)
);

OR2x2_ASAP7_75t_SL g745 ( 
.A(n_601),
.B(n_448),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_518),
.B(n_275),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_518),
.B(n_505),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_505),
.B(n_434),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_L g749 ( 
.A1(n_519),
.A2(n_165),
.B1(n_170),
.B2(n_183),
.C(n_185),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_560),
.B(n_415),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_571),
.B(n_415),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_460),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_571),
.B(n_415),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_593),
.B(n_409),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_505),
.B(n_434),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_585),
.B(n_448),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_552),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_593),
.B(n_409),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_462),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_598),
.B(n_413),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_598),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_499),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_546),
.B(n_434),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_462),
.B(n_275),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_546),
.B(n_434),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_L g766 ( 
.A(n_555),
.B(n_279),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_606),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_546),
.B(n_464),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_462),
.B(n_279),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_606),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_507),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_575),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_464),
.B(n_413),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_462),
.B(n_245),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_575),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_464),
.B(n_420),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_580),
.Y(n_777)
);

BUFx12f_ASAP7_75t_L g778 ( 
.A(n_622),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_773),
.A2(n_555),
.B(n_546),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_629),
.A2(n_672),
.B(n_617),
.C(n_680),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_622),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_776),
.A2(n_546),
.B(n_567),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_768),
.A2(n_464),
.B(n_511),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_607),
.B(n_662),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_634),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_660),
.B(n_677),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_669),
.B(n_511),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_768),
.A2(n_464),
.B(n_511),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_SL g790 ( 
.A(n_625),
.B(n_472),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_637),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_668),
.A2(n_538),
.B(n_511),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_736),
.A2(n_592),
.B(n_511),
.C(n_538),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_611),
.B(n_552),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_656),
.B(n_538),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_654),
.A2(n_538),
.B(n_474),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_660),
.B(n_457),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_629),
.A2(n_476),
.B(n_473),
.C(n_578),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_679),
.B(n_484),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_673),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_625),
.A2(n_538),
.B(n_500),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_658),
.B(n_580),
.Y(n_802)
);

A2O1A1Ixp33_ASAP7_75t_L g803 ( 
.A1(n_672),
.A2(n_558),
.B(n_517),
.C(n_537),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_613),
.B(n_587),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_625),
.A2(n_545),
.B(n_500),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_664),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_625),
.A2(n_545),
.B(n_500),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_615),
.B(n_587),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_736),
.A2(n_653),
.B(n_657),
.C(n_654),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_647),
.A2(n_666),
.B(n_633),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_659),
.B(n_517),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_680),
.A2(n_701),
.B(n_653),
.C(n_692),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_702),
.B(n_677),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_694),
.B(n_595),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_671),
.B(n_595),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_657),
.A2(n_602),
.B(n_597),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_681),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_711),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_631),
.B(n_649),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_647),
.A2(n_594),
.B(n_545),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_631),
.B(n_597),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_716),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_633),
.A2(n_603),
.B(n_602),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_674),
.B(n_504),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_729),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_647),
.Y(n_826)
);

O2A1O1Ixp5_ASAP7_75t_L g827 ( 
.A1(n_697),
.A2(n_603),
.B(n_420),
.C(n_534),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_647),
.A2(n_500),
.B(n_599),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_675),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_730),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_666),
.A2(n_545),
.B(n_599),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_761),
.Y(n_832)
);

AO21x1_ASAP7_75t_L g833 ( 
.A1(n_697),
.A2(n_535),
.B(n_534),
.Y(n_833)
);

AOI21xp33_ASAP7_75t_L g834 ( 
.A1(n_705),
.A2(n_584),
.B(n_548),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_757),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_666),
.A2(n_599),
.B(n_594),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_666),
.B(n_457),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_767),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_770),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_638),
.A2(n_599),
.B(n_594),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_649),
.B(n_600),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_639),
.B(n_537),
.Y(n_842)
);

INVx4_ASAP7_75t_L g843 ( 
.A(n_670),
.Y(n_843)
);

AO21x1_ASAP7_75t_L g844 ( 
.A1(n_706),
.A2(n_709),
.B(n_743),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_701),
.A2(n_547),
.B(n_584),
.C(n_548),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_614),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_772),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_754),
.A2(n_594),
.B(n_532),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_646),
.B(n_547),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_609),
.B(n_165),
.Y(n_850)
);

O2A1O1Ixp33_ASAP7_75t_L g851 ( 
.A1(n_706),
.A2(n_507),
.B(n_527),
.C(n_574),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_709),
.A2(n_527),
.B(n_529),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_609),
.B(n_170),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_758),
.A2(n_532),
.B(n_469),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_722),
.B(n_457),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_743),
.B(n_457),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_760),
.B(n_600),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_670),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_651),
.A2(n_529),
.B(n_535),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_746),
.B(n_600),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_692),
.A2(n_747),
.B1(n_759),
.B2(n_728),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_748),
.A2(n_532),
.B(n_495),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_652),
.A2(n_553),
.B(n_574),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_748),
.A2(n_532),
.B(n_495),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_642),
.B(n_245),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_746),
.B(n_469),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_775),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_636),
.B(n_515),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_747),
.B(n_619),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_714),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_703),
.A2(n_579),
.B1(n_483),
.B2(n_477),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_608),
.A2(n_553),
.B(n_569),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_777),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_664),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_712),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_619),
.B(n_515),
.Y(n_876)
);

AOI21x1_ASAP7_75t_L g877 ( 
.A1(n_755),
.A2(n_765),
.B(n_763),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_621),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_627),
.B(n_469),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_626),
.A2(n_477),
.B1(n_483),
.B2(n_579),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_645),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_610),
.A2(n_563),
.B(n_569),
.C(n_568),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_640),
.B(n_469),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_624),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_641),
.A2(n_282),
.B1(n_298),
.B2(n_294),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_755),
.A2(n_532),
.B(n_495),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_763),
.A2(n_532),
.B(n_495),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_643),
.A2(n_282),
.B1(n_298),
.B2(n_294),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_650),
.B(n_520),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_610),
.A2(n_551),
.B(n_568),
.C(n_564),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_765),
.A2(n_544),
.B(n_550),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_623),
.B(n_520),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_676),
.B(n_520),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_719),
.A2(n_544),
.B(n_550),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_684),
.B(n_183),
.Y(n_895)
);

NAND2x1_ASAP7_75t_L g896 ( 
.A(n_670),
.B(n_520),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_731),
.B(n_544),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_705),
.B(n_544),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_684),
.B(n_550),
.Y(n_899)
);

OAI21xp33_ASAP7_75t_L g900 ( 
.A1(n_749),
.A2(n_718),
.B(n_712),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_718),
.B(n_742),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_720),
.A2(n_551),
.B(n_564),
.C(n_563),
.Y(n_902)
);

AOI21x1_ASAP7_75t_L g903 ( 
.A1(n_741),
.A2(n_561),
.B(n_390),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_714),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_735),
.A2(n_550),
.B(n_561),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_714),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_655),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_744),
.B(n_185),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_665),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_766),
.A2(n_515),
.B(n_390),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_700),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_648),
.A2(n_579),
.B(n_483),
.Y(n_912)
);

BUFx8_ASAP7_75t_L g913 ( 
.A(n_756),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_628),
.A2(n_515),
.B(n_390),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_667),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_733),
.B(n_189),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_742),
.A2(n_234),
.B(n_224),
.C(n_197),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_630),
.A2(n_632),
.B(n_618),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_764),
.B(n_579),
.Y(n_919)
);

INVx1_ASAP7_75t_SL g920 ( 
.A(n_645),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_626),
.A2(n_483),
.B1(n_477),
.B2(n_579),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_695),
.A2(n_432),
.B(n_431),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_764),
.B(n_579),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_661),
.A2(n_234),
.B(n_224),
.C(n_197),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_769),
.B(n_477),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_741),
.A2(n_431),
.B(n_432),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_686),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_670),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_688),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_769),
.B(n_720),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_726),
.A2(n_431),
.B(n_432),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_745),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_L g933 ( 
.A1(n_648),
.A2(n_483),
.B(n_477),
.Y(n_933)
);

AO21x1_ASAP7_75t_L g934 ( 
.A1(n_721),
.A2(n_723),
.B(n_740),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_774),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_726),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_SL g937 ( 
.A(n_635),
.B(n_304),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_726),
.A2(n_431),
.B(n_432),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_723),
.A2(n_740),
.B(n_663),
.C(n_753),
.Y(n_939)
);

AOI22x1_ASAP7_75t_L g940 ( 
.A1(n_717),
.A2(n_304),
.B1(n_189),
.B2(n_307),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_648),
.B(n_193),
.Y(n_941)
);

O2A1O1Ixp5_ASAP7_75t_L g942 ( 
.A1(n_678),
.A2(n_428),
.B(n_437),
.C(n_429),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_738),
.A2(n_309),
.B1(n_254),
.B2(n_255),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_703),
.B(n_483),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_682),
.A2(n_193),
.B(n_309),
.C(n_254),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_689),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_683),
.A2(n_483),
.B(n_477),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_698),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_726),
.A2(n_436),
.B(n_433),
.Y(n_949)
);

BUFx4f_ASAP7_75t_L g950 ( 
.A(n_738),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_752),
.A2(n_436),
.B(n_433),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_752),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_703),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_717),
.B(n_433),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_693),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_685),
.A2(n_687),
.B(n_696),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_690),
.A2(n_436),
.B(n_433),
.Y(n_957)
);

NOR2x1p5_ASAP7_75t_L g958 ( 
.A(n_717),
.B(n_255),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_704),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_725),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_739),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_691),
.A2(n_437),
.B(n_429),
.C(n_436),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_762),
.B(n_434),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_699),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_800),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_800),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_846),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_875),
.B(n_707),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_819),
.B(n_771),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_900),
.A2(n_751),
.B(n_750),
.C(n_737),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_901),
.B(n_708),
.Y(n_971)
);

AOI22xp33_ASAP7_75t_SL g972 ( 
.A1(n_895),
.A2(n_245),
.B1(n_260),
.B2(n_269),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_835),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_SL g974 ( 
.A1(n_932),
.A2(n_260),
.B1(n_269),
.B2(n_270),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_780),
.B(n_713),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_846),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_785),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_928),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_779),
.A2(n_732),
.B(n_727),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_780),
.A2(n_812),
.B1(n_787),
.B2(n_798),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_782),
.A2(n_724),
.B(n_715),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_895),
.B(n_734),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_829),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_911),
.B(n_612),
.Y(n_984)
);

O2A1O1Ixp5_ASAP7_75t_L g985 ( 
.A1(n_844),
.A2(n_620),
.B(n_616),
.C(n_710),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_928),
.Y(n_986)
);

INVx2_ASAP7_75t_SL g987 ( 
.A(n_791),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_930),
.B(n_710),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_908),
.A2(n_710),
.B1(n_389),
.B2(n_434),
.Y(n_989)
);

OAI21x1_ASAP7_75t_L g990 ( 
.A1(n_903),
.A2(n_710),
.B(n_389),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_787),
.B(n_307),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_865),
.B(n_270),
.Y(n_992)
);

NAND2x1p5_ASAP7_75t_L g993 ( 
.A(n_826),
.B(n_434),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_786),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_909),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_840),
.A2(n_710),
.B(n_389),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_802),
.B(n_434),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_801),
.A2(n_419),
.B(n_404),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_824),
.B(n_290),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_810),
.A2(n_419),
.B(n_404),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_824),
.B(n_794),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_826),
.B(n_434),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_797),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_964),
.B(n_290),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_792),
.A2(n_419),
.B(n_404),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_R g1006 ( 
.A(n_778),
.B(n_281),
.Y(n_1006)
);

OR2x6_ASAP7_75t_SL g1007 ( 
.A(n_799),
.B(n_277),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_SL g1008 ( 
.A(n_812),
.B(n_277),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_797),
.A2(n_419),
.B(n_404),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_913),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_959),
.B(n_281),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_781),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_SL g1013 ( 
.A(n_917),
.B(n_3),
.C(n_4),
.Y(n_1013)
);

INVxp33_ASAP7_75t_SL g1014 ( 
.A(n_920),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_935),
.B(n_63),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_817),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_964),
.B(n_419),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_813),
.B(n_389),
.Y(n_1018)
);

O2A1O1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_917),
.A2(n_11),
.B(n_12),
.C(n_15),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_904),
.B(n_16),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_881),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_804),
.A2(n_419),
.B(n_404),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_908),
.A2(n_419),
.B(n_404),
.C(n_399),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_811),
.B(n_419),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_830),
.B(n_419),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_809),
.A2(n_389),
.B(n_419),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_928),
.Y(n_1027)
);

OR2x6_ASAP7_75t_L g1028 ( 
.A(n_781),
.B(n_404),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_791),
.Y(n_1029)
);

O2A1O1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_945),
.A2(n_916),
.B(n_924),
.C(n_953),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_916),
.A2(n_389),
.B1(n_404),
.B2(n_21),
.Y(n_1031)
);

AO22x1_ASAP7_75t_L g1032 ( 
.A1(n_913),
.A2(n_389),
.B1(n_18),
.B2(n_26),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_855),
.B(n_71),
.Y(n_1033)
);

NAND2x1p5_ASAP7_75t_L g1034 ( 
.A(n_843),
.B(n_404),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_928),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_808),
.A2(n_404),
.B(n_66),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_941),
.B(n_17),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_839),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_SL g1039 ( 
.A(n_937),
.B(n_17),
.C(n_27),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_818),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_952),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_822),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_945),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_924),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_955),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_955),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_850),
.B(n_33),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_850),
.B(n_35),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_861),
.A2(n_35),
.B(n_38),
.C(n_39),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_798),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_853),
.B(n_41),
.Y(n_1051)
);

AOI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_842),
.A2(n_389),
.B1(n_93),
.B2(n_101),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_842),
.A2(n_389),
.B1(n_92),
.B2(n_105),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_943),
.B(n_48),
.C(n_50),
.Y(n_1054)
);

NOR2xp67_ASAP7_75t_SL g1055 ( 
.A(n_843),
.B(n_48),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_858),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_853),
.B(n_51),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_L g1058 ( 
.A1(n_876),
.A2(n_389),
.B(n_133),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_805),
.A2(n_108),
.B(n_155),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_825),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_849),
.A2(n_389),
.B1(n_85),
.B2(n_137),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_795),
.B(n_81),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_832),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_R g1064 ( 
.A(n_870),
.B(n_78),
.Y(n_1064)
);

NOR3xp33_ASAP7_75t_SL g1065 ( 
.A(n_885),
.B(n_53),
.C(n_54),
.Y(n_1065)
);

CKINVDCx14_ASAP7_75t_R g1066 ( 
.A(n_855),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_807),
.A2(n_142),
.B(n_59),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_788),
.A2(n_56),
.B(n_65),
.C(n_74),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_796),
.A2(n_140),
.B1(n_145),
.B2(n_147),
.Y(n_1069)
);

OR2x6_ASAP7_75t_L g1070 ( 
.A(n_811),
.B(n_151),
.Y(n_1070)
);

O2A1O1Ixp5_ASAP7_75t_L g1071 ( 
.A1(n_869),
.A2(n_152),
.B(n_934),
.C(n_841),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_952),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_820),
.A2(n_836),
.B(n_831),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_828),
.A2(n_815),
.B(n_869),
.Y(n_1074)
);

A2O1A1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_849),
.A2(n_790),
.B(n_834),
.C(n_793),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_906),
.B(n_838),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_847),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_867),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_910),
.A2(n_918),
.B(n_898),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_940),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_821),
.B(n_960),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_961),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_950),
.B(n_860),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_857),
.A2(n_845),
.B1(n_803),
.B2(n_958),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_950),
.B(n_939),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_845),
.A2(n_803),
.B1(n_871),
.B2(n_856),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_858),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_888),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_783),
.A2(n_789),
.B(n_893),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_806),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_873),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_866),
.B(n_897),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_952),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_899),
.B(n_856),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_961),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_952),
.Y(n_1096)
);

BUFx3_ASAP7_75t_L g1097 ( 
.A(n_907),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_915),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_806),
.B(n_874),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_927),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_871),
.A2(n_944),
.B1(n_954),
.B2(n_814),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_946),
.B(n_892),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_929),
.B(n_948),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_936),
.B(n_874),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_936),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_946),
.B(n_879),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_876),
.A2(n_894),
.B(n_868),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_L g1108 ( 
.A(n_919),
.B(n_923),
.C(n_925),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_883),
.B(n_889),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_868),
.B(n_884),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1079),
.A2(n_872),
.B(n_905),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1001),
.B(n_878),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1047),
.A2(n_942),
.B(n_837),
.C(n_962),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_973),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1073),
.A2(n_863),
.B(n_859),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_977),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_968),
.B(n_854),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_1029),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_1056),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_983),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1089),
.A2(n_823),
.B(n_848),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_971),
.B(n_816),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1074),
.A2(n_914),
.B(n_837),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_982),
.B(n_956),
.Y(n_1124)
);

AO32x2_ASAP7_75t_L g1125 ( 
.A1(n_980),
.A2(n_833),
.A3(n_827),
.B1(n_877),
.B2(n_882),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1045),
.Y(n_1126)
);

AOI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_972),
.A2(n_890),
.B1(n_902),
.B2(n_957),
.C(n_926),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_995),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1048),
.A2(n_933),
.B(n_912),
.C(n_851),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_L g1130 ( 
.A1(n_1107),
.A2(n_852),
.B(n_891),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1092),
.A2(n_896),
.B(n_947),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_994),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1092),
.A2(n_862),
.B(n_864),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1081),
.B(n_951),
.Y(n_1134)
);

AO32x2_ASAP7_75t_L g1135 ( 
.A1(n_980),
.A2(n_880),
.A3(n_921),
.B1(n_963),
.B2(n_922),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1084),
.A2(n_931),
.A3(n_938),
.B(n_949),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_1012),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1057),
.A2(n_886),
.B(n_887),
.C(n_1030),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1099),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_SL g1140 ( 
.A1(n_1069),
.A2(n_1085),
.B(n_1083),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_1046),
.Y(n_1141)
);

BUFx2_ASAP7_75t_R g1142 ( 
.A(n_1021),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1109),
.A2(n_979),
.B(n_981),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1050),
.A2(n_1051),
.B1(n_1003),
.B2(n_975),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_978),
.Y(n_1145)
);

NAND3xp33_ASAP7_75t_L g1146 ( 
.A(n_1065),
.B(n_1008),
.C(n_1054),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1016),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_L g1148 ( 
.A1(n_1005),
.A2(n_998),
.B(n_996),
.Y(n_1148)
);

BUFx4f_ASAP7_75t_SL g1149 ( 
.A(n_1010),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1008),
.A2(n_1088),
.B(n_1071),
.C(n_991),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_1014),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_978),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_987),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_975),
.A2(n_1094),
.B(n_1075),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1069),
.A2(n_1049),
.B(n_1084),
.C(n_1062),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1026),
.A2(n_1000),
.B(n_985),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1004),
.B(n_999),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1038),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1050),
.A2(n_1039),
.B(n_1019),
.C(n_1044),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1108),
.A2(n_1086),
.B(n_1094),
.Y(n_1160)
);

OAI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1037),
.A2(n_1070),
.B1(n_1011),
.B2(n_1080),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1026),
.A2(n_990),
.B(n_1009),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1022),
.A2(n_1058),
.B(n_988),
.Y(n_1163)
);

AOI221xp5_ASAP7_75t_SL g1164 ( 
.A1(n_1043),
.A2(n_1086),
.B1(n_1101),
.B2(n_1031),
.C(n_969),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1023),
.A2(n_1101),
.A3(n_1062),
.B(n_1110),
.Y(n_1165)
);

INVxp67_ASAP7_75t_L g1166 ( 
.A(n_1076),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1077),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_974),
.A2(n_1020),
.B1(n_992),
.B2(n_1013),
.C(n_1091),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_970),
.A2(n_997),
.B(n_1018),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_L g1170 ( 
.A(n_984),
.B(n_1068),
.C(n_1042),
.Y(n_1170)
);

AO21x1_ASAP7_75t_L g1171 ( 
.A1(n_1036),
.A2(n_1102),
.B(n_1067),
.Y(n_1171)
);

AND2x4_ASAP7_75t_SL g1172 ( 
.A(n_1087),
.B(n_1033),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1102),
.A2(n_1106),
.B(n_1017),
.Y(n_1173)
);

OAI221xp5_ASAP7_75t_SL g1174 ( 
.A1(n_1070),
.A2(n_1053),
.B1(n_1052),
.B2(n_1061),
.C(n_1007),
.Y(n_1174)
);

AO21x2_ASAP7_75t_L g1175 ( 
.A1(n_1059),
.A2(n_1025),
.B(n_966),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1082),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_993),
.A2(n_1002),
.B(n_1034),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_965),
.B(n_967),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1056),
.A2(n_1027),
.B(n_1099),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_976),
.B(n_1100),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1103),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1078),
.A2(n_1063),
.B(n_1060),
.C(n_1040),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_SL g1183 ( 
.A1(n_1033),
.A2(n_1070),
.B(n_1087),
.Y(n_1183)
);

CKINVDCx11_ASAP7_75t_R g1184 ( 
.A(n_1028),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1056),
.A2(n_1027),
.B(n_1024),
.Y(n_1185)
);

NAND3xp33_ASAP7_75t_L g1186 ( 
.A(n_1055),
.B(n_1098),
.C(n_1097),
.Y(n_1186)
);

INVx3_ASAP7_75t_L g1187 ( 
.A(n_1041),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1095),
.A2(n_1015),
.B(n_1028),
.C(n_1090),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_993),
.A2(n_1002),
.B(n_1034),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1056),
.A2(n_1027),
.B(n_1090),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1015),
.B(n_1105),
.Y(n_1191)
);

INVx3_ASAP7_75t_SL g1192 ( 
.A(n_1028),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1027),
.A2(n_989),
.B(n_1035),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1066),
.A2(n_1032),
.B(n_1064),
.C(n_1006),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1035),
.A2(n_1104),
.B(n_1041),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1041),
.A2(n_1072),
.B(n_1093),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_SL g1197 ( 
.A(n_978),
.B(n_986),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_986),
.A2(n_1072),
.B(n_1093),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1072),
.A2(n_1093),
.B(n_1096),
.Y(n_1199)
);

AO31x2_ASAP7_75t_L g1200 ( 
.A1(n_986),
.A2(n_1084),
.A3(n_980),
.B(n_1086),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1096),
.A2(n_901),
.B1(n_1008),
.B2(n_895),
.Y(n_1201)
);

NAND3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1096),
.B(n_900),
.C(n_901),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1001),
.B(n_784),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1084),
.A2(n_980),
.A3(n_1086),
.B(n_844),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_973),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_1047),
.A2(n_900),
.B(n_780),
.C(n_901),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1047),
.A2(n_900),
.B(n_780),
.C(n_901),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1001),
.B(n_784),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1001),
.B(n_784),
.Y(n_1209)
);

AOI221x1_ASAP7_75t_L g1210 ( 
.A1(n_980),
.A2(n_1050),
.B1(n_900),
.B2(n_780),
.C(n_1084),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1014),
.B(n_662),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1073),
.A2(n_1107),
.B(n_979),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_973),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_971),
.B(n_780),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_980),
.A2(n_780),
.B(n_1084),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_977),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1014),
.B(n_662),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_980),
.A2(n_780),
.B(n_1084),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1099),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1073),
.A2(n_1107),
.B(n_979),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_980),
.A2(n_780),
.B(n_1084),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_978),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_971),
.B(n_780),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1047),
.A2(n_901),
.B(n_900),
.C(n_674),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1001),
.B(n_784),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_977),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_983),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1084),
.A2(n_980),
.A3(n_1086),
.B(n_844),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_973),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_980),
.A2(n_780),
.B1(n_812),
.B2(n_787),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1029),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1047),
.A2(n_900),
.B(n_780),
.C(n_901),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1014),
.B(n_662),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_973),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1047),
.A2(n_901),
.B(n_900),
.C(n_674),
.Y(n_1242)
);

A2O1A1Ixp33_ASAP7_75t_L g1243 ( 
.A1(n_1047),
.A2(n_900),
.B(n_780),
.C(n_901),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1047),
.A2(n_900),
.B(n_780),
.C(n_901),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_983),
.B(n_875),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1247)
);

AOI221x1_ASAP7_75t_L g1248 ( 
.A1(n_980),
.A2(n_1050),
.B1(n_900),
.B2(n_780),
.C(n_1084),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_980),
.A2(n_780),
.B(n_1084),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1079),
.A2(n_647),
.B(n_625),
.Y(n_1250)
);

AO31x2_ASAP7_75t_L g1251 ( 
.A1(n_1084),
.A2(n_980),
.A3(n_1086),
.B(n_844),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1047),
.A2(n_901),
.B(n_900),
.C(n_674),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_SL g1253 ( 
.A1(n_1069),
.A2(n_787),
.B(n_780),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_995),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1011),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_R g1256 ( 
.A(n_1010),
.B(n_406),
.Y(n_1256)
);

BUFx2_ASAP7_75t_L g1257 ( 
.A(n_1205),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1116),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1166),
.A2(n_1211),
.B1(n_1223),
.B2(n_1240),
.Y(n_1259)
);

OAI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_1245),
.A2(n_1155),
.B1(n_1157),
.B2(n_1146),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1146),
.A2(n_1227),
.B1(n_1216),
.B2(n_1249),
.Y(n_1261)
);

BUFx2_ASAP7_75t_SL g1262 ( 
.A(n_1241),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1137),
.Y(n_1263)
);

BUFx4f_ASAP7_75t_SL g1264 ( 
.A(n_1114),
.Y(n_1264)
);

BUFx4_ASAP7_75t_R g1265 ( 
.A(n_1255),
.Y(n_1265)
);

CKINVDCx8_ASAP7_75t_R g1266 ( 
.A(n_1120),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1132),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1145),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1210),
.A2(n_1248),
.B1(n_1237),
.B2(n_1227),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1209),
.B(n_1232),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1216),
.A2(n_1224),
.B1(n_1249),
.B2(n_1237),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_SL g1273 ( 
.A1(n_1224),
.A2(n_1201),
.B1(n_1144),
.B2(n_1160),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1234),
.Y(n_1274)
);

INVx8_ASAP7_75t_L g1275 ( 
.A(n_1145),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1144),
.A2(n_1161),
.B1(n_1160),
.B2(n_1168),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1147),
.Y(n_1277)
);

INVx1_ASAP7_75t_SL g1278 ( 
.A(n_1114),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1213),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1236),
.Y(n_1280)
);

INVx6_ASAP7_75t_L g1281 ( 
.A(n_1119),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1158),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1167),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1222),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1202),
.A2(n_1229),
.B1(n_1214),
.B2(n_1170),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1174),
.A2(n_1170),
.B1(n_1243),
.B2(n_1206),
.Y(n_1286)
);

INVx1_ASAP7_75t_SL g1287 ( 
.A(n_1126),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1255),
.A2(n_1186),
.B1(n_1229),
.B2(n_1214),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1233),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1254),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1181),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1151),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1178),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1126),
.A2(n_1186),
.B1(n_1117),
.B2(n_1122),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1180),
.Y(n_1295)
);

BUFx8_ASAP7_75t_L g1296 ( 
.A(n_1141),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1180),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1159),
.A2(n_1242),
.B(n_1231),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1112),
.B(n_1252),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1178),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1253),
.A2(n_1149),
.B1(n_1197),
.B2(n_1154),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1145),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1182),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1142),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1134),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1184),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1207),
.B(n_1239),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1139),
.B(n_1225),
.Y(n_1308)
);

BUFx12f_ASAP7_75t_L g1309 ( 
.A(n_1176),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1139),
.Y(n_1310)
);

OAI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1124),
.A2(n_1197),
.B1(n_1192),
.B2(n_1118),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1119),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1169),
.A2(n_1124),
.B1(n_1127),
.B2(n_1171),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1225),
.Y(n_1314)
);

INVx6_ASAP7_75t_L g1315 ( 
.A(n_1191),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1238),
.A2(n_1153),
.B1(n_1169),
.B2(n_1173),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_1191),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1200),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1164),
.A2(n_1244),
.B1(n_1172),
.B2(n_1150),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1187),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1164),
.A2(n_1175),
.B1(n_1131),
.B2(n_1143),
.Y(n_1321)
);

OAI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1193),
.A2(n_1140),
.B1(n_1195),
.B2(n_1185),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1152),
.Y(n_1323)
);

INVx1_ASAP7_75t_SL g1324 ( 
.A(n_1187),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1183),
.A2(n_1188),
.B1(n_1194),
.B2(n_1138),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1152),
.Y(n_1326)
);

CKINVDCx6p67_ASAP7_75t_R g1327 ( 
.A(n_1228),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1196),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1228),
.Y(n_1329)
);

OAI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1195),
.A2(n_1179),
.B1(n_1228),
.B2(n_1204),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1199),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1199),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1204),
.Y(n_1333)
);

OR2x2_ASAP7_75t_L g1334 ( 
.A(n_1204),
.B(n_1251),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1175),
.A2(n_1133),
.B1(n_1111),
.B2(n_1115),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1156),
.B2(n_1121),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1235),
.A2(n_1251),
.B1(n_1250),
.B2(n_1221),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1235),
.A2(n_1220),
.B1(n_1247),
.B2(n_1246),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1198),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1177),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1136),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1215),
.A2(n_1230),
.B1(n_1219),
.B2(n_1218),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1256),
.Y(n_1343)
);

INVx6_ASAP7_75t_L g1344 ( 
.A(n_1190),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1165),
.Y(n_1345)
);

INVx2_ASAP7_75t_SL g1346 ( 
.A(n_1189),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_1123),
.Y(n_1347)
);

INVxp33_ASAP7_75t_SL g1348 ( 
.A(n_1217),
.Y(n_1348)
);

BUFx10_ASAP7_75t_L g1349 ( 
.A(n_1129),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1165),
.B(n_1113),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1135),
.A2(n_1125),
.B1(n_1162),
.B2(n_1130),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1212),
.A2(n_1226),
.B1(n_1148),
.B2(n_1163),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1135),
.A2(n_700),
.B1(n_756),
.B2(n_900),
.Y(n_1353)
);

CKINVDCx6p67_ASAP7_75t_R g1354 ( 
.A(n_1135),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1125),
.B(n_1203),
.Y(n_1355)
);

INVx4_ASAP7_75t_L g1356 ( 
.A(n_1125),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1128),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1146),
.A2(n_900),
.B1(n_895),
.B2(n_901),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1119),
.Y(n_1361)
);

BUFx2_ASAP7_75t_R g1362 ( 
.A(n_1120),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1128),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1241),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1116),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1114),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1241),
.Y(n_1367)
);

CKINVDCx8_ASAP7_75t_R g1368 ( 
.A(n_1120),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1146),
.A2(n_1008),
.B1(n_1050),
.B2(n_895),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1146),
.A2(n_1008),
.B1(n_901),
.B2(n_1050),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1146),
.A2(n_900),
.B1(n_895),
.B2(n_901),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1241),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1137),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1145),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1211),
.A2(n_700),
.B1(n_756),
.B2(n_900),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1128),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1128),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1128),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1166),
.A2(n_901),
.B1(n_674),
.B2(n_662),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1146),
.A2(n_900),
.B1(n_895),
.B2(n_901),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1161),
.A2(n_700),
.B(n_756),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1166),
.A2(n_901),
.B1(n_674),
.B2(n_662),
.Y(n_1382)
);

OAI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1146),
.A2(n_1008),
.B1(n_901),
.B2(n_1050),
.Y(n_1383)
);

CKINVDCx11_ASAP7_75t_R g1384 ( 
.A(n_1114),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1146),
.A2(n_900),
.B1(n_895),
.B2(n_901),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1203),
.B(n_1208),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1281),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1340),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1318),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1335),
.A2(n_1321),
.B(n_1341),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1346),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1355),
.B(n_1354),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1318),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1347),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1333),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1286),
.A2(n_1260),
.B1(n_1325),
.B2(n_1307),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1334),
.B(n_1345),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1316),
.A2(n_1269),
.B(n_1350),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1258),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1328),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1273),
.B(n_1272),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1299),
.B(n_1358),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1276),
.A2(n_1369),
.B1(n_1272),
.B2(n_1261),
.Y(n_1403)
);

AO21x2_ASAP7_75t_L g1404 ( 
.A1(n_1316),
.A2(n_1269),
.B(n_1351),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1267),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1356),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1335),
.A2(n_1321),
.B(n_1313),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1273),
.B(n_1261),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1270),
.B(n_1271),
.Y(n_1409)
);

OAI21xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1276),
.A2(n_1319),
.B(n_1358),
.Y(n_1410)
);

INVx5_ASAP7_75t_L g1411 ( 
.A(n_1344),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1369),
.A2(n_1371),
.B1(n_1380),
.B2(n_1385),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1356),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1371),
.A2(n_1380),
.B1(n_1385),
.B2(n_1370),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1305),
.B(n_1353),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1293),
.B(n_1300),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1298),
.A2(n_1383),
.B(n_1370),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1277),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1349),
.B(n_1285),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1282),
.Y(n_1420)
);

INVx11_ASAP7_75t_L g1421 ( 
.A(n_1296),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1283),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1284),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1295),
.B(n_1297),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1285),
.B(n_1313),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1289),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1365),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1287),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1339),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1336),
.Y(n_1430)
);

INVx2_ASAP7_75t_SL g1431 ( 
.A(n_1281),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_SL g1432 ( 
.A1(n_1303),
.A2(n_1331),
.B(n_1332),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1349),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1320),
.Y(n_1434)
);

INVx2_ASAP7_75t_SL g1435 ( 
.A(n_1281),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1291),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1257),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1274),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1383),
.A2(n_1375),
.B1(n_1288),
.B2(n_1301),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1279),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1312),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1336),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1351),
.Y(n_1443)
);

INVx2_ASAP7_75t_SL g1444 ( 
.A(n_1312),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1337),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1381),
.A2(n_1348),
.B1(n_1259),
.B2(n_1264),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1386),
.B(n_1359),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1337),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1278),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1379),
.A2(n_1382),
.B1(n_1317),
.B2(n_1366),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1290),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_SL g1452 ( 
.A(n_1292),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1357),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1363),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1376),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1377),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1378),
.Y(n_1457)
);

INVxp33_ASAP7_75t_L g1458 ( 
.A(n_1360),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1330),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1344),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1330),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1311),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1294),
.A2(n_1288),
.B1(n_1322),
.B2(n_1311),
.C(n_1301),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1308),
.B(n_1310),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1338),
.A2(n_1342),
.B(n_1352),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1344),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1294),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1352),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1338),
.Y(n_1469)
);

OA21x2_ASAP7_75t_L g1470 ( 
.A1(n_1342),
.A2(n_1314),
.B(n_1322),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1280),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1312),
.A2(n_1361),
.B(n_1265),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1268),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1268),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1324),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1302),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1264),
.A2(n_1304),
.B1(n_1315),
.B2(n_1309),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1361),
.B(n_1302),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1374),
.Y(n_1479)
);

INVx4_ASAP7_75t_L g1480 ( 
.A(n_1275),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1262),
.B(n_1275),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1407),
.A2(n_1329),
.B(n_1326),
.Y(n_1482)
);

NOR2x1_ASAP7_75t_SL g1483 ( 
.A(n_1411),
.B(n_1263),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1411),
.A2(n_1465),
.B(n_1463),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1417),
.A2(n_1373),
.B(n_1364),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1389),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1464),
.B(n_1384),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1472),
.B(n_1265),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_SL g1489 ( 
.A1(n_1432),
.A2(n_1306),
.B(n_1362),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_SL g1490 ( 
.A1(n_1432),
.A2(n_1296),
.B(n_1327),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1402),
.B(n_1367),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1410),
.B(n_1367),
.Y(n_1492)
);

O2A1O1Ixp33_ASAP7_75t_SL g1493 ( 
.A1(n_1425),
.A2(n_1343),
.B(n_1275),
.C(n_1323),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1464),
.B(n_1367),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1410),
.A2(n_1372),
.B1(n_1343),
.B2(n_1368),
.C(n_1266),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1462),
.B(n_1323),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1388),
.B(n_1418),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1429),
.Y(n_1498)
);

AND2x4_ASAP7_75t_L g1499 ( 
.A(n_1388),
.B(n_1420),
.Y(n_1499)
);

OAI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1396),
.A2(n_1414),
.B(n_1412),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1394),
.B(n_1392),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_1433),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1394),
.B(n_1392),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1419),
.B(n_1458),
.Y(n_1504)
);

NOR2x1_ASAP7_75t_SL g1505 ( 
.A(n_1411),
.B(n_1481),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1420),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1399),
.B(n_1405),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_SL g1508 ( 
.A(n_1452),
.B(n_1438),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1439),
.A2(n_1403),
.B(n_1446),
.Y(n_1509)
);

AOI211xp5_ASAP7_75t_L g1510 ( 
.A1(n_1408),
.A2(n_1467),
.B(n_1401),
.C(n_1419),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1425),
.A2(n_1408),
.B1(n_1401),
.B2(n_1450),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1433),
.A2(n_1450),
.B(n_1415),
.Y(n_1512)
);

AO21x2_ASAP7_75t_L g1513 ( 
.A1(n_1390),
.A2(n_1404),
.B(n_1468),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1422),
.B(n_1427),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1436),
.B(n_1409),
.Y(n_1515)
);

AO32x2_ASAP7_75t_L g1516 ( 
.A1(n_1443),
.A2(n_1406),
.A3(n_1413),
.B1(n_1404),
.B2(n_1389),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1416),
.B(n_1428),
.Y(n_1517)
);

AND2x4_ASAP7_75t_L g1518 ( 
.A(n_1388),
.B(n_1423),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1471),
.A2(n_1447),
.B1(n_1477),
.B2(n_1440),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1437),
.B(n_1449),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1426),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1421),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1471),
.B(n_1434),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1481),
.A2(n_1469),
.B1(n_1387),
.B2(n_1441),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1421),
.A2(n_1475),
.B1(n_1481),
.B2(n_1469),
.Y(n_1525)
);

AO32x2_ASAP7_75t_L g1526 ( 
.A1(n_1443),
.A2(n_1413),
.A3(n_1406),
.B1(n_1404),
.B2(n_1398),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1388),
.B(n_1426),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1470),
.B(n_1445),
.C(n_1448),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1398),
.A2(n_1448),
.B1(n_1445),
.B2(n_1461),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1397),
.B(n_1459),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1424),
.B(n_1453),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_SL g1533 ( 
.A1(n_1481),
.A2(n_1387),
.B(n_1441),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1453),
.B(n_1455),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1466),
.A2(n_1460),
.B(n_1470),
.Y(n_1535)
);

A2O1A1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1459),
.A2(n_1461),
.B(n_1430),
.C(n_1442),
.Y(n_1536)
);

NAND3xp33_ASAP7_75t_L g1537 ( 
.A(n_1470),
.B(n_1466),
.C(n_1468),
.Y(n_1537)
);

AND4x1_ASAP7_75t_L g1538 ( 
.A(n_1473),
.B(n_1476),
.C(n_1479),
.D(n_1474),
.Y(n_1538)
);

OAI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1466),
.A2(n_1460),
.B(n_1470),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1486),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1521),
.B(n_1398),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1500),
.A2(n_1465),
.B1(n_1430),
.B2(n_1442),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1482),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1498),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1465),
.Y(n_1545)
);

OAI221xp5_ASAP7_75t_L g1546 ( 
.A1(n_1509),
.A2(n_1465),
.B1(n_1460),
.B2(n_1411),
.C(n_1456),
.Y(n_1546)
);

AOI21xp5_ASAP7_75t_SL g1547 ( 
.A1(n_1495),
.A2(n_1441),
.B(n_1444),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1482),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1400),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1506),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1400),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1497),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1507),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1507),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1516),
.B(n_1400),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1516),
.B(n_1482),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1530),
.B(n_1397),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1521),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1537),
.B(n_1393),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1526),
.B(n_1535),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1514),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1529),
.B(n_1395),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1497),
.B(n_1391),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1497),
.Y(n_1564)
);

INVxp67_ASAP7_75t_L g1565 ( 
.A(n_1504),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1495),
.A2(n_1456),
.B1(n_1455),
.B2(n_1457),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1564),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1549),
.B(n_1526),
.Y(n_1568)
);

AND2x4_ASAP7_75t_L g1569 ( 
.A(n_1552),
.B(n_1505),
.Y(n_1569)
);

INVx5_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

OAI31xp33_ASAP7_75t_L g1571 ( 
.A1(n_1546),
.A2(n_1511),
.A3(n_1492),
.B(n_1519),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1564),
.B(n_1523),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1564),
.B(n_1501),
.Y(n_1573)
);

INVx4_ASAP7_75t_L g1574 ( 
.A(n_1563),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1557),
.B(n_1528),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1564),
.B(n_1503),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1558),
.B(n_1515),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1558),
.B(n_1536),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1565),
.B(n_1499),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1565),
.B(n_1499),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1552),
.B(n_1499),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1550),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1544),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1549),
.B(n_1527),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1543),
.Y(n_1585)
);

NAND4xp25_ASAP7_75t_L g1586 ( 
.A(n_1542),
.B(n_1510),
.C(n_1512),
.D(n_1492),
.Y(n_1586)
);

NAND4xp25_ASAP7_75t_SL g1587 ( 
.A(n_1547),
.B(n_1484),
.C(n_1485),
.D(n_1536),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1540),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1550),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1491),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1550),
.Y(n_1591)
);

AOI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1542),
.A2(n_1546),
.B1(n_1484),
.B2(n_1560),
.C(n_1562),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1554),
.B(n_1518),
.Y(n_1593)
);

OAI33xp33_ASAP7_75t_L g1594 ( 
.A1(n_1541),
.A2(n_1517),
.A3(n_1531),
.B1(n_1525),
.B2(n_1532),
.B3(n_1534),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1543),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1566),
.B(n_1538),
.C(n_1520),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1566),
.A2(n_1524),
.B1(n_1502),
.B2(n_1488),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1557),
.B(n_1539),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1545),
.A2(n_1488),
.B1(n_1496),
.B2(n_1520),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1575),
.B(n_1541),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1568),
.B(n_1560),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1568),
.B(n_1560),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1582),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1583),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1575),
.B(n_1556),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1595),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1577),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1560),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1582),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1578),
.B(n_1561),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1584),
.B(n_1556),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1584),
.B(n_1556),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1574),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1584),
.B(n_1570),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1589),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1574),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1598),
.B(n_1540),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1595),
.B(n_1548),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1591),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1583),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1585),
.B(n_1548),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1570),
.B(n_1549),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1583),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1598),
.B(n_1585),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1570),
.B(n_1551),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1570),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1588),
.B(n_1548),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1574),
.B(n_1551),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1591),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1574),
.B(n_1551),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1567),
.B(n_1555),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1606),
.Y(n_1635)
);

OAI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1607),
.A2(n_1586),
.B1(n_1596),
.B2(n_1599),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1606),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1610),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1607),
.B(n_1590),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1610),
.B(n_1596),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1616),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1615),
.B(n_1569),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1623),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1600),
.B(n_1614),
.Y(n_1644)
);

INVxp67_ASAP7_75t_SL g1645 ( 
.A(n_1619),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1619),
.B(n_1588),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1623),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1614),
.A2(n_1587),
.B1(n_1592),
.B2(n_1597),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1615),
.B(n_1569),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1600),
.B(n_1627),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1616),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1623),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1569),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1616),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1632),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1627),
.B(n_1571),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1632),
.Y(n_1657)
);

NAND4xp25_ASAP7_75t_L g1658 ( 
.A(n_1605),
.B(n_1592),
.C(n_1571),
.D(n_1586),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1605),
.B(n_1559),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1605),
.B(n_1579),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1613),
.B(n_1522),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1630),
.B(n_1579),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1630),
.B(n_1580),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1601),
.B(n_1569),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1630),
.B(n_1559),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1601),
.B(n_1581),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1632),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1603),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1601),
.B(n_1580),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1603),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1624),
.A2(n_1587),
.B(n_1545),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1609),
.Y(n_1672)
);

NAND2x1p5_ASAP7_75t_L g1673 ( 
.A(n_1629),
.B(n_1559),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1613),
.B(n_1522),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1602),
.B(n_1608),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1602),
.B(n_1581),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1651),
.Y(n_1677)
);

OAI21xp33_ASAP7_75t_L g1678 ( 
.A1(n_1658),
.A2(n_1599),
.B(n_1545),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1673),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1651),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1650),
.B(n_1620),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1629),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1655),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1655),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1672),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1675),
.B(n_1602),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1672),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1639),
.B(n_1572),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1641),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1664),
.B(n_1608),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1636),
.B(n_1572),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1664),
.B(n_1608),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1640),
.B(n_1573),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1656),
.B(n_1573),
.Y(n_1694)
);

OAI31xp33_ASAP7_75t_L g1695 ( 
.A1(n_1671),
.A2(n_1638),
.A3(n_1597),
.B(n_1673),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1673),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1648),
.B(n_1576),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1645),
.B(n_1576),
.Y(n_1699)
);

INVxp67_ASAP7_75t_L g1700 ( 
.A(n_1661),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1654),
.Y(n_1701)
);

NOR2x1_ASAP7_75t_L g1702 ( 
.A(n_1674),
.B(n_1613),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1644),
.B(n_1593),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1704)
);

AOI211xp5_ASAP7_75t_L g1705 ( 
.A1(n_1650),
.A2(n_1594),
.B(n_1545),
.C(n_1493),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1649),
.B(n_1618),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1669),
.B(n_1620),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1657),
.Y(n_1708)
);

INVxp67_ASAP7_75t_L g1709 ( 
.A(n_1646),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1667),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1649),
.B(n_1611),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1678),
.A2(n_1594),
.B1(n_1653),
.B2(n_1663),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1709),
.B(n_1666),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1682),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1698),
.B(n_1666),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1702),
.B(n_1653),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1696),
.B(n_1676),
.Y(n_1717)
);

AOI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1700),
.A2(n_1662),
.B1(n_1637),
.B2(n_1635),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1694),
.B(n_1676),
.Y(n_1719)
);

INVx1_ASAP7_75t_SL g1720 ( 
.A(n_1681),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1697),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1681),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1695),
.A2(n_1635),
.B1(n_1637),
.B2(n_1647),
.C(n_1643),
.Y(n_1723)
);

O2A1O1Ixp5_ASAP7_75t_L g1724 ( 
.A1(n_1697),
.A2(n_1691),
.B(n_1682),
.C(n_1679),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1705),
.B(n_1643),
.Y(n_1725)
);

O2A1O1Ixp33_ASAP7_75t_L g1726 ( 
.A1(n_1697),
.A2(n_1629),
.B(n_1652),
.C(n_1647),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1693),
.B(n_1652),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1682),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1688),
.B(n_1660),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1677),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1677),
.Y(n_1731)
);

NOR2xp33_ASAP7_75t_L g1732 ( 
.A(n_1699),
.B(n_1508),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1696),
.B(n_1704),
.Y(n_1733)
);

NAND2xp33_ASAP7_75t_L g1734 ( 
.A(n_1679),
.B(n_1487),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1685),
.Y(n_1735)
);

NAND4xp25_ASAP7_75t_L g1736 ( 
.A(n_1707),
.B(n_1704),
.C(n_1706),
.D(n_1708),
.Y(n_1736)
);

OAI222xp33_ASAP7_75t_L g1737 ( 
.A1(n_1707),
.A2(n_1646),
.B1(n_1659),
.B2(n_1617),
.C1(n_1665),
.C2(n_1624),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1730),
.Y(n_1738)
);

NAND2xp33_ASAP7_75t_L g1739 ( 
.A(n_1720),
.B(n_1706),
.Y(n_1739)
);

INVxp33_ASAP7_75t_L g1740 ( 
.A(n_1732),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1723),
.A2(n_1690),
.B1(n_1692),
.B2(n_1686),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1734),
.A2(n_1690),
.B1(n_1692),
.B2(n_1686),
.Y(n_1742)
);

XNOR2xp5_ASAP7_75t_L g1743 ( 
.A(n_1718),
.B(n_1494),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1731),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1724),
.A2(n_1689),
.B(n_1710),
.Y(n_1745)
);

OAI22xp33_ASAP7_75t_SL g1746 ( 
.A1(n_1725),
.A2(n_1665),
.B1(n_1659),
.B2(n_1708),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1735),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1735),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1722),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_SL g1751 ( 
.A1(n_1716),
.A2(n_1617),
.B1(n_1624),
.B2(n_1625),
.Y(n_1751)
);

OAI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1736),
.A2(n_1620),
.B1(n_1559),
.B2(n_1685),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1714),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1714),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1728),
.Y(n_1755)
);

OAI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1740),
.A2(n_1715),
.B(n_1712),
.Y(n_1756)
);

NOR2xp33_ASAP7_75t_L g1757 ( 
.A(n_1749),
.B(n_1734),
.Y(n_1757)
);

OAI321xp33_ASAP7_75t_L g1758 ( 
.A1(n_1752),
.A2(n_1726),
.A3(n_1721),
.B1(n_1733),
.B2(n_1727),
.C(n_1719),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1753),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1754),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1747),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1755),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1739),
.B(n_1732),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1748),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1738),
.Y(n_1765)
);

AOI321xp33_ASAP7_75t_L g1766 ( 
.A1(n_1758),
.A2(n_1746),
.A3(n_1750),
.B1(n_1752),
.B2(n_1741),
.C(n_1742),
.Y(n_1766)
);

NAND4xp25_ASAP7_75t_L g1767 ( 
.A(n_1757),
.B(n_1745),
.C(n_1744),
.D(n_1751),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_L g1768 ( 
.A(n_1756),
.B(n_1728),
.C(n_1737),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1763),
.B(n_1757),
.C(n_1764),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1760),
.A2(n_1751),
.B1(n_1716),
.B2(n_1743),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1759),
.B(n_1716),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1729),
.Y(n_1772)
);

NAND4xp25_ASAP7_75t_L g1773 ( 
.A(n_1761),
.B(n_1765),
.C(n_1721),
.D(n_1717),
.Y(n_1773)
);

OAI321xp33_ASAP7_75t_L g1774 ( 
.A1(n_1761),
.A2(n_1687),
.A3(n_1683),
.B1(n_1684),
.B2(n_1680),
.C(n_1689),
.Y(n_1774)
);

OAI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1766),
.A2(n_1687),
.B(n_1710),
.C(n_1701),
.Y(n_1775)
);

AOI211xp5_ASAP7_75t_L g1776 ( 
.A1(n_1767),
.A2(n_1701),
.B(n_1684),
.C(n_1683),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1770),
.A2(n_1680),
.B(n_1703),
.Y(n_1777)
);

NAND2xp33_ASAP7_75t_R g1778 ( 
.A(n_1771),
.B(n_1711),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_SL g1779 ( 
.A1(n_1774),
.A2(n_1489),
.B(n_1670),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1775),
.A2(n_1768),
.B(n_1769),
.C(n_1773),
.Y(n_1780)
);

AOI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1776),
.A2(n_1772),
.B(n_1493),
.C(n_1711),
.Y(n_1781)
);

OAI221xp5_ASAP7_75t_SL g1782 ( 
.A1(n_1777),
.A2(n_1617),
.B1(n_1613),
.B2(n_1628),
.C(n_1625),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1778),
.A2(n_1613),
.B1(n_1668),
.B2(n_1625),
.Y(n_1783)
);

OAI211xp5_ASAP7_75t_L g1784 ( 
.A1(n_1779),
.A2(n_1533),
.B(n_1628),
.C(n_1480),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1778),
.Y(n_1785)
);

NAND4xp75_ASAP7_75t_L g1786 ( 
.A(n_1785),
.B(n_1628),
.C(n_1633),
.D(n_1611),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1780),
.B(n_1611),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1781),
.B(n_1612),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1783),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1784),
.Y(n_1790)
);

AOI222xp33_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1782),
.B1(n_1633),
.B2(n_1631),
.C1(n_1612),
.C2(n_1634),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1788),
.B(n_1604),
.Y(n_1792)
);

NOR2x1_ASAP7_75t_L g1793 ( 
.A(n_1789),
.B(n_1631),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1793),
.B(n_1790),
.Y(n_1794)
);

OA22x2_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1792),
.B1(n_1787),
.B2(n_1786),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1795),
.B(n_1791),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1795),
.Y(n_1797)
);

NOR3x1_ASAP7_75t_L g1798 ( 
.A(n_1796),
.B(n_1435),
.C(n_1431),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1797),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1604),
.B(n_1626),
.Y(n_1800)
);

OAI21x1_ASAP7_75t_SL g1801 ( 
.A1(n_1798),
.A2(n_1490),
.B(n_1483),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1800),
.Y(n_1802)
);

AOI31xp33_ASAP7_75t_L g1803 ( 
.A1(n_1802),
.A2(n_1801),
.A3(n_1444),
.B(n_1435),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1803),
.Y(n_1804)
);

AOI221xp5_ASAP7_75t_L g1805 ( 
.A1(n_1804),
.A2(n_1604),
.B1(n_1622),
.B2(n_1626),
.C(n_1621),
.Y(n_1805)
);

AOI211xp5_ASAP7_75t_L g1806 ( 
.A1(n_1805),
.A2(n_1431),
.B(n_1478),
.C(n_1604),
.Y(n_1806)
);


endmodule