module real_aes_18173_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_87;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_0), .A2(n_3), .B1(n_244), .B2(n_245), .Y(n_243) );
INVx1_ASAP7_75t_L g540 ( .A(n_1), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_2), .A2(n_16), .B1(n_171), .B2(n_180), .Y(n_188) );
AND2x2_ASAP7_75t_L g464 ( .A(n_4), .B(n_65), .Y(n_464) );
INVx1_ASAP7_75t_L g497 ( .A(n_4), .Y(n_497) );
AND2x2_ASAP7_75t_L g515 ( .A(n_4), .B(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g131 ( .A1(n_5), .A2(n_42), .B1(n_91), .B2(n_132), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_6), .A2(n_10), .B1(n_110), .B2(n_111), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_7), .Y(n_179) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_8), .Y(n_93) );
INVx1_ASAP7_75t_L g649 ( .A(n_9), .Y(n_649) );
INVx1_ASAP7_75t_L g472 ( .A(n_11), .Y(n_472) );
INVx1_ASAP7_75t_L g555 ( .A(n_11), .Y(n_555) );
INVx2_ASAP7_75t_L g478 ( .A(n_12), .Y(n_478) );
INVx1_ASAP7_75t_L g537 ( .A(n_13), .Y(n_537) );
OAI322xp33_ASAP7_75t_L g547 ( .A1(n_13), .A2(n_548), .A3(n_562), .B1(n_566), .B2(n_576), .C1(n_592), .C2(n_600), .Y(n_547) );
OAI21x1_ASAP7_75t_L g119 ( .A1(n_14), .A2(n_40), .B(n_120), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_15), .Y(n_193) );
AOI221xp5_ASAP7_75t_L g522 ( .A1(n_17), .A2(n_48), .B1(n_523), .B2(n_524), .C(n_528), .Y(n_522) );
INVx1_ASAP7_75t_L g573 ( .A(n_17), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_18), .B(n_95), .Y(n_200) );
INVx4_ASAP7_75t_R g154 ( .A(n_19), .Y(n_154) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_19), .A2(n_154), .B1(n_646), .B2(n_647), .Y(n_645) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_20), .B(n_171), .Y(n_206) );
INVx1_ASAP7_75t_L g249 ( .A(n_21), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_SL g177 ( .A1(n_22), .A2(n_94), .B(n_110), .C(n_178), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_23), .A2(n_37), .B1(n_110), .B2(n_114), .Y(n_189) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_24), .A2(n_652), .B1(n_653), .B2(n_654), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g653 ( .A(n_24), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_25), .A2(n_34), .B1(n_499), .B2(n_504), .Y(n_498) );
INVxp33_ASAP7_75t_L g567 ( .A(n_25), .Y(n_567) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_26), .Y(n_174) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_27), .A2(n_28), .B1(n_499), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g583 ( .A(n_27), .Y(n_583) );
INVxp67_ASAP7_75t_L g557 ( .A(n_28), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_29), .A2(n_454), .B1(n_657), .B2(n_677), .Y(n_676) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_29), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_30), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g565 ( .A(n_30), .Y(n_565) );
INVx1_ASAP7_75t_L g599 ( .A(n_30), .Y(n_599) );
INVx1_ASAP7_75t_L g203 ( .A(n_31), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_32), .B(n_110), .Y(n_205) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_33), .A2(n_50), .B1(n_483), .B2(n_487), .C(n_493), .Y(n_482) );
INVxp67_ASAP7_75t_L g580 ( .A(n_33), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_34), .A2(n_48), .B1(n_585), .B2(n_589), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_35), .Y(n_222) );
INVx2_ASAP7_75t_L g666 ( .A(n_36), .Y(n_666) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_38), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_39), .A2(n_68), .B1(n_110), .B2(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g511 ( .A(n_41), .Y(n_511) );
BUFx3_ASAP7_75t_L g474 ( .A(n_43), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_44), .Y(n_122) );
AND2x4_ASAP7_75t_L g85 ( .A(n_45), .B(n_86), .Y(n_85) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_45), .Y(n_675) );
INVx1_ASAP7_75t_L g120 ( .A(n_46), .Y(n_120) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_47), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_49), .A2(n_71), .B1(n_114), .B2(n_242), .Y(n_241) );
INVxp67_ASAP7_75t_L g549 ( .A(n_50), .Y(n_549) );
AO22x1_ASAP7_75t_L g135 ( .A1(n_51), .A2(n_58), .B1(n_136), .B2(n_138), .Y(n_135) );
INVx1_ASAP7_75t_L g86 ( .A(n_52), .Y(n_86) );
AND2x2_ASAP7_75t_L g181 ( .A(n_53), .B(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g521 ( .A(n_54), .Y(n_521) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_55), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_56), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_57), .B(n_132), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_59), .B(n_171), .Y(n_223) );
INVx1_ASAP7_75t_L g691 ( .A(n_59), .Y(n_691) );
INVx2_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_61), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_62), .B(n_182), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_63), .B(n_118), .Y(n_133) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_64), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g643 ( .A(n_64), .Y(n_643) );
BUFx3_ASAP7_75t_L g496 ( .A(n_65), .Y(n_496) );
INVx1_ASAP7_75t_L g516 ( .A(n_65), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g617 ( .A(n_66), .Y(n_617) );
INVx1_ASAP7_75t_L g517 ( .A(n_67), .Y(n_517) );
OAI211xp5_ASAP7_75t_L g618 ( .A1(n_67), .A2(n_619), .B(n_624), .C(n_635), .Y(n_618) );
INVx1_ASAP7_75t_L g467 ( .A(n_69), .Y(n_467) );
INVx2_ASAP7_75t_L g546 ( .A(n_69), .Y(n_546) );
INVx1_ASAP7_75t_L g598 ( .A(n_69), .Y(n_598) );
BUFx2_ASAP7_75t_L g652 ( .A(n_70), .Y(n_652) );
BUFx2_ASAP7_75t_L g647 ( .A(n_71), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_72), .B(n_182), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_73), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_74), .A2(n_116), .B(n_132), .C(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g158 ( .A(n_75), .B(n_159), .Y(n_158) );
BUFx2_ASAP7_75t_L g642 ( .A(n_76), .Y(n_642) );
NAND2xp33_ASAP7_75t_L g227 ( .A(n_77), .B(n_155), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_96), .B(n_452), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_83), .B(n_87), .Y(n_82) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_83), .A2(n_149), .B(n_152), .Y(n_148) );
INVx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
AO31x2_ASAP7_75t_L g107 ( .A1(n_84), .A2(n_108), .A3(n_117), .B(n_121), .Y(n_107) );
BUFx10_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
BUFx10_ASAP7_75t_L g191 ( .A(n_85), .Y(n_191) );
INVx1_ASAP7_75t_L g247 ( .A(n_85), .Y(n_247) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_86), .Y(n_673) );
AOI21xp5_ASAP7_75t_SL g693 ( .A1(n_87), .A2(n_681), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g87 ( .A(n_88), .B(n_94), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_92), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx3_ASAP7_75t_L g110 ( .A(n_93), .Y(n_110) );
BUFx6f_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
INVx1_ASAP7_75t_L g132 ( .A(n_93), .Y(n_132) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_93), .Y(n_137) );
INVx1_ASAP7_75t_L g139 ( .A(n_93), .Y(n_139) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_93), .Y(n_156) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_93), .Y(n_171) );
INVx1_ASAP7_75t_L g173 ( .A(n_93), .Y(n_173) );
INVx2_ASAP7_75t_L g180 ( .A(n_93), .Y(n_180) );
INVx6_ASAP7_75t_L g112 ( .A(n_94), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_94), .B(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_94), .A2(n_227), .B(n_228), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_94), .A2(n_127), .B(n_135), .C(n_141), .Y(n_270) );
BUFx8_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g116 ( .A(n_95), .Y(n_116) );
INVx2_ASAP7_75t_L g130 ( .A(n_95), .Y(n_130) );
INVx1_ASAP7_75t_L g176 ( .A(n_95), .Y(n_176) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
NOR2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_366), .Y(n_98) );
NAND4xp75_ASAP7_75t_L g99 ( .A(n_100), .B(n_271), .C(n_313), .D(n_337), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI211xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_160), .B(n_208), .C(n_250), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g357 ( .A(n_104), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g451 ( .A(n_104), .B(n_388), .Y(n_451) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_124), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_L g266 ( .A(n_106), .B(n_218), .Y(n_266) );
AND2x2_ASAP7_75t_L g307 ( .A(n_106), .B(n_268), .Y(n_307) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g214 ( .A(n_107), .B(n_144), .Y(n_214) );
OR2x2_ASAP7_75t_L g232 ( .A(n_107), .B(n_144), .Y(n_232) );
INVx2_ASAP7_75t_L g258 ( .A(n_107), .Y(n_258) );
AND2x2_ASAP7_75t_L g288 ( .A(n_107), .B(n_218), .Y(n_288) );
AND2x2_ASAP7_75t_L g317 ( .A(n_107), .B(n_143), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_107), .B(n_269), .Y(n_353) );
OAI22x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_112), .B1(n_113), .B2(n_115), .Y(n_108) );
INVx4_ASAP7_75t_L g111 ( .A(n_110), .Y(n_111) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_111), .A2(n_222), .B(n_223), .C(n_224), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g187 ( .A1(n_112), .A2(n_128), .B1(n_188), .B2(n_189), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_112), .A2(n_115), .B1(n_241), .B2(n_243), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_114), .B(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g244 ( .A(n_114), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_115), .B(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g123 ( .A(n_118), .Y(n_123) );
OAI21xp33_ASAP7_75t_L g141 ( .A1(n_118), .A2(n_133), .B(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g147 ( .A(n_118), .Y(n_147) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_119), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx2_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
BUFx2_ASAP7_75t_L g166 ( .A(n_123), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_123), .B(n_193), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_123), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g330 ( .A(n_124), .B(n_259), .Y(n_330) );
INVx2_ASAP7_75t_L g425 ( .A(n_124), .Y(n_425) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_143), .Y(n_124) );
INVx2_ASAP7_75t_L g213 ( .A(n_125), .Y(n_213) );
AND2x4_ASAP7_75t_L g256 ( .A(n_125), .B(n_144), .Y(n_256) );
AOI21x1_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_134), .B(n_140), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI21x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B(n_133), .Y(n_127) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_128), .A2(n_205), .B(n_206), .Y(n_204) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g225 ( .A(n_130), .Y(n_225) );
INVxp67_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
OAI21xp33_ASAP7_75t_SL g199 ( .A1(n_138), .A2(n_200), .B(n_201), .Y(n_199) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_142), .A2(n_168), .B(n_177), .Y(n_167) );
AND2x2_ASAP7_75t_L g415 ( .A(n_143), .B(n_213), .Y(n_415) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g279 ( .A(n_144), .Y(n_279) );
AND2x2_ASAP7_75t_L g336 ( .A(n_144), .B(n_218), .Y(n_336) );
AND2x2_ASAP7_75t_L g351 ( .A(n_144), .B(n_259), .Y(n_351) );
AND2x2_ASAP7_75t_L g373 ( .A(n_144), .B(n_213), .Y(n_373) );
AO21x2_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_148), .B(n_158), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI22xp33_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B1(n_156), .B2(n_157), .Y(n_153) );
INVx2_ASAP7_75t_L g242 ( .A(n_155), .Y(n_242) );
OAI211xp5_ASAP7_75t_SL g420 ( .A1(n_160), .A2(n_421), .B(n_423), .C(n_430), .Y(n_420) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_194), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OR2x2_ASAP7_75t_L g407 ( .A(n_163), .B(n_343), .Y(n_407) );
OR2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_184), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_164), .B(n_196), .Y(n_306) );
INVxp67_ASAP7_75t_L g320 ( .A(n_164), .Y(n_320) );
AND2x2_ASAP7_75t_L g340 ( .A(n_164), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_164), .B(n_253), .Y(n_347) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g236 ( .A(n_165), .Y(n_236) );
AOI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_181), .Y(n_165) );
AO31x2_ASAP7_75t_L g239 ( .A1(n_166), .A2(n_240), .A3(n_246), .B(n_248), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_172), .B(n_175), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx2_ASAP7_75t_L g245 ( .A(n_173), .Y(n_245) );
BUFx4f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_176), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx2_ASAP7_75t_L g190 ( .A(n_182), .Y(n_190) );
NOR2x1_ASAP7_75t_L g229 ( .A(n_182), .B(n_230), .Y(n_229) );
INVx4_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g207 ( .A(n_183), .B(n_191), .Y(n_207) );
OR2x2_ASAP7_75t_L g281 ( .A(n_184), .B(n_263), .Y(n_281) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
OR2x2_ASAP7_75t_L g329 ( .A(n_185), .B(n_236), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_185), .B(n_239), .Y(n_335) );
INVx2_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g235 ( .A(n_186), .B(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g304 ( .A(n_186), .B(n_239), .Y(n_304) );
BUFx2_ASAP7_75t_L g311 ( .A(n_186), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_186), .B(n_239), .Y(n_391) );
AO31x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_190), .A3(n_191), .B(n_192), .Y(n_186) );
INVx1_ASAP7_75t_L g230 ( .A(n_191), .Y(n_230) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x4_ASAP7_75t_L g321 ( .A(n_195), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g450 ( .A(n_195), .B(n_235), .Y(n_450) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx3_ASAP7_75t_L g253 ( .A(n_196), .Y(n_253) );
AND2x2_ASAP7_75t_L g264 ( .A(n_196), .B(n_239), .Y(n_264) );
AND2x2_ASAP7_75t_L g310 ( .A(n_196), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g343 ( .A(n_196), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_196), .B(n_254), .Y(n_360) );
AND2x2_ASAP7_75t_L g399 ( .A(n_196), .B(n_400), .Y(n_399) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_204), .B(n_207), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_215), .B(n_233), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_210), .A2(n_378), .B1(n_379), .B2(n_381), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_214), .Y(n_210) );
AND2x2_ASAP7_75t_L g375 ( .A(n_211), .B(n_266), .Y(n_375) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g290 ( .A(n_212), .Y(n_290) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g439 ( .A(n_213), .B(n_259), .Y(n_439) );
AND2x2_ASAP7_75t_L g403 ( .A(n_214), .B(n_298), .Y(n_403) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_231), .Y(n_215) );
OR2x2_ASAP7_75t_L g300 ( .A(n_216), .B(n_277), .Y(n_300) );
OR2x2_ASAP7_75t_L g412 ( .A(n_216), .B(n_232), .Y(n_412) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
BUFx3_ASAP7_75t_L g341 ( .A(n_218), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
OAI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_226), .B(n_229), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_222), .A2(n_454), .B1(n_657), .B2(n_689), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_222), .Y(n_689) );
INVx2_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
OR2x2_ASAP7_75t_L g409 ( .A(n_232), .B(n_268), .Y(n_409) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_237), .Y(n_234) );
AND2x2_ASAP7_75t_L g251 ( .A(n_235), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g292 ( .A(n_235), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g429 ( .A(n_235), .Y(n_429) );
INVx1_ASAP7_75t_L g448 ( .A(n_235), .Y(n_448) );
INVx2_ASAP7_75t_L g263 ( .A(n_236), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_236), .B(n_239), .Y(n_312) );
INVx1_ASAP7_75t_L g376 ( .A(n_237), .Y(n_376) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g437 ( .A(n_238), .Y(n_437) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g254 ( .A(n_239), .Y(n_254) );
INVx1_ASAP7_75t_L g344 ( .A(n_239), .Y(n_344) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_255), .B1(n_260), .B2(n_265), .Y(n_250) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx2_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
AND2x2_ASAP7_75t_L g295 ( .A(n_253), .B(n_280), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_253), .B(n_263), .Y(n_355) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx3_ASAP7_75t_L g286 ( .A(n_256), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_256), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g380 ( .A(n_256), .B(n_364), .Y(n_380) );
INVx1_ASAP7_75t_L g284 ( .A(n_257), .Y(n_284) );
AOI222xp33_ASAP7_75t_L g294 ( .A1(n_257), .A2(n_295), .B1(n_296), .B2(n_301), .C1(n_307), .C2(n_308), .Y(n_294) );
OAI21xp33_ASAP7_75t_SL g324 ( .A1(n_257), .A2(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g348 ( .A(n_257), .B(n_267), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_257), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OR2x2_ASAP7_75t_L g277 ( .A(n_258), .B(n_269), .Y(n_277) );
INVx1_ASAP7_75t_L g365 ( .A(n_258), .Y(n_365) );
BUFx2_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_262), .B(n_303), .Y(n_332) );
OR2x2_ASAP7_75t_L g444 ( .A(n_262), .B(n_304), .Y(n_444) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g327 ( .A(n_264), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g442 ( .A(n_264), .Y(n_442) );
OAI31xp33_ASAP7_75t_L g423 ( .A1(n_265), .A2(n_424), .A3(n_426), .B(n_427), .Y(n_423) );
AND2x4_ASAP7_75t_SL g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_266), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_294), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_280), .B(n_282), .Y(n_272) );
NOR2x1_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x6_ASAP7_75t_L g393 ( .A(n_275), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g325 ( .A(n_278), .Y(n_325) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g416 ( .A(n_279), .B(n_353), .Y(n_416) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_281), .A2(n_370), .B1(n_372), .B2(n_374), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g430 ( .A1(n_281), .A2(n_342), .B(n_404), .C(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B(n_291), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND4xp25_ASAP7_75t_L g383 ( .A(n_286), .B(n_384), .C(n_385), .D(n_387), .Y(n_383) );
NAND2x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_288), .B(n_290), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_288), .B(n_373), .Y(n_396) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g362 ( .A(n_293), .B(n_322), .Y(n_362) );
NAND2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_300), .Y(n_296) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_300), .A2(n_444), .B1(n_445), .B2(n_447), .Y(n_443) );
AOI221x1_ASAP7_75t_L g382 ( .A1(n_301), .A2(n_383), .B1(n_389), .B2(n_392), .C(n_395), .Y(n_382) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g322 ( .A(n_304), .Y(n_322) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g334 ( .A(n_306), .B(n_335), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g397 ( .A(n_307), .B(n_388), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_L g410 ( .A1(n_308), .A2(n_392), .B(n_411), .C(n_413), .Y(n_410) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx2_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_323), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_315), .A2(n_333), .B1(n_403), .B2(n_404), .C(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g339 ( .A(n_317), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_317), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g438 ( .A(n_317), .B(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2x1_ASAP7_75t_L g417 ( .A(n_320), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g441 ( .A(n_320), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g381 ( .A(n_321), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B1(n_330), .B2(n_331), .C1(n_333), .C2(n_336), .Y(n_323) );
INVx1_ASAP7_75t_L g408 ( .A(n_327), .Y(n_408) );
INVx1_ASAP7_75t_L g371 ( .A(n_328), .Y(n_371) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g405 ( .A(n_329), .Y(n_405) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g346 ( .A(n_335), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g400 ( .A(n_335), .Y(n_400) );
AND2x2_ASAP7_75t_L g363 ( .A(n_336), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_356), .Y(n_337) );
AOI222xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_342), .B1(n_345), .B2(n_348), .C1(n_349), .C2(n_354), .Y(n_338) );
INVx3_ASAP7_75t_L g388 ( .A(n_341), .Y(n_388) );
BUFx2_ASAP7_75t_L g446 ( .A(n_341), .Y(n_446) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g418 ( .A(n_343), .Y(n_418) );
OR2x2_ASAP7_75t_L g428 ( .A(n_343), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
INVx2_ASAP7_75t_SL g386 ( .A(n_351), .Y(n_386) );
AND2x2_ASAP7_75t_L g431 ( .A(n_352), .B(n_388), .Y(n_431) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
INVxp67_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g390 ( .A(n_355), .B(n_391), .Y(n_390) );
NOR2x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_361), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
OR2x2_ASAP7_75t_L g447 ( .A(n_360), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
INVx1_ASAP7_75t_L g378 ( .A(n_362), .Y(n_378) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x2_ASAP7_75t_L g385 ( .A(n_365), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g435 ( .A(n_365), .Y(n_435) );
NAND4xp75_ASAP7_75t_L g366 ( .A(n_367), .B(n_401), .C(n_419), .D(n_432), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_382), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_369), .A2(n_376), .B(n_377), .Y(n_368) );
INVxp33_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_371), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
AND2x2_ASAP7_75t_L g434 ( .A(n_373), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g404 ( .A(n_376), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OAI22xp33_ASAP7_75t_SL g413 ( .A1(n_390), .A2(n_414), .B1(n_416), .B2(n_417), .Y(n_413) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI21xp33_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g426 ( .A(n_397), .Y(n_426) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_410), .Y(n_401) );
AOI21xp5_ASAP7_75t_SL g406 ( .A1(n_407), .A2(n_408), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx3_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_449), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_438), .B2(n_440), .C(n_443), .Y(n_433) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
OAI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_659), .B1(n_676), .B2(n_678), .C(n_682), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_638), .B1(n_657), .B2(n_658), .Y(n_453) );
INVx1_ASAP7_75t_L g657 ( .A(n_454), .Y(n_657) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_604), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_479), .B1(n_480), .B2(n_541), .C(n_547), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_468), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_465), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_464), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g485 ( .A(n_463), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g491 ( .A(n_463), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g502 ( .A(n_463), .Y(n_502) );
INVx2_ASAP7_75t_L g507 ( .A(n_463), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_464), .B(n_509), .Y(n_508) );
AND2x6_ASAP7_75t_L g533 ( .A(n_464), .B(n_484), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_464), .B(n_501), .Y(n_616) );
INVxp67_ASAP7_75t_L g610 ( .A(n_465), .Y(n_610) );
BUFx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g476 ( .A(n_466), .Y(n_476) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx3_ASAP7_75t_L g575 ( .A(n_469), .Y(n_575) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_472), .B(n_474), .Y(n_561) );
INVx2_ASAP7_75t_L g591 ( .A(n_472), .Y(n_591) );
INVx2_ASAP7_75t_L g628 ( .A(n_473), .Y(n_628) );
BUFx6f_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g556 ( .A(n_474), .Y(n_556) );
OR2x2_ASAP7_75t_L g571 ( .A(n_474), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_L g590 ( .A(n_474), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g602 ( .A(n_475), .Y(n_602) );
OR2x2_ASAP7_75t_L g613 ( .A(n_475), .B(n_559), .Y(n_613) );
INVx1_ASAP7_75t_L g623 ( .A(n_475), .Y(n_623) );
OR2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
OR2x2_ASAP7_75t_L g563 ( .A(n_476), .B(n_564), .Y(n_563) );
NAND2xp33_ASAP7_75t_SL g564 ( .A(n_478), .B(n_565), .Y(n_564) );
INVx3_ASAP7_75t_L g596 ( .A(n_478), .Y(n_596) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_518), .C(n_534), .Y(n_480) );
AOI222xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_498), .B1(n_508), .B2(n_511), .C1(n_512), .C2(n_517), .Y(n_481) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x4_ASAP7_75t_SL g520 ( .A(n_484), .B(n_515), .Y(n_520) );
BUFx3_ASAP7_75t_L g523 ( .A(n_484), .Y(n_523) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g492 ( .A(n_486), .Y(n_492) );
INVx1_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
AND2x2_ASAP7_75t_L g506 ( .A(n_486), .B(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g510 ( .A(n_486), .Y(n_510) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g536 ( .A(n_490), .B(n_515), .Y(n_536) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g527 ( .A(n_491), .Y(n_527) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g530 ( .A(n_496), .B(n_497), .Y(n_530) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g514 ( .A(n_501), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_505), .Y(n_532) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_506), .Y(n_539) );
BUFx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_511), .A2(n_521), .B1(n_625), .B2(n_630), .Y(n_624) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_L g538 ( .A(n_515), .B(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_521), .B1(n_522), .B2(n_531), .C(n_533), .Y(n_518) );
BUFx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
HB1xp67_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_537), .B1(n_538), .B2(n_540), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_540), .A2(n_605), .B1(n_611), .B2(n_617), .C(n_618), .Y(n_604) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_550), .B1(n_557), .B2(n_558), .Y(n_548) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_553), .Y(n_579) );
BUFx8_ASAP7_75t_L g603 ( .A(n_553), .Y(n_603) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g572 ( .A(n_555), .Y(n_572) );
AND2x4_ASAP7_75t_L g587 ( .A(n_556), .B(n_588), .Y(n_587) );
BUFx3_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g582 ( .A(n_561), .Y(n_582) );
BUFx8_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g671 ( .A(n_564), .Y(n_671) );
INVx1_ASAP7_75t_L g609 ( .A(n_565), .Y(n_609) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B1(n_573), .B2(n_574), .Y(n_566) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx4f_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g621 ( .A(n_571), .Y(n_621) );
INVx1_ASAP7_75t_L g588 ( .A(n_572), .Y(n_588) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B1(n_581), .B2(n_583), .C(n_584), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
BUFx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx8_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx8_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_587), .B(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
BUFx2_ASAP7_75t_L g637 ( .A(n_590), .Y(n_637) );
INVx1_ASAP7_75t_L g634 ( .A(n_591), .Y(n_634) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NAND3x1_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .C(n_599), .Y(n_595) );
AND2x4_ASAP7_75t_L g608 ( .A(n_596), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g615 ( .A(n_598), .Y(n_615) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_603), .Y(n_601) );
INVx3_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x6_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
AND2x4_ASAP7_75t_L g629 ( .A(n_608), .B(n_615), .Y(n_629) );
AND2x6_ASAP7_75t_L g665 ( .A(n_608), .B(n_627), .Y(n_665) );
INVx8_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
OR2x6_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
INVx2_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2x1_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND3xp33_ASAP7_75t_L g667 ( .A(n_627), .B(n_668), .C(n_671), .Y(n_667) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x4_ASAP7_75t_L g630 ( .A(n_629), .B(n_631), .Y(n_630) );
AND2x4_ASAP7_75t_L g636 ( .A(n_629), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
CKINVDCx14_ASAP7_75t_R g658 ( .A(n_638), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B1(n_648), .B2(n_656), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
XOR2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_645), .Y(n_640) );
INVx1_ASAP7_75t_L g644 ( .A(n_642), .Y(n_644) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g656 ( .A(n_648), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_651), .B2(n_655), .Y(n_648) );
INVx1_ASAP7_75t_SL g655 ( .A(n_649), .Y(n_655) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g654 ( .A(n_652), .Y(n_654) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx3_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx12f_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
BUFx8_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_667), .C(n_672), .Y(n_663) );
AND2x2_ASAP7_75t_L g687 ( .A(n_664), .B(n_667), .Y(n_687) );
INVx4_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g670 ( .A(n_666), .Y(n_670) );
INVx2_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g686 ( .A(n_672), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
BUFx2_ASAP7_75t_L g681 ( .A(n_673), .Y(n_681) );
AND2x2_ASAP7_75t_L g694 ( .A(n_673), .B(n_674), .Y(n_694) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g680 ( .A(n_675), .B(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx4f_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_688), .B1(n_690), .B2(n_692), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OR2x6_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx2_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
endmodule