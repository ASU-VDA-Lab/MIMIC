module fake_netlist_6_2596_n_202 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_202);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_202;

wire n_52;
wire n_119;
wire n_146;
wire n_46;
wire n_91;
wire n_163;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_199;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_195;
wire n_189;
wire n_32;
wire n_85;
wire n_66;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_197;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_196;
wire n_200;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_198;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_201;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

OR2x6_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_2),
.Y(n_67)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx5p33_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_46),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_70),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_54),
.A2(n_52),
.B1(n_49),
.B2(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_49),
.Y(n_87)
);

NAND2x1p5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_47),
.Y(n_88)
);

NAND2xp33_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_45),
.Y(n_89)
);

NOR2xp67_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_18),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_74),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_56),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_61),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_58),
.B(n_60),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_63),
.B1(n_67),
.B2(n_72),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_89),
.A2(n_73),
.B(n_45),
.C(n_34),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_74),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_67),
.Y(n_103)
);

OAI21x1_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_88),
.B(n_87),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

AO31x2_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_34),
.A3(n_102),
.B(n_79),
.Y(n_107)
);

OAI21x1_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_88),
.B(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_110),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_100),
.B(n_94),
.C(n_103),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_83),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_105),
.Y(n_117)
);

CKINVDCx11_ASAP7_75t_R g118 ( 
.A(n_106),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_108),
.B(n_104),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_99),
.B1(n_85),
.B2(n_83),
.C(n_77),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_122),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_116),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_116),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NOR2x1p5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_59),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_124),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_113),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_107),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_130),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_114),
.B(n_131),
.C(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_137),
.B(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_127),
.B1(n_134),
.B2(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_130),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_127),
.B(n_90),
.C(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_143),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_140),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_138),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_107),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_SL g161 ( 
.A(n_145),
.B(n_131),
.Y(n_161)
);

OAI221xp5_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_150),
.B1(n_81),
.B2(n_91),
.C(n_132),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_134),
.B1(n_144),
.B2(n_152),
.Y(n_163)
);

OAI221xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_91),
.B1(n_81),
.B2(n_62),
.C(n_88),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_153),
.A2(n_83),
.B(n_85),
.Y(n_165)
);

NAND4xp25_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_98),
.C(n_79),
.D(n_76),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_129),
.Y(n_167)
);

AOI222xp33_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_85),
.B1(n_133),
.B2(n_125),
.C1(n_8),
.C2(n_9),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_156),
.A2(n_104),
.B(n_108),
.Y(n_169)
);

AOI211xp5_ASAP7_75t_L g170 ( 
.A1(n_157),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_154),
.A2(n_133),
.B(n_109),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_154),
.Y(n_172)
);

NAND3x2_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_159),
.C(n_7),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_159),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_109),
.B1(n_104),
.B2(n_111),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_107),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_169),
.Y(n_177)
);

OAI321xp33_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_111),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C(n_14),
.Y(n_178)
);

NAND4xp25_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_6),
.C(n_10),
.D(n_11),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_172),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_174),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_177),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_173),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_175),
.Y(n_187)
);

AND2x4_ASAP7_75t_SL g188 ( 
.A(n_182),
.B(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_165),
.C(n_171),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_14),
.B1(n_111),
.B2(n_86),
.C(n_93),
.Y(n_192)
);

NAND4xp25_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_106),
.C(n_107),
.D(n_112),
.Y(n_193)
);

OR3x1_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_107),
.C(n_21),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_187),
.B1(n_184),
.B2(n_185),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_180),
.B1(n_106),
.B2(n_25),
.Y(n_197)
);

OR3x2_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_193),
.C(n_189),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_192),
.B(n_191),
.C(n_28),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_197),
.A2(n_19),
.B(n_24),
.C(n_30),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_199),
.B1(n_200),
.B2(n_96),
.Y(n_201)
);

NOR4xp25_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_96),
.C(n_108),
.D(n_199),
.Y(n_202)
);


endmodule