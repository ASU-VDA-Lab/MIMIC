module fake_jpeg_31321_n_62 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx16_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_2),
.Y(n_9)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_6),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_9),
.A2(n_0),
.B(n_2),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_21),
.C(n_28),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_18),
.B(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_22),
.Y(n_32)
);

OR2x2_ASAP7_75t_SL g21 ( 
.A(n_10),
.B(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_SL g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_7),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_25),
.B(n_8),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_26),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_9),
.B(n_3),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_15),
.B1(n_14),
.B2(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_35),
.B(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_16),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_37),
.B(n_40),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_21),
.C(n_28),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_35),
.C(n_11),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_43),
.B1(n_34),
.B2(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

A2O1A1O1Ixp25_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_43),
.B(n_22),
.C(n_24),
.D(n_34),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_37),
.C(n_11),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_50),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_42),
.C(n_14),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_14),
.C(n_15),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_45),
.B(n_22),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_52),
.A2(n_46),
.B1(n_29),
.B2(n_15),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_55),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_54),
.A2(n_12),
.B(n_16),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_12),
.B(n_5),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_29),
.C(n_17),
.Y(n_58)
);

BUFx24_ASAP7_75t_SL g60 ( 
.A(n_58),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_60),
.B(n_59),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_24),
.Y(n_62)
);


endmodule