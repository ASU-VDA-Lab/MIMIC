module fake_jpeg_1540_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_1),
.B(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_0),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_16),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_12),
.B(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_18),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_20),
.B1(n_21),
.B2(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_3),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_10),
.C(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_15),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_27),
.B2(n_17),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_11),
.B(n_14),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_33),
.C(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_28),
.B(n_22),
.C(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_39),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_31),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_5),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_18),
.B1(n_4),
.B2(n_5),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_18),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.C(n_46),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_40),
.Y(n_46)
);

OAI221xp5_ASAP7_75t_SL g48 ( 
.A1(n_47),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.C(n_46),
.Y(n_48)
);


endmodule