module fake_jpeg_24710_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx8_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_37),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_22),
.B1(n_35),
.B2(n_23),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_52),
.A2(n_55),
.B1(n_61),
.B2(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_23),
.B1(n_29),
.B2(n_32),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_59),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_71),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_23),
.B1(n_35),
.B2(n_22),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_19),
.B1(n_36),
.B2(n_32),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_67),
.B(n_73),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx4f_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_35),
.B1(n_22),
.B2(n_26),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_78),
.B1(n_30),
.B2(n_21),
.Y(n_113)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_38),
.B(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_43),
.B(n_19),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_33),
.B1(n_26),
.B2(n_27),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_79),
.A2(n_24),
.B1(n_20),
.B2(n_27),
.Y(n_93)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_81),
.Y(n_119)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_38),
.B(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

NAND2xp33_ASAP7_75t_SL g84 ( 
.A(n_42),
.B(n_20),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_84),
.A2(n_20),
.B(n_33),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_39),
.B(n_37),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_31),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_44),
.B1(n_26),
.B2(n_27),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_88),
.A2(n_96),
.B1(n_116),
.B2(n_111),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_36),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_105),
.Y(n_124)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_97),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_28),
.B(n_97),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_33),
.B(n_78),
.C(n_52),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_99),
.A2(n_88),
.B1(n_72),
.B2(n_62),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_46),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_120),
.Y(n_127)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_31),
.A3(n_28),
.B1(n_21),
.B2(n_42),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_42),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_79),
.B1(n_66),
.B2(n_54),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_130),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_114),
.A2(n_49),
.B1(n_72),
.B2(n_74),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_122),
.A2(n_125),
.B1(n_133),
.B2(n_143),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_74),
.B1(n_62),
.B2(n_54),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_152),
.B1(n_132),
.B2(n_123),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_49),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_66),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_138),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_101),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_42),
.C(n_46),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_120),
.C(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_140),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_40),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_40),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_148),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_28),
.B1(n_21),
.B2(n_40),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_144),
.A2(n_109),
.B(n_110),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_17),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_149),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_39),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_2),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_169),
.C(n_135),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_159),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_152),
.B(n_108),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_164),
.B(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_165),
.B(n_168),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_166),
.A2(n_144),
.B(n_143),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_39),
.C(n_68),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_176),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_107),
.B1(n_106),
.B2(n_91),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_171),
.A2(n_177),
.B1(n_126),
.B2(n_149),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_17),
.C(n_16),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_179),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_92),
.Y(n_175)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_175),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_92),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_139),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_137),
.B(n_91),
.Y(n_182)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_183),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_R g227 ( 
.A(n_184),
.B(n_158),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_132),
.B1(n_123),
.B2(n_146),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_177),
.B1(n_183),
.B2(n_158),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_187),
.A2(n_171),
.B1(n_167),
.B2(n_170),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_121),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_197),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_136),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_151),
.B(n_140),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_157),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_206),
.Y(n_220)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_205),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_153),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_213),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_190),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_167),
.B1(n_195),
.B2(n_179),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_215),
.A2(n_219),
.B(n_221),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_159),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_217),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_165),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_198),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_169),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_197),
.C(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_193),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_227),
.B1(n_160),
.B2(n_162),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_157),
.Y(n_225)
);

AOI21x1_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_160),
.B(n_156),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_226),
.A2(n_208),
.B1(n_212),
.B2(n_217),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_208),
.A2(n_186),
.B1(n_206),
.B2(n_168),
.Y(n_228)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_230),
.B(n_233),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_232),
.C(n_240),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_222),
.C(n_218),
.Y(n_232)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_188),
.A3(n_194),
.B1(n_207),
.B2(n_205),
.C1(n_185),
.C2(n_180),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_239),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_216),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_201),
.B1(n_193),
.B2(n_202),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_203),
.C(n_199),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_155),
.C(n_148),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_240),
.C(n_237),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_161),
.B(n_3),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_243),
.A2(n_2),
.B(n_4),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_248),
.Y(n_259)
);

AOI321xp33_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_225),
.A3(n_215),
.B1(n_209),
.B2(n_224),
.C(n_211),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_247),
.A2(n_241),
.B(n_239),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_211),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_254),
.C(n_10),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_9),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_223),
.B(n_6),
.C(n_7),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_242),
.B(n_8),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_223),
.C(n_107),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_257),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_5),
.C(n_7),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_233),
.B1(n_236),
.B2(n_229),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_252),
.B1(n_249),
.B2(n_248),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_260),
.A2(n_11),
.B(n_12),
.Y(n_274)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_261),
.B(n_266),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_265),
.B(n_264),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_263),
.A2(n_253),
.B1(n_262),
.B2(n_265),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_8),
.B(n_9),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_244),
.C(n_250),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_270),
.A2(n_264),
.B1(n_261),
.B2(n_269),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_272),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_260),
.A2(n_252),
.B(n_249),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_274),
.B(n_258),
.Y(n_277)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_279),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_267),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_273),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_281),
.B(n_277),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_278),
.A2(n_259),
.B(n_12),
.Y(n_281)
);

OAI321xp33_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_285),
.A3(n_286),
.B1(n_11),
.B2(n_13),
.C(n_14),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_259),
.C(n_12),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_11),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_13),
.C(n_15),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_15),
.Y(n_289)
);


endmodule