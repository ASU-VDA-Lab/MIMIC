module fake_jpeg_26894_n_49 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_49);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_49;

wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_4),
.B(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_1),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_28),
.C(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_2),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_23),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_32),
.B(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

OA21x2_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_20),
.B(n_3),
.Y(n_38)
);

AOI32xp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_20),
.A3(n_24),
.B1(n_22),
.B2(n_7),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_9),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_12),
.B1(n_15),
.B2(n_5),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_8),
.C(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_44),
.B(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_45),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_46),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_42),
.C(n_43),
.Y(n_48)
);

AOI31xp33_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_39),
.A3(n_40),
.B(n_31),
.Y(n_49)
);


endmodule