module fake_jpeg_9336_n_110 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx9p33_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_9),
.C(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_23),
.B(n_25),
.Y(n_36)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_26),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_12),
.B(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_13),
.B1(n_16),
.B2(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_29),
.A2(n_37),
.B1(n_27),
.B2(n_21),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_20),
.B1(n_17),
.B2(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_17),
.B1(n_20),
.B2(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_22),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_26),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_40),
.B(n_42),
.Y(n_65)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_49),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_30),
.B1(n_20),
.B2(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_25),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_3),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_55),
.Y(n_70)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_29),
.B(n_37),
.C(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_61),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_53),
.B(n_39),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_54),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_62),
.A2(n_44),
.B(n_39),
.C(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_70),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_4),
.Y(n_67)
);

NOR2xp67_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_9),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_4),
.C(n_5),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_43),
.C(n_6),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_76),
.B(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND3xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_47),
.C(n_44),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_68),
.C(n_65),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_41),
.B1(n_51),
.B2(n_5),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_62),
.B1(n_60),
.B2(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_88),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_66),
.B1(n_57),
.B2(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_89),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_83),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_90),
.B(n_93),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_85),
.B(n_79),
.C(n_87),
.D(n_89),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_84),
.B(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_58),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_98),
.B(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_5),
.Y(n_105)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_92),
.A3(n_94),
.B1(n_95),
.B2(n_67),
.C1(n_83),
.C2(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_102),
.A2(n_103),
.B1(n_74),
.B2(n_77),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_74),
.A3(n_61),
.B1(n_82),
.B2(n_58),
.C1(n_65),
.C2(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_105),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_64),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_64),
.C(n_7),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_7),
.B(n_106),
.C(n_64),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_107),
.Y(n_110)
);


endmodule