module real_aes_18428_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_884;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AND2x4_ASAP7_75t_L g883 ( .A(n_0), .B(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_1), .A2(n_34), .B1(n_144), .B2(n_156), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_2), .A2(n_9), .B1(n_549), .B2(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g884 ( .A(n_3), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_4), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_5), .A2(n_10), .B1(n_559), .B2(n_560), .Y(n_558) );
OR2x2_ASAP7_75t_L g124 ( .A(n_6), .B(n_30), .Y(n_124) );
BUFx2_ASAP7_75t_L g877 ( .A(n_6), .Y(n_877) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_7), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_8), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_11), .B(n_195), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g865 ( .A(n_12), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_13), .A2(n_101), .B1(n_192), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_14), .A2(n_31), .B1(n_572), .B2(n_573), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_15), .B(n_195), .Y(n_614) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_16), .A2(n_45), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_17), .B(n_284), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g554 ( .A(n_18), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g859 ( .A1(n_19), .A2(n_94), .B1(n_860), .B2(n_861), .Y(n_859) );
INVx1_ASAP7_75t_L g861 ( .A(n_19), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_20), .A2(n_38), .B1(n_182), .B2(n_200), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g176 ( .A(n_21), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_22), .A2(n_43), .B1(n_182), .B2(n_549), .Y(n_584) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_23), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_24), .B(n_572), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_25), .B(n_147), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_26), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_27), .B(n_205), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_28), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g113 ( .A1(n_29), .A2(n_82), .B1(n_114), .B2(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
HB1xp67_ASAP7_75t_L g879 ( .A(n_30), .Y(n_879) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_32), .A2(n_85), .B1(n_144), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_33), .A2(n_37), .B1(n_144), .B2(n_562), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_35), .A2(n_48), .B1(n_549), .B2(n_551), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_36), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_39), .B(n_195), .Y(n_245) );
INVx2_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_41), .B(n_196), .Y(n_279) );
INVx1_ASAP7_75t_L g122 ( .A(n_42), .Y(n_122) );
BUFx3_ASAP7_75t_L g524 ( .A(n_42), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_44), .B(n_164), .Y(n_286) );
AND2x2_ASAP7_75t_L g184 ( .A(n_46), .B(n_164), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_47), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_49), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_50), .B(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_51), .A2(n_78), .B1(n_508), .B2(n_509), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_51), .Y(n_508) );
XNOR2x1_ASAP7_75t_L g531 ( .A(n_51), .B(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_52), .A2(n_68), .B1(n_200), .B2(n_551), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_53), .A2(n_72), .B1(n_144), .B2(n_562), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_54), .B(n_155), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_55), .A2(n_149), .B(n_174), .C(n_175), .Y(n_173) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_56), .A2(n_98), .B1(n_549), .B2(n_560), .Y(n_623) );
INVx1_ASAP7_75t_L g140 ( .A(n_57), .Y(n_140) );
AND2x4_ASAP7_75t_L g161 ( .A(n_58), .B(n_162), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_59), .A2(n_60), .B1(n_182), .B2(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_61), .B(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_62), .B(n_164), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_63), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_64), .B(n_182), .Y(n_248) );
INVx1_ASAP7_75t_L g162 ( .A(n_65), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_66), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_67), .B(n_205), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_69), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_70), .B(n_144), .Y(n_143) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_71), .B(n_156), .C(n_196), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_73), .A2(n_105), .B1(n_872), .B2(n_886), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_74), .B(n_144), .Y(n_226) );
INVx2_ASAP7_75t_L g151 ( .A(n_75), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_76), .B(n_195), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_77), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g509 ( .A(n_78), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_79), .B(n_202), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_80), .A2(n_97), .B1(n_174), .B2(n_182), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_81), .Y(n_588) );
INVx1_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g856 ( .A1(n_83), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
CKINVDCx5p33_ASAP7_75t_R g857 ( .A(n_83), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_84), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_86), .A2(n_91), .B1(n_147), .B2(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_87), .B(n_195), .Y(n_194) );
NAND2xp33_ASAP7_75t_SL g218 ( .A(n_88), .B(n_201), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_89), .B(n_193), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_90), .B(n_205), .Y(n_619) );
CKINVDCx5p33_ASAP7_75t_R g566 ( .A(n_92), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_93), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g530 ( .A(n_93), .Y(n_530) );
INVx1_ASAP7_75t_L g860 ( .A(n_94), .Y(n_860) );
NAND2xp33_ASAP7_75t_L g617 ( .A(n_95), .B(n_195), .Y(n_617) );
NAND2xp33_ASAP7_75t_L g227 ( .A(n_96), .B(n_201), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_99), .B(n_164), .Y(n_163) );
NAND3xp33_ASAP7_75t_L g214 ( .A(n_100), .B(n_201), .C(n_213), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_102), .B(n_144), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_103), .B(n_147), .Y(n_153) );
AO221x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B1(n_519), .B2(n_525), .C(n_864), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x6_ASAP7_75t_SL g521 ( .A(n_108), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_109), .B(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_516), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_125), .B(n_510), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .Y(n_112) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_113), .B(n_517), .C(n_518), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_116), .Y(n_518) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx12f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
CKINVDCx8_ASAP7_75t_R g515 ( .A(n_119), .Y(n_515) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_122), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_123), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR2x1_ASAP7_75t_L g871 ( .A(n_124), .B(n_524), .Y(n_871) );
XOR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_507), .Y(n_125) );
XNOR2x1_ASAP7_75t_L g517 ( .A(n_126), .B(n_507), .Y(n_517) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g532 ( .A(n_127), .Y(n_532) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_402), .Y(n_127) );
NOR2x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_337), .Y(n_128) );
NAND3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_260), .C(n_310), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_185), .B(n_220), .C(n_237), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OR2x2_ASAP7_75t_L g476 ( .A(n_132), .B(n_395), .Y(n_476) );
OR2x2_ASAP7_75t_L g487 ( .A(n_132), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_133), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g378 ( .A(n_133), .B(n_267), .Y(n_378) );
AND2x2_ASAP7_75t_L g499 ( .A(n_133), .B(n_309), .Y(n_499) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_165), .Y(n_133) );
INVx2_ASAP7_75t_L g329 ( .A(n_134), .Y(n_329) );
AND2x2_ASAP7_75t_L g344 ( .A(n_134), .B(n_296), .Y(n_344) );
AND2x2_ASAP7_75t_L g353 ( .A(n_134), .B(n_222), .Y(n_353) );
AND2x2_ASAP7_75t_L g422 ( .A(n_134), .B(n_308), .Y(n_422) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g235 ( .A(n_135), .Y(n_235) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_141), .B(n_163), .Y(n_135) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_136), .A2(n_189), .B(n_204), .Y(n_188) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_136), .A2(n_189), .B(n_204), .Y(n_303) );
OAI21xp33_ASAP7_75t_SL g394 ( .A1(n_136), .A2(n_141), .B(n_163), .Y(n_394) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_137), .B(n_554), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_137), .B(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g169 ( .A(n_138), .Y(n_169) );
INVx2_ASAP7_75t_L g259 ( .A(n_138), .Y(n_259) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_139), .Y(n_206) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_152), .B(n_160), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_149), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_144), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_180) );
INVx1_ASAP7_75t_L g551 ( .A(n_144), .Y(n_551) );
INVx1_ASAP7_75t_L g560 ( .A(n_144), .Y(n_560) );
INVx4_ASAP7_75t_L g562 ( .A(n_144), .Y(n_562) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx1_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
INVx2_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
INVx1_ASAP7_75t_L g193 ( .A(n_145), .Y(n_193) );
BUFx6f_ASAP7_75t_L g195 ( .A(n_145), .Y(n_195) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_145), .Y(n_201) );
INVx1_ASAP7_75t_L g217 ( .A(n_145), .Y(n_217) );
INVx1_ASAP7_75t_L g256 ( .A(n_145), .Y(n_256) );
INVx1_ASAP7_75t_L g559 ( .A(n_147), .Y(n_559) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_149), .A2(n_216), .B(n_218), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_149), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_149), .A2(n_244), .B(n_245), .Y(n_243) );
BUFx4f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g159 ( .A(n_151), .Y(n_159) );
BUFx8_ASAP7_75t_L g196 ( .A(n_151), .Y(n_196) );
INVx1_ASAP7_75t_L g213 ( .A(n_151), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_157), .Y(n_152) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_160), .A2(n_190), .B(n_197), .Y(n_189) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_211), .B(n_215), .Y(n_210) );
AND2x4_ASAP7_75t_SL g232 ( .A(n_160), .B(n_206), .Y(n_232) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_160), .A2(n_243), .B(n_246), .Y(n_242) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_160), .A2(n_278), .B(n_281), .Y(n_277) );
BUFx10_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx10_ASAP7_75t_L g171 ( .A(n_161), .Y(n_171) );
INVx1_ASAP7_75t_L g586 ( .A(n_161), .Y(n_586) );
AND2x2_ASAP7_75t_L g393 ( .A(n_165), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g236 ( .A(n_166), .B(n_208), .Y(n_236) );
INVx2_ASAP7_75t_L g265 ( .A(n_166), .Y(n_265) );
AOI21x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_172), .B(n_184), .Y(n_166) );
NOR2xp67_ASAP7_75t_SL g167 ( .A(n_168), .B(n_170), .Y(n_167) );
INVx2_ASAP7_75t_L g552 ( .A(n_168), .Y(n_552) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO31x2_ASAP7_75t_L g250 ( .A1(n_169), .A2(n_171), .A3(n_251), .B(n_257), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g565 ( .A(n_169), .B(n_566), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_169), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g546 ( .A(n_170), .Y(n_546) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO31x2_ASAP7_75t_L g556 ( .A1(n_171), .A2(n_557), .A3(n_564), .B(n_565), .Y(n_556) );
AO31x2_ASAP7_75t_L g569 ( .A1(n_171), .A2(n_570), .A3(n_576), .B(n_577), .Y(n_569) );
AO31x2_ASAP7_75t_L g632 ( .A1(n_171), .A2(n_633), .A3(n_636), .B(n_637), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_178), .Y(n_172) );
INVx1_ASAP7_75t_L g230 ( .A(n_174), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
INVx2_ASAP7_75t_SL g602 ( .A(n_177), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_179), .A2(n_252), .B1(n_254), .B2(n_255), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_179), .A2(n_254), .B1(n_548), .B2(n_550), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g570 ( .A1(n_179), .A2(n_254), .B1(n_571), .B2(n_574), .Y(n_570) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_179), .A2(n_254), .B1(n_583), .B2(n_584), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_179), .A2(n_254), .B1(n_634), .B2(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g253 ( .A(n_182), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g278 ( .A1(n_182), .A2(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g430 ( .A(n_185), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_207), .Y(n_186) );
INVx1_ASAP7_75t_L g450 ( .A(n_187), .Y(n_450) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g288 ( .A(n_188), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g371 ( .A(n_188), .B(n_276), .Y(n_371) );
O2A1O1Ixp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_194), .C(n_196), .Y(n_190) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_195), .A2(n_212), .B(n_214), .Y(n_211) );
INVx1_ASAP7_75t_L g284 ( .A(n_195), .Y(n_284) );
INVx3_ASAP7_75t_L g549 ( .A(n_195), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_196), .A2(n_247), .B(n_248), .Y(n_246) );
INVx6_ASAP7_75t_L g254 ( .A(n_196), .Y(n_254) );
O2A1O1Ixp5_ASAP7_75t_L g612 ( .A1(n_196), .A2(n_562), .B(n_613), .C(n_614), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_202), .Y(n_197) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g572 ( .A(n_201), .Y(n_572) );
INVx2_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_203), .A2(n_229), .B1(n_230), .B2(n_231), .Y(n_228) );
INVx2_ASAP7_75t_L g636 ( .A(n_205), .Y(n_636) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_SL g209 ( .A(n_206), .Y(n_209) );
INVx2_ASAP7_75t_L g241 ( .A(n_206), .Y(n_241) );
BUFx3_ASAP7_75t_L g576 ( .A(n_206), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_206), .B(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g610 ( .A(n_206), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_206), .B(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_206), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g297 ( .A(n_207), .B(n_235), .Y(n_297) );
INVxp67_ASAP7_75t_L g446 ( .A(n_207), .Y(n_446) );
OR2x2_ASAP7_75t_L g488 ( .A(n_207), .B(n_222), .Y(n_488) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_219), .Y(n_208) );
INVx1_ASAP7_75t_L g285 ( .A(n_213), .Y(n_285) );
INVx1_ASAP7_75t_SL g563 ( .A(n_213), .Y(n_563) );
INVx1_ASAP7_75t_L g604 ( .A(n_213), .Y(n_604) );
INVx1_ASAP7_75t_L g573 ( .A(n_217), .Y(n_573) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_233), .Y(n_220) );
INVx1_ASAP7_75t_L g343 ( .A(n_221), .Y(n_343) );
AND2x2_ASAP7_75t_L g497 ( .A(n_221), .B(n_393), .Y(n_497) );
BUFx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g268 ( .A(n_222), .Y(n_268) );
INVx4_ASAP7_75t_L g308 ( .A(n_222), .Y(n_308) );
AND2x4_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
OAI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_228), .B(n_232), .Y(n_224) );
AND2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g324 ( .A(n_234), .B(n_307), .Y(n_324) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g361 ( .A(n_235), .B(n_309), .Y(n_361) );
INVx2_ASAP7_75t_L g327 ( .A(n_236), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_236), .B(n_332), .Y(n_495) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_239), .B(n_408), .Y(n_407) );
BUFx2_ASAP7_75t_L g480 ( .A(n_239), .Y(n_480) );
AND2x2_ASAP7_75t_L g494 ( .A(n_239), .B(n_316), .Y(n_494) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_250), .Y(n_239) );
INVx1_ASAP7_75t_L g274 ( .A(n_240), .Y(n_274) );
AND2x2_ASAP7_75t_L g429 ( .A(n_240), .B(n_336), .Y(n_429) );
OR2x2_ASAP7_75t_L g466 ( .A(n_240), .B(n_250), .Y(n_466) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_249), .Y(n_240) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_241), .A2(n_277), .B(n_286), .Y(n_276) );
OA21x2_ASAP7_75t_L g289 ( .A1(n_241), .A2(n_277), .B(n_286), .Y(n_289) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_241), .A2(n_242), .B(n_249), .Y(n_292) );
AND2x2_ASAP7_75t_L g275 ( .A(n_250), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g290 ( .A(n_250), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g336 ( .A(n_250), .Y(n_336) );
OR2x2_ASAP7_75t_L g349 ( .A(n_250), .B(n_289), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_250), .B(n_289), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_254), .A2(n_558), .B1(n_561), .B2(n_563), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_254), .A2(n_601), .B1(n_603), .B2(n_604), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_254), .A2(n_616), .B(n_617), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_254), .A2(n_563), .B1(n_623), .B2(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g575 ( .A(n_256), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
BUFx2_ASAP7_75t_L g564 ( .A(n_259), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_270), .B(n_293), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AOI31xp33_ASAP7_75t_L g339 ( .A1(n_262), .A2(n_340), .A3(n_342), .B(n_345), .Y(n_339) );
OR2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
AND2x2_ASAP7_75t_L g352 ( .A(n_263), .B(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g362 ( .A(n_264), .Y(n_362) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_264), .Y(n_368) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g296 ( .A(n_265), .Y(n_296) );
AND2x2_ASAP7_75t_L g325 ( .A(n_265), .B(n_309), .Y(n_325) );
INVx2_ASAP7_75t_L g375 ( .A(n_265), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_266), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g400 ( .A(n_267), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g449 ( .A(n_267), .B(n_450), .Y(n_449) );
AOI33xp33_ASAP7_75t_L g504 ( .A1(n_267), .A2(n_334), .A3(n_344), .B1(n_371), .B2(n_480), .B3(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx2_ASAP7_75t_L g309 ( .A(n_269), .Y(n_309) );
INVx1_ASAP7_75t_L g396 ( .A(n_269), .Y(n_396) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_272), .B(n_287), .Y(n_271) );
INVx2_ASAP7_75t_L g304 ( .A(n_272), .Y(n_304) );
AND2x2_ASAP7_75t_L g385 ( .A(n_272), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
INVx1_ASAP7_75t_L g347 ( .A(n_273), .Y(n_347) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g415 ( .A(n_274), .B(n_302), .Y(n_415) );
AND2x2_ASAP7_75t_L g365 ( .A(n_275), .B(n_359), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_275), .B(n_383), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_275), .B(n_415), .Y(n_464) );
AND2x2_ASAP7_75t_L g301 ( .A(n_276), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g320 ( .A(n_276), .B(n_315), .Y(n_320) );
INVx1_ASAP7_75t_L g335 ( .A(n_276), .Y(n_335) );
AOI21x1_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_285), .Y(n_281) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
INVx1_ASAP7_75t_L g390 ( .A(n_288), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_288), .B(n_483), .Y(n_485) );
AND2x2_ASAP7_75t_L g498 ( .A(n_288), .B(n_314), .Y(n_498) );
AND2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_302), .Y(n_316) );
INVx2_ASAP7_75t_L g298 ( .A(n_290), .Y(n_298) );
AND2x2_ASAP7_75t_L g412 ( .A(n_290), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g471 ( .A(n_290), .B(n_383), .Y(n_471) );
BUFx2_ASAP7_75t_L g453 ( .A(n_291), .Y(n_453) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx3_ASAP7_75t_L g315 ( .A(n_292), .Y(n_315) );
OAI32xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_298), .A3(n_299), .B1(n_304), .B2(n_305), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g401 ( .A(n_296), .Y(n_401) );
AND2x2_ASAP7_75t_L g431 ( .A(n_296), .B(n_353), .Y(n_431) );
AND2x2_ASAP7_75t_L g373 ( .A(n_297), .B(n_374), .Y(n_373) );
AND3x2_ASAP7_75t_L g380 ( .A(n_297), .B(n_307), .C(n_375), .Y(n_380) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_300), .A2(n_322), .B1(n_331), .B2(n_333), .Y(n_330) );
OAI322xp33_ASAP7_75t_L g478 ( .A1(n_300), .A2(n_399), .A3(n_479), .B1(n_480), .B2(n_481), .C1(n_482), .C2(n_485), .Y(n_478) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g500 ( .A(n_301), .B(n_483), .Y(n_500) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_302), .Y(n_319) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_302), .Y(n_359) );
BUFx3_ASAP7_75t_L g383 ( .A(n_302), .Y(n_383) );
INVx1_ASAP7_75t_L g409 ( .A(n_302), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_302), .Y(n_413) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g367 ( .A(n_306), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g418 ( .A(n_307), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_307), .B(n_375), .Y(n_469) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2x1_ASAP7_75t_L g328 ( .A(n_308), .B(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
AND2x2_ASAP7_75t_L g374 ( .A(n_308), .B(n_375), .Y(n_374) );
OR2x2_ASAP7_75t_L g395 ( .A(n_308), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_309), .B(n_422), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_317), .B(n_321), .C(n_330), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AOI31xp33_ASAP7_75t_L g472 ( .A1(n_312), .A2(n_473), .A3(n_475), .B(n_476), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_316), .Y(n_312) );
AND2x4_ASAP7_75t_L g425 ( .A(n_313), .B(n_334), .Y(n_425) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g441 ( .A(n_315), .B(n_335), .Y(n_441) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
NAND2x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_326), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g481 ( .A(n_324), .Y(n_481) );
AND2x2_ASAP7_75t_L g341 ( .A(n_325), .B(n_332), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_326), .A2(n_411), .B1(n_414), .B2(n_416), .Y(n_410) );
OR2x6_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_SL g468 ( .A(n_329), .Y(n_468) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g438 ( .A(n_334), .B(n_383), .Y(n_438) );
INVx2_ASAP7_75t_L g484 ( .A(n_334), .Y(n_484) );
AND2x4_ASAP7_75t_L g492 ( .A(n_334), .B(n_413), .Y(n_492) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND3xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_354), .C(n_384), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_350), .Y(n_338) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_341), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
AND2x4_ASAP7_75t_L g405 ( .A(n_343), .B(n_360), .Y(n_405) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_346), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g436 ( .A(n_348), .B(n_415), .Y(n_436) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_349), .Y(n_356) );
INVx1_ASAP7_75t_L g474 ( .A(n_349), .Y(n_474) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g503 ( .A(n_352), .Y(n_503) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_360), .B(n_363), .C(n_376), .Y(n_354) );
NOR3x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .C(n_358), .Y(n_355) );
NAND2x1_ASAP7_75t_L g424 ( .A(n_358), .B(n_425), .Y(n_424) );
BUFx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2x1p5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_362), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_366), .B1(n_369), .B2(n_372), .Y(n_363) );
INVxp67_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g457 ( .A(n_368), .Y(n_457) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g452 ( .A(n_371), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g506 ( .A(n_374), .Y(n_506) );
AOI21xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g460 ( .A(n_381), .Y(n_460) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx2_ASAP7_75t_L g387 ( .A(n_383), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_383), .B(n_441), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B(n_389), .Y(n_384) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_387), .B(n_474), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B1(n_397), .B2(n_399), .Y(n_389) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g442 ( .A(n_392), .Y(n_442) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g417 ( .A(n_393), .B(n_418), .Y(n_417) );
BUFx2_ASAP7_75t_L g434 ( .A(n_394), .Y(n_434) );
INVx1_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_458), .Y(n_402) );
NAND3xp33_ASAP7_75t_SL g403 ( .A(n_404), .B(n_419), .C(n_432), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g465 ( .A(n_408), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2x1p5_ASAP7_75t_L g462 ( .A(n_417), .B(n_445), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B1(n_426), .B2(n_430), .Y(n_419) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g475 ( .A(n_425), .Y(n_475) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g447 ( .A1(n_427), .A2(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_443), .B1(n_447), .B2(n_455), .Y(n_432) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_437), .Y(n_433) );
INVxp67_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_442), .Y(n_437) );
INVx1_ASAP7_75t_L g502 ( .A(n_438), .Y(n_502) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
INVx2_ASAP7_75t_L g483 ( .A(n_453), .Y(n_483) );
INVxp67_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_459), .B(n_477), .Y(n_458) );
AOI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_463), .C(n_472), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B(n_467), .C(n_470), .Y(n_463) );
OR2x2_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .C(n_501), .Y(n_477) );
OR2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_484), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_489), .B1(n_493), .B2(n_495), .C(n_496), .Y(n_486) );
NOR2xp67_ASAP7_75t_L g489 ( .A(n_490), .B(n_492), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
OAI21xp33_ASAP7_75t_SL g501 ( .A1(n_502), .A2(n_503), .B(n_504), .Y(n_501) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g864 ( .A1(n_511), .A2(n_865), .B(n_866), .Y(n_864) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx4_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
OAI22x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_855), .B1(n_856), .B2(n_862), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_531), .B(n_533), .Y(n_526) );
AOI21x1_ASAP7_75t_L g863 ( .A1(n_527), .A2(n_531), .B(n_533), .Y(n_863) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx8_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g870 ( .A(n_529), .B(n_871), .Y(n_870) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g537 ( .A(n_530), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g881 ( .A(n_537), .B(n_882), .C(n_885), .Y(n_881) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_764), .Y(n_538) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_703), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_541), .B(n_654), .C(n_673), .D(n_684), .Y(n_540) );
O2A1O1Ixp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_589), .B(n_596), .C(n_627), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_567), .Y(n_542) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_543), .B(n_719), .C(n_720), .Y(n_718) );
AND2x2_ASAP7_75t_L g800 ( .A(n_543), .B(n_682), .Y(n_800) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
AND2x2_ASAP7_75t_L g644 ( .A(n_544), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g662 ( .A(n_544), .B(n_663), .Y(n_662) );
INVx3_ASAP7_75t_L g679 ( .A(n_544), .Y(n_679) );
AND2x2_ASAP7_75t_L g724 ( .A(n_544), .B(n_569), .Y(n_724) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g593 ( .A(n_545), .Y(n_593) );
AND2x4_ASAP7_75t_L g672 ( .A(n_545), .B(n_663), .Y(n_672) );
AO31x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .A3(n_552), .B(n_553), .Y(n_545) );
AO31x2_ASAP7_75t_L g621 ( .A1(n_546), .A2(n_564), .A3(n_622), .B(n_625), .Y(n_621) );
AO31x2_ASAP7_75t_L g581 ( .A1(n_552), .A2(n_582), .A3(n_585), .B(n_587), .Y(n_581) );
AND2x2_ASAP7_75t_L g594 ( .A(n_555), .B(n_595), .Y(n_594) );
AND2x4_ASAP7_75t_L g647 ( .A(n_555), .B(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_555), .Y(n_670) );
INVx1_ASAP7_75t_L g681 ( .A(n_555), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_555), .B(n_579), .Y(n_690) );
INVx2_ASAP7_75t_L g697 ( .A(n_555), .Y(n_697) );
INVx4_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g642 ( .A(n_556), .B(n_569), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_556), .B(n_649), .Y(n_715) );
AND2x2_ASAP7_75t_L g723 ( .A(n_556), .B(n_581), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_556), .B(n_770), .Y(n_769) );
BUFx2_ASAP7_75t_L g776 ( .A(n_556), .Y(n_776) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g792 ( .A(n_568), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_579), .Y(n_568) );
INVx1_ASAP7_75t_L g595 ( .A(n_569), .Y(n_595) );
INVx1_ASAP7_75t_L g649 ( .A(n_569), .Y(n_649) );
INVx2_ASAP7_75t_L g683 ( .A(n_569), .Y(n_683) );
OR2x2_ASAP7_75t_L g687 ( .A(n_569), .B(n_581), .Y(n_687) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_569), .Y(n_736) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_576), .A2(n_585), .A3(n_600), .B(n_605), .Y(n_599) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g709 ( .A(n_580), .B(n_593), .Y(n_709) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_581), .Y(n_645) );
INVx2_ASAP7_75t_L g663 ( .A(n_581), .Y(n_663) );
AND2x4_ASAP7_75t_L g682 ( .A(n_581), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g770 ( .A(n_581), .Y(n_770) );
INVx2_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx2_ASAP7_75t_SL g618 ( .A(n_586), .Y(n_618) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_594), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g688 ( .A(n_592), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_592), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g751 ( .A(n_593), .Y(n_751) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_607), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_598), .B(n_608), .Y(n_701) );
INVx1_ASAP7_75t_L g799 ( .A(n_598), .Y(n_799) );
BUFx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g639 ( .A(n_599), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g653 ( .A(n_599), .B(n_632), .Y(n_653) );
AND2x4_ASAP7_75t_L g676 ( .A(n_599), .B(n_620), .Y(n_676) );
INVx2_ASAP7_75t_L g693 ( .A(n_599), .Y(n_693) );
AND2x2_ASAP7_75t_L g719 ( .A(n_599), .B(n_621), .Y(n_719) );
INVx1_ASAP7_75t_L g784 ( .A(n_599), .Y(n_784) );
AND2x2_ASAP7_75t_L g744 ( .A(n_607), .B(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_620), .Y(n_607) );
AND2x2_ASAP7_75t_L g710 ( .A(n_608), .B(n_667), .Y(n_710) );
AND2x4_ASAP7_75t_L g726 ( .A(n_608), .B(n_693), .Y(n_726) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
BUFx2_ASAP7_75t_L g720 ( .A(n_609), .Y(n_720) );
OAI21x1_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_619), .Y(n_609) );
OAI21x1_ASAP7_75t_L g641 ( .A1(n_610), .A2(n_611), .B(n_619), .Y(n_641) );
OAI21x1_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B(n_618), .Y(n_611) );
INVx2_ASAP7_75t_L g652 ( .A(n_620), .Y(n_652) );
INVx3_ASAP7_75t_L g658 ( .A(n_620), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_620), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_620), .B(n_787), .Y(n_786) );
INVx3_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g692 ( .A(n_621), .B(n_693), .Y(n_692) );
BUFx2_ASAP7_75t_L g816 ( .A(n_621), .Y(n_816) );
OAI33xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_642), .A3(n_643), .B1(n_644), .B2(n_646), .B3(n_650), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_639), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g750 ( .A(n_631), .B(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g659 ( .A(n_632), .B(n_641), .Y(n_659) );
INVx2_ASAP7_75t_L g667 ( .A(n_632), .Y(n_667) );
INVx1_ASAP7_75t_L g675 ( .A(n_632), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_639), .A2(n_695), .B1(n_698), .B2(n_702), .Y(n_694) );
OR2x2_ASAP7_75t_L g834 ( .A(n_639), .B(n_652), .Y(n_834) );
AND2x4_ASAP7_75t_L g738 ( .A(n_640), .B(n_700), .Y(n_738) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_641), .B(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_642), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g702 ( .A(n_642), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_642), .B(n_678), .Y(n_780) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g753 ( .A(n_644), .Y(n_753) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g811 ( .A(n_647), .B(n_679), .Y(n_811) );
NAND2x1_ASAP7_75t_L g829 ( .A(n_647), .B(n_678), .Y(n_829) );
AND2x2_ASAP7_75t_L g853 ( .A(n_647), .B(n_672), .Y(n_853) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g843 ( .A(n_651), .B(n_720), .Y(n_843) );
NOR2x1p5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
AND2x2_ASAP7_75t_L g777 ( .A(n_652), .B(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g745 ( .A(n_653), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_660), .B1(n_664), .B2(n_668), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
AND2x2_ASAP7_75t_L g752 ( .A(n_657), .B(n_720), .Y(n_752) );
AND2x2_ASAP7_75t_L g789 ( .A(n_657), .B(n_738), .Y(n_789) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x4_ASAP7_75t_L g664 ( .A(n_658), .B(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_658), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g830 ( .A(n_658), .B(n_659), .Y(n_830) );
AND2x2_ASAP7_75t_L g691 ( .A(n_659), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g810 ( .A(n_659), .B(n_676), .Y(n_810) );
AND2x2_ASAP7_75t_L g854 ( .A(n_659), .B(n_719), .Y(n_854) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI222xp33_ASAP7_75t_L g788 ( .A1(n_664), .A2(n_789), .B1(n_790), .B2(n_793), .C1(n_795), .C2(n_796), .Y(n_788) );
AND2x2_ASAP7_75t_L g711 ( .A(n_665), .B(n_679), .Y(n_711) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g742 ( .A(n_666), .Y(n_742) );
INVxp67_ASAP7_75t_SL g787 ( .A(n_666), .Y(n_787) );
INVx2_ASAP7_75t_L g700 ( .A(n_667), .Y(n_700) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g757 ( .A(n_670), .Y(n_757) );
INVx2_ASAP7_75t_L g763 ( .A(n_671), .Y(n_763) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x4_ASAP7_75t_L g747 ( .A(n_672), .B(n_736), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
AND2x4_ASAP7_75t_L g778 ( .A(n_675), .B(n_726), .Y(n_778) );
INVx2_ASAP7_75t_L g825 ( .A(n_675), .Y(n_825) );
AND2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
INVx4_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OR2x2_ASAP7_75t_L g768 ( .A(n_679), .B(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g802 ( .A(n_679), .B(n_687), .Y(n_802) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
INVx1_ASAP7_75t_L g707 ( .A(n_681), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_682), .B(n_772), .Y(n_771) );
AND2x4_ASAP7_75t_L g814 ( .A(n_682), .B(n_730), .Y(n_814) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_689), .B(n_691), .C(n_694), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
OR2x2_ASAP7_75t_L g695 ( .A(n_687), .B(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g731 ( .A(n_687), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_688), .B(n_723), .Y(n_827) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g803 ( .A(n_690), .B(n_772), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_692), .B(n_742), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_692), .A2(n_708), .B1(n_750), .B2(n_752), .Y(n_749) );
AND2x2_ASAP7_75t_L g755 ( .A(n_692), .B(n_720), .Y(n_755) );
AND2x2_ASAP7_75t_L g824 ( .A(n_692), .B(n_825), .Y(n_824) );
O2A1O1Ixp33_ASAP7_75t_L g817 ( .A1(n_695), .A2(n_797), .B(n_818), .C(n_821), .Y(n_817) );
INVx2_ASAP7_75t_L g730 ( .A(n_697), .Y(n_730) );
OR2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVx1_ASAP7_75t_L g808 ( .A(n_700), .Y(n_808) );
INVx1_ASAP7_75t_L g733 ( .A(n_701), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_702), .A2(n_749), .B1(n_753), .B2(n_754), .Y(n_748) );
NAND3xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_716), .C(n_739), .Y(n_703) );
AO22x1_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B1(n_711), .B2(n_712), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_709), .Y(n_842) );
OR2x2_ASAP7_75t_L g849 ( .A(n_709), .B(n_730), .Y(n_849) );
AND2x2_ASAP7_75t_L g761 ( .A(n_710), .B(n_719), .Y(n_761) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g837 ( .A(n_715), .Y(n_837) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_721), .C(n_727), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g759 ( .A(n_719), .Y(n_759) );
AND2x4_ASAP7_75t_SL g795 ( .A(n_719), .B(n_738), .Y(n_795) );
INVx1_ASAP7_75t_SL g806 ( .A(n_719), .Y(n_806) );
OR2x2_ASAP7_75t_L g758 ( .A(n_720), .B(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
AND2x4_ASAP7_75t_L g735 ( .A(n_723), .B(n_736), .Y(n_735) );
AND2x2_ASAP7_75t_L g793 ( .A(n_724), .B(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g815 ( .A(n_726), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g840 ( .A(n_726), .B(n_820), .Y(n_840) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_732), .B1(n_734), .B2(n_737), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
AND2x4_ASAP7_75t_L g775 ( .A(n_731), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g797 ( .A(n_731), .Y(n_797) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g852 ( .A(n_735), .B(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_748), .C(n_756), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_743), .B(n_746), .Y(n_740) );
INVx1_ASAP7_75t_L g821 ( .A(n_742), .Y(n_821) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AOI222xp33_ASAP7_75t_L g844 ( .A1(n_747), .A2(n_845), .B1(n_848), .B2(n_850), .C1(n_852), .C2(n_854), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_750), .B(n_840), .Y(n_839) );
INVx3_ASAP7_75t_L g773 ( .A(n_751), .Y(n_773) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_758), .B(n_760), .C(n_762), .Y(n_756) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_822), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_766), .B(n_788), .C(n_798), .D(n_809), .Y(n_765) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_777), .B1(n_779), .B2(n_781), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .C(n_774), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_768), .B(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g794 ( .A(n_770), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_772), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AND2x4_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
AND2x2_ASAP7_75t_L g819 ( .A(n_784), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g833 ( .A(n_785), .Y(n_833) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_786), .Y(n_851) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx3_ASAP7_75t_L g846 ( .A(n_795), .Y(n_846) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_800), .B(n_801), .C(n_807), .Y(n_798) );
AOI21xp33_ASAP7_75t_SL g801 ( .A1(n_802), .A2(n_803), .B(n_804), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_802), .B(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_811), .B1(n_812), .B2(n_815), .C(n_817), .Y(n_809) );
INVx1_ASAP7_75t_L g847 ( .A(n_810), .Y(n_847) );
AOI31xp33_ASAP7_75t_L g831 ( .A1(n_813), .A2(n_832), .A3(n_833), .B(n_834), .Y(n_831) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g820 ( .A(n_816), .Y(n_820) );
INVxp67_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND3xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_835), .C(n_844), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_826), .B1(n_828), .B2(n_830), .C(n_831), .Y(n_823) );
INVx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_SL g832 ( .A(n_830), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_836), .A2(n_838), .B1(n_841), .B2(n_843), .Y(n_835) );
HB1xp67_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
BUFx10_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
BUFx6f_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_873), .Y(n_887) );
INVx8_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OR2x6_ASAP7_75t_L g874 ( .A(n_875), .B(n_880), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NOR2xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
INVxp33_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
INVx2_ASAP7_75t_SL g882 ( .A(n_883), .Y(n_882) );
INVx4_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
endmodule