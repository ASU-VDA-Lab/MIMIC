module fake_aes_339_n_1174 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_1174);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_1174;
wire n_1173;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1124;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_1158;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_252;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_1122;
wire n_528;
wire n_383;
wire n_288;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_1128;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_1118;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_1161;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_1163;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_1121;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_769;
wire n_927;
wire n_596;
wire n_286;
wire n_246;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_1097;
wire n_572;
wire n_1017;
wire n_324;
wire n_1078;
wire n_773;
wire n_1094;
wire n_1125;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_847;
wire n_1169;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_1042;
wire n_975;
wire n_1060;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_955;
wire n_479;
wire n_623;
wire n_593;
wire n_945;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_529;
wire n_312;
wire n_1132;
wire n_1011;
wire n_1025;
wire n_880;
wire n_1101;
wire n_1155;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_844;
wire n_818;
wire n_1160;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1063;
wire n_767;
wire n_828;
wire n_1138;
wire n_293;
wire n_1014;
wire n_506;
wire n_533;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_1171;
wire n_665;
wire n_571;
wire n_1154;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_950;
wire n_935;
wire n_460;
wire n_1046;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_1076;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_1145;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_1167;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_1140;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_1147;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_1130;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_1129;
wire n_450;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_446;
wire n_420;
wire n_621;
wire n_423;
wire n_342;
wire n_666;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_1157;
wire n_974;
wire n_1153;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_956;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_1135;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_1144;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_1152;
wire n_681;
wire n_1139;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_1149;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_1170;
wire n_419;
wire n_851;
wire n_1119;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_908;
wire n_1133;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_1159;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1131;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1069;
wire n_1021;
wire n_811;
wire n_1123;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_1156;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_1043;
wire n_1141;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_1172;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_1136;
wire n_397;
wire n_1142;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_1027;
wire n_1007;
wire n_859;
wire n_1117;
wire n_1040;
wire n_1165;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_1143;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_1168;
wire n_377;
wire n_510;
wire n_343;
wire n_1112;
wire n_1075;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1164;
wire n_1038;
wire n_341;
wire n_1162;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_1073;
wire n_323;
wire n_868;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_266;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_1150;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_1104;
wire n_742;
wire n_1120;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_1134;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_1146;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_1137;
wire n_781;
wire n_916;
wire n_421;
wire n_1148;
wire n_709;
wire n_739;
wire n_1166;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_257;
wire n_992;
wire n_1127;
wire n_269;
BUFx3_ASAP7_75t_L g242 ( .A(n_103), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_2), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_193), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_223), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_128), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_74), .Y(n_247) );
NOR2xp67_ASAP7_75t_L g248 ( .A(n_8), .B(n_122), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_82), .Y(n_249) );
NOR2xp67_ASAP7_75t_L g250 ( .A(n_145), .B(n_123), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
INVxp67_ASAP7_75t_SL g252 ( .A(n_141), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_70), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_62), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g255 ( .A(n_0), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_56), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_96), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_232), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_136), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_194), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_8), .Y(n_261) );
INVx1_ASAP7_75t_SL g262 ( .A(n_80), .Y(n_262) );
CKINVDCx20_ASAP7_75t_R g263 ( .A(n_87), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_44), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_28), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_85), .Y(n_266) );
CKINVDCx6p67_ASAP7_75t_R g267 ( .A(n_94), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_212), .Y(n_268) );
INVxp33_ASAP7_75t_SL g269 ( .A(n_135), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_234), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_191), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_2), .B(n_28), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_14), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_20), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_138), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_63), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_42), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_7), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_18), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_156), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_107), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_166), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_101), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_97), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_236), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_77), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_59), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_216), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_150), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_21), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_181), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_153), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_131), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_209), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_25), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_182), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_51), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_109), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_14), .B(n_5), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_39), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_47), .Y(n_301) );
CKINVDCx16_ASAP7_75t_R g302 ( .A(n_224), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_124), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_227), .Y(n_304) );
INVxp33_ASAP7_75t_L g305 ( .A(n_214), .Y(n_305) );
OR2x2_ASAP7_75t_L g306 ( .A(n_52), .B(n_155), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_238), .Y(n_307) );
BUFx5_ASAP7_75t_L g308 ( .A(n_118), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_104), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_208), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_89), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_116), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_59), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_29), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_110), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_159), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_207), .Y(n_317) );
INVxp67_ASAP7_75t_L g318 ( .A(n_37), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_167), .Y(n_319) );
CKINVDCx14_ASAP7_75t_R g320 ( .A(n_42), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_149), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_5), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_1), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_140), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_29), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_38), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_168), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_171), .Y(n_328) );
CKINVDCx20_ASAP7_75t_R g329 ( .A(n_139), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_72), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_213), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_130), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_47), .Y(n_333) );
INVxp67_ASAP7_75t_L g334 ( .A(n_184), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_137), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_95), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_205), .Y(n_337) );
INVxp33_ASAP7_75t_SL g338 ( .A(n_225), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_36), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_0), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_226), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_230), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_148), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_1), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_211), .Y(n_345) );
INVx2_ASAP7_75t_SL g346 ( .A(n_83), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_13), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_79), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_52), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_151), .Y(n_350) );
CKINVDCx11_ASAP7_75t_R g351 ( .A(n_56), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_219), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_11), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_200), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_18), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_60), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_48), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_169), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_229), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_41), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_48), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_81), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_65), .Y(n_363) );
INVxp67_ASAP7_75t_L g364 ( .A(n_102), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_64), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_120), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_203), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_134), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_76), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_84), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_30), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_39), .Y(n_372) );
INVxp33_ASAP7_75t_L g373 ( .A(n_174), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_21), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_32), .Y(n_375) );
INVxp33_ASAP7_75t_SL g376 ( .A(n_196), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_308), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_372), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_305), .B(n_3), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_246), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_308), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_246), .B(n_3), .Y(n_382) );
NAND2xp5_ASAP7_75t_SL g383 ( .A(n_305), .B(n_4), .Y(n_383) );
BUFx2_ASAP7_75t_L g384 ( .A(n_320), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_320), .A2(n_4), .B1(n_6), .B2(n_7), .Y(n_385) );
INVx3_ASAP7_75t_L g386 ( .A(n_246), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_251), .B(n_6), .Y(n_387) );
AND2x2_ASAP7_75t_SL g388 ( .A(n_283), .B(n_75), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_263), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_345), .B(n_9), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_359), .B(n_10), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_256), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_256), .Y(n_394) );
OA21x2_ASAP7_75t_L g395 ( .A1(n_259), .A2(n_12), .B(n_13), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_308), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_349), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_349), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_242), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_346), .B(n_12), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_259), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_308), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_242), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_373), .B(n_15), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_308), .Y(n_405) );
OAI22xp5_ASAP7_75t_SL g406 ( .A1(n_254), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_244), .Y(n_407) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_351), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_323), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_308), .Y(n_410) );
INVx2_ASAP7_75t_SL g411 ( .A(n_266), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_253), .B(n_16), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_382), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_380), .B(n_373), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_380), .Y(n_416) );
BUFx3_ASAP7_75t_L g417 ( .A(n_382), .Y(n_417) );
INVx4_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_382), .B(n_268), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_395), .A2(n_265), .B1(n_273), .B2(n_261), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_384), .B(n_267), .Y(n_422) );
INVx4_ASAP7_75t_L g423 ( .A(n_382), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_377), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_377), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_384), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_386), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_381), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_395), .A2(n_277), .B1(n_278), .B2(n_276), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
NOR2x1p5_ASAP7_75t_L g432 ( .A(n_391), .B(n_267), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_380), .B(n_268), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_409), .B(n_302), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_409), .B(n_404), .Y(n_435) );
AND2x2_ASAP7_75t_SL g436 ( .A(n_388), .B(n_316), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_380), .B(n_285), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_386), .B(n_279), .Y(n_438) );
NOR2x1p5_ASAP7_75t_L g439 ( .A(n_391), .B(n_243), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_409), .B(n_257), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_395), .A2(n_287), .B1(n_297), .B2(n_295), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_381), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_404), .B(n_243), .Y(n_443) );
INVx4_ASAP7_75t_L g444 ( .A(n_386), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_411), .B(n_255), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_392), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_411), .B(n_255), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_386), .B(n_257), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_386), .Y(n_449) );
INVx3_ASAP7_75t_L g450 ( .A(n_381), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_387), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_388), .A2(n_263), .B1(n_284), .B2(n_275), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_399), .Y(n_453) );
OR2x6_ASAP7_75t_L g454 ( .A(n_389), .B(n_306), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_411), .B(n_260), .Y(n_455) );
NOR2x1p5_ASAP7_75t_L g456 ( .A(n_392), .B(n_408), .Y(n_456) );
CKINVDCx11_ASAP7_75t_R g457 ( .A(n_408), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_402), .Y(n_458) );
INVx4_ASAP7_75t_L g459 ( .A(n_387), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_454), .B(n_406), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_418), .B(n_388), .Y(n_461) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_436), .A2(n_388), .B1(n_387), .B2(n_383), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_448), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_436), .A2(n_387), .B1(n_395), .B2(n_407), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_446), .B(n_387), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_418), .B(n_402), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_457), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_440), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_436), .A2(n_395), .B1(n_407), .B2(n_383), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_446), .B(n_400), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_444), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_418), .B(n_402), .Y(n_473) );
BUFx3_ASAP7_75t_L g474 ( .A(n_414), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_422), .B(n_379), .Y(n_475) );
AOI22xp5_ASAP7_75t_SL g476 ( .A1(n_434), .A2(n_254), .B1(n_361), .B2(n_389), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_415), .B(n_403), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_427), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_448), .B(n_403), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_422), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_434), .B(n_264), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_422), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_427), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_423), .B(n_396), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_436), .A2(n_385), .B1(n_275), .B2(n_328), .Y(n_485) );
NAND2xp33_ASAP7_75t_L g486 ( .A(n_420), .B(n_260), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_455), .B(n_403), .Y(n_487) );
INVx5_ASAP7_75t_L g488 ( .A(n_423), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_452), .A2(n_385), .B1(n_361), .B2(n_284), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_444), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_451), .A2(n_395), .B1(n_394), .B2(n_412), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_434), .B(n_264), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_423), .B(n_396), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_423), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_428), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_451), .A2(n_394), .B1(n_397), .B2(n_393), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_435), .A2(n_329), .B1(n_342), .B2(n_328), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_449), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_455), .B(n_394), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_440), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_449), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_449), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_449), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_445), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_445), .Y(n_506) );
OAI21xp5_ASAP7_75t_L g507 ( .A1(n_442), .A2(n_410), .B(n_405), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_414), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_435), .A2(n_342), .B1(n_343), .B2(n_329), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_423), .B(n_405), .Y(n_510) );
NOR2x1p5_ASAP7_75t_L g511 ( .A(n_445), .B(n_290), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_459), .A2(n_394), .B1(n_397), .B2(n_393), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_435), .B(n_398), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g514 ( .A(n_457), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_459), .A2(n_398), .B1(n_338), .B2(n_376), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_459), .A2(n_338), .B1(n_376), .B2(n_269), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_459), .A2(n_269), .B1(n_410), .B2(n_405), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_414), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_439), .B(n_378), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_447), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_431), .B(n_319), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_431), .B(n_298), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_414), .Y(n_524) );
O2A1O1Ixp5_ASAP7_75t_L g525 ( .A1(n_419), .A2(n_252), .B(n_249), .C(n_245), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_443), .B(n_290), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_443), .B(n_334), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_438), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_438), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_452), .A2(n_362), .B1(n_343), .B2(n_299), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_439), .B(n_378), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_459), .B(n_364), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_438), .B(n_350), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_417), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_417), .B(n_352), .Y(n_535) );
NAND3xp33_ASAP7_75t_SL g536 ( .A(n_462), .B(n_362), .C(n_355), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_498), .B(n_454), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_528), .Y(n_538) );
NOR3xp33_ASAP7_75t_L g539 ( .A(n_489), .B(n_406), .C(n_351), .Y(n_539) );
NOR2xp67_ASAP7_75t_L g540 ( .A(n_485), .B(n_420), .Y(n_540) );
BUFx8_ASAP7_75t_SL g541 ( .A(n_467), .Y(n_541) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_505), .A2(n_454), .B(n_437), .C(n_433), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_466), .A2(n_416), .B(n_430), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_464), .A2(n_454), .B1(n_430), .B2(n_441), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_483), .B(n_432), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_480), .B(n_454), .Y(n_546) );
OR2x6_ASAP7_75t_SL g547 ( .A(n_467), .B(n_514), .Y(n_547) );
NAND2x1p5_ASAP7_75t_L g548 ( .A(n_483), .B(n_432), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_471), .B(n_437), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_506), .A2(n_454), .B1(n_401), .B2(n_272), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_529), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_530), .B(n_468), .C(n_481), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_480), .B(n_355), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_461), .A2(n_456), .B1(n_450), .B2(n_421), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_500), .Y(n_556) );
BUFx3_ASAP7_75t_L g557 ( .A(n_519), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_463), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_482), .B(n_456), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_461), .A2(n_450), .B1(n_421), .B2(n_424), .Y(n_560) );
AOI221xp5_ASAP7_75t_L g561 ( .A1(n_521), .A2(n_318), .B1(n_371), .B2(n_314), .C(n_274), .Y(n_561) );
O2A1O1Ixp33_ASAP7_75t_L g562 ( .A1(n_513), .A2(n_313), .B(n_322), .C(n_300), .Y(n_562) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_509), .B(n_325), .Y(n_563) );
AOI21x1_ASAP7_75t_L g564 ( .A1(n_479), .A2(n_424), .B(n_413), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_495), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_470), .A2(n_401), .B1(n_326), .B2(n_333), .Y(n_566) );
O2A1O1Ixp5_ASAP7_75t_L g567 ( .A1(n_525), .A2(n_413), .B(n_426), .C(n_425), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_473), .A2(n_425), .B(n_413), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_493), .B(n_247), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_482), .B(n_330), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_495), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_488), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_495), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_465), .B(n_450), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_534), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_501), .B(n_301), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
BUFx2_ASAP7_75t_L g578 ( .A(n_475), .Y(n_578) );
NOR2xp33_ASAP7_75t_R g579 ( .A(n_486), .B(n_352), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_475), .B(n_527), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_534), .Y(n_581) );
NOR2xp33_ASAP7_75t_SL g582 ( .A(n_488), .B(n_426), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_534), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_475), .B(n_458), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_476), .B(n_339), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_516), .B(n_429), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_522), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_519), .B(n_429), .Y(n_588) );
INVxp67_ASAP7_75t_L g589 ( .A(n_511), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_484), .A2(n_458), .B(n_410), .Y(n_590) );
INVx4_ASAP7_75t_L g591 ( .A(n_534), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_523), .B(n_360), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_519), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_518), .Y(n_594) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_474), .Y(n_595) );
A2O1A1Ixp33_ASAP7_75t_SL g596 ( .A1(n_535), .A2(n_401), .B(n_390), .C(n_289), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_460), .A2(n_401), .B1(n_344), .B2(n_347), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_460), .A2(n_401), .B1(n_353), .B2(n_356), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_508), .B(n_270), .Y(n_599) );
OR2x6_ASAP7_75t_SL g600 ( .A(n_460), .B(n_363), .Y(n_600) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_533), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_474), .Y(n_602) );
NOR3xp33_ASAP7_75t_SL g603 ( .A(n_460), .B(n_375), .C(n_374), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_531), .B(n_390), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g605 ( .A(n_508), .B(n_271), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_486), .A2(n_357), .B1(n_365), .B2(n_340), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_531), .Y(n_607) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_507), .A2(n_289), .B(n_285), .Y(n_608) );
BUFx6f_ASAP7_75t_L g609 ( .A(n_469), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_494), .A2(n_453), .B(n_280), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_515), .Y(n_611) );
BUFx3_ASAP7_75t_L g612 ( .A(n_491), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_518), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_532), .A2(n_258), .B1(n_286), .B2(n_282), .Y(n_614) );
NAND2xp5_ASAP7_75t_SL g615 ( .A(n_469), .B(n_281), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_510), .A2(n_453), .B(n_291), .Y(n_616) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_487), .A2(n_293), .B(n_294), .C(n_288), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_491), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_472), .B(n_304), .Y(n_619) );
INVx5_ASAP7_75t_L g620 ( .A(n_472), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_517), .B(n_17), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_524), .A2(n_307), .B1(n_310), .B2(n_309), .Y(n_622) );
O2A1O1Ixp33_ASAP7_75t_L g623 ( .A1(n_477), .A2(n_312), .B(n_315), .C(n_311), .Y(n_623) );
BUFx8_ASAP7_75t_SL g624 ( .A(n_496), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g625 ( .A1(n_524), .A2(n_321), .B1(n_327), .B2(n_324), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_497), .B(n_331), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_496), .B(n_19), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_492), .A2(n_248), .B1(n_335), .B2(n_332), .Y(n_628) );
AOI21x1_ASAP7_75t_L g629 ( .A1(n_502), .A2(n_250), .B(n_337), .Y(n_629) );
INVx5_ASAP7_75t_L g630 ( .A(n_490), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_512), .B(n_367), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_504), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_503), .A2(n_358), .B(n_368), .C(n_348), .Y(n_633) );
O2A1O1Ixp33_ASAP7_75t_SL g634 ( .A1(n_499), .A2(n_262), .B(n_292), .C(n_366), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_466), .A2(n_303), .B(n_296), .Y(n_635) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_572), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_604), .Y(n_637) );
AND2x4_ASAP7_75t_L g638 ( .A(n_552), .B(n_303), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_543), .A2(n_336), .B(n_317), .Y(n_639) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_568), .A2(n_336), .B(n_317), .Y(n_640) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_572), .Y(n_641) );
OAI21x1_ASAP7_75t_L g642 ( .A1(n_608), .A2(n_354), .B(n_341), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_611), .B(n_22), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_564), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_542), .A2(n_370), .B(n_369), .C(n_341), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_580), .B(n_553), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_609), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_624), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_540), .B(n_22), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_577), .Y(n_650) );
AO21x1_ASAP7_75t_L g651 ( .A1(n_628), .A2(n_399), .B(n_78), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_539), .A2(n_399), .B1(n_24), .B2(n_25), .C(n_26), .Y(n_652) );
AO31x2_ASAP7_75t_L g653 ( .A1(n_566), .A2(n_23), .A3(n_24), .B(n_26), .Y(n_653) );
O2A1O1Ixp33_ASAP7_75t_L g654 ( .A1(n_550), .A2(n_23), .B(n_27), .C(n_30), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_584), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_609), .Y(n_656) );
OAI22x1_ASAP7_75t_L g657 ( .A1(n_600), .A2(n_27), .B1(n_31), .B2(n_32), .Y(n_657) );
BUFx10_ASAP7_75t_L g658 ( .A(n_545), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_596), .A2(n_129), .B(n_240), .C(n_239), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_537), .B(n_31), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_587), .A2(n_33), .B1(n_34), .B2(n_35), .C(n_36), .Y(n_661) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_592), .B(n_33), .C(n_34), .Y(n_662) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_541), .B(n_35), .Y(n_663) );
INVx3_ASAP7_75t_L g664 ( .A(n_557), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_549), .B(n_37), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_546), .B(n_578), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_550), .A2(n_38), .B(n_40), .C(n_41), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_601), .B(n_40), .Y(n_668) );
INVx3_ASAP7_75t_L g669 ( .A(n_545), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_570), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_563), .A2(n_43), .B1(n_44), .B2(n_45), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_556), .B(n_43), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_570), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_589), .B(n_45), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_588), .Y(n_675) );
AO31x2_ASAP7_75t_L g676 ( .A1(n_566), .A2(n_46), .A3(n_49), .B(n_50), .Y(n_676) );
OAI21x1_ASAP7_75t_L g677 ( .A1(n_610), .A2(n_88), .B(n_86), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_561), .A2(n_46), .B1(n_49), .B2(n_50), .C(n_51), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_558), .Y(n_679) );
NAND2x1p5_ASAP7_75t_L g680 ( .A(n_591), .B(n_53), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_597), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_681) );
NOR2x1p5_ASAP7_75t_L g682 ( .A(n_536), .B(n_54), .Y(n_682) );
INVx4_ASAP7_75t_L g683 ( .A(n_595), .Y(n_683) );
CKINVDCx6p67_ASAP7_75t_R g684 ( .A(n_547), .Y(n_684) );
AO21x2_ASAP7_75t_L g685 ( .A1(n_579), .A2(n_91), .B(n_90), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_585), .A2(n_55), .B1(n_57), .B2(n_58), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_562), .A2(n_57), .B(n_58), .C(n_60), .Y(n_687) );
NOR2xp33_ASAP7_75t_SL g688 ( .A(n_582), .B(n_61), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_576), .Y(n_689) );
AO32x2_ASAP7_75t_L g690 ( .A1(n_597), .A2(n_61), .A3(n_62), .B1(n_63), .B2(n_64), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_590), .A2(n_152), .B(n_237), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_619), .Y(n_692) );
NAND2xp33_ASAP7_75t_L g693 ( .A(n_544), .B(n_92), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g694 ( .A1(n_598), .A2(n_66), .B(n_67), .C(n_68), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_619), .Y(n_695) );
INVx3_ASAP7_75t_SL g696 ( .A(n_607), .Y(n_696) );
CKINVDCx16_ASAP7_75t_R g697 ( .A(n_598), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_593), .Y(n_698) );
BUFx2_ASAP7_75t_L g699 ( .A(n_595), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_569), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_544), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_559), .B(n_69), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_538), .Y(n_703) );
INVx2_ASAP7_75t_L g704 ( .A(n_594), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_551), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_621), .A2(n_70), .B1(n_71), .B2(n_72), .Y(n_706) );
NOR2x1_ASAP7_75t_R g707 ( .A(n_559), .B(n_71), .Y(n_707) );
O2A1O1Ixp33_ASAP7_75t_L g708 ( .A1(n_633), .A2(n_73), .B(n_74), .C(n_93), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_548), .B(n_73), .Y(n_709) );
AO31x2_ASAP7_75t_L g710 ( .A1(n_635), .A2(n_98), .A3(n_99), .B(n_100), .Y(n_710) );
AOI31xp67_ASAP7_75t_L g711 ( .A1(n_575), .A2(n_105), .A3(n_106), .B(n_108), .Y(n_711) );
O2A1O1Ixp33_ASAP7_75t_L g712 ( .A1(n_586), .A2(n_111), .B(n_112), .C(n_113), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g713 ( .A1(n_606), .A2(n_114), .B(n_115), .C(n_117), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_554), .A2(n_119), .B(n_121), .Y(n_714) );
AO31x2_ASAP7_75t_L g715 ( .A1(n_616), .A2(n_125), .A3(n_126), .B(n_127), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_555), .B(n_132), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_548), .B(n_133), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_614), .A2(n_142), .B1(n_143), .B2(n_144), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_627), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_574), .A2(n_146), .B1(n_147), .B2(n_154), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_560), .A2(n_157), .B(n_158), .Y(n_721) );
AO31x2_ASAP7_75t_L g722 ( .A1(n_581), .A2(n_160), .A3(n_161), .B(n_162), .Y(n_722) );
OAI22x1_ASAP7_75t_L g723 ( .A1(n_603), .A2(n_163), .B1(n_164), .B2(n_165), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_565), .Y(n_724) );
AO31x2_ASAP7_75t_L g725 ( .A1(n_583), .A2(n_170), .A3(n_172), .B(n_173), .Y(n_725) );
OAI22xp33_ASAP7_75t_L g726 ( .A1(n_622), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_726) );
NAND2x1p5_ASAP7_75t_L g727 ( .A(n_602), .B(n_178), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g728 ( .A1(n_626), .A2(n_179), .B1(n_180), .B2(n_183), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_571), .Y(n_729) );
OAI21xp5_ASAP7_75t_L g730 ( .A1(n_573), .A2(n_185), .B(n_186), .Y(n_730) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_613), .A2(n_187), .B(n_188), .Y(n_731) );
AO31x2_ASAP7_75t_L g732 ( .A1(n_631), .A2(n_189), .A3(n_190), .B(n_192), .Y(n_732) );
AO31x2_ASAP7_75t_L g733 ( .A1(n_634), .A2(n_195), .A3(n_197), .B(n_198), .Y(n_733) );
BUFx3_ASAP7_75t_L g734 ( .A(n_620), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_620), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_615), .A2(n_199), .B(n_201), .Y(n_736) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_599), .A2(n_202), .B(n_204), .C(n_206), .Y(n_737) );
AO32x2_ASAP7_75t_L g738 ( .A1(n_625), .A2(n_210), .A3(n_217), .B1(n_218), .B2(n_220), .Y(n_738) );
BUFx3_ASAP7_75t_L g739 ( .A(n_620), .Y(n_739) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_630), .A2(n_221), .B1(n_222), .B2(n_228), .Y(n_740) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_605), .A2(n_231), .B(n_233), .C(n_235), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_618), .B(n_241), .Y(n_742) );
AND2x4_ASAP7_75t_L g743 ( .A(n_630), .B(n_612), .Y(n_743) );
INVx2_ASAP7_75t_SL g744 ( .A(n_630), .Y(n_744) );
OAI21xp5_ASAP7_75t_L g745 ( .A1(n_632), .A2(n_543), .B(n_567), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_632), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g747 ( .A1(n_632), .A2(n_542), .B(n_617), .C(n_623), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_703), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_697), .B(n_700), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_646), .B(n_692), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_705), .Y(n_751) );
INVx3_ASAP7_75t_L g752 ( .A(n_743), .Y(n_752) );
AO31x2_ASAP7_75t_L g753 ( .A1(n_651), .A2(n_645), .A3(n_639), .B(n_747), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_679), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_650), .B(n_638), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_734), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_696), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_695), .B(n_655), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_702), .B(n_638), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_689), .B(n_637), .Y(n_760) );
OR2x6_ASAP7_75t_L g761 ( .A(n_648), .B(n_680), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_640), .A2(n_659), .B(n_665), .Y(n_762) );
OA21x2_ASAP7_75t_L g763 ( .A1(n_731), .A2(n_730), .B(n_677), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_672), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_684), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g766 ( .A1(n_649), .A2(n_719), .B(n_721), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_660), .A2(n_643), .B1(n_682), .B2(n_670), .Y(n_767) );
NOR2x1_ASAP7_75t_L g768 ( .A(n_739), .B(n_662), .Y(n_768) );
HB1xp67_ASAP7_75t_L g769 ( .A(n_743), .Y(n_769) );
AOI21xp33_ASAP7_75t_L g770 ( .A1(n_654), .A2(n_667), .B(n_687), .Y(n_770) );
OAI221xp5_ASAP7_75t_SL g771 ( .A1(n_671), .A2(n_652), .B1(n_686), .B2(n_678), .C(n_681), .Y(n_771) );
AND2x2_ASAP7_75t_L g772 ( .A(n_657), .B(n_673), .Y(n_772) );
INVxp67_ASAP7_75t_L g773 ( .A(n_707), .Y(n_773) );
BUFx2_ASAP7_75t_L g774 ( .A(n_744), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_704), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_675), .B(n_666), .Y(n_776) );
AND2x2_ASAP7_75t_L g777 ( .A(n_669), .B(n_658), .Y(n_777) );
AO31x2_ASAP7_75t_L g778 ( .A1(n_701), .A2(n_723), .A3(n_720), .B(n_713), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g779 ( .A1(n_742), .A2(n_706), .B1(n_727), .B2(n_661), .Y(n_779) );
A2O1A1Ixp33_ASAP7_75t_L g780 ( .A1(n_708), .A2(n_694), .B(n_717), .C(n_709), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_658), .B(n_698), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_668), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_724), .B(n_729), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_664), .B(n_674), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_735), .B(n_746), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g786 ( .A(n_688), .B(n_636), .Y(n_786) );
A2O1A1Ixp33_ASAP7_75t_L g787 ( .A1(n_737), .A2(n_741), .B(n_712), .C(n_714), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_653), .Y(n_788) );
A2O1A1Ixp33_ASAP7_75t_L g789 ( .A1(n_728), .A2(n_736), .B(n_716), .C(n_691), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_647), .B(n_656), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_699), .B(n_641), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_641), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_663), .A2(n_683), .B1(n_718), .B2(n_726), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_740), .A2(n_685), .B(n_683), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_690), .Y(n_795) );
OR2x2_ASAP7_75t_L g796 ( .A(n_676), .B(n_732), .Y(n_796) );
AO21x2_ASAP7_75t_L g797 ( .A1(n_711), .A2(n_733), .B(n_732), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_733), .B(n_732), .Y(n_798) );
OR2x6_ASAP7_75t_L g799 ( .A(n_690), .B(n_738), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_733), .B(n_715), .Y(n_800) );
A2O1A1Ixp33_ASAP7_75t_L g801 ( .A1(n_738), .A2(n_710), .B(n_722), .C(n_725), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_710), .B(n_722), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_710), .B(n_722), .Y(n_803) );
AND2x4_ASAP7_75t_L g804 ( .A(n_725), .B(n_743), .Y(n_804) );
OAI21xp33_ASAP7_75t_L g805 ( .A1(n_646), .A2(n_483), .B(n_478), .Y(n_805) );
NAND2x1p5_ASAP7_75t_L g806 ( .A(n_734), .B(n_739), .Y(n_806) );
OAI21xp5_ASAP7_75t_L g807 ( .A1(n_646), .A2(n_544), .B(n_542), .Y(n_807) );
NOR2xp67_ASAP7_75t_SL g808 ( .A(n_697), .B(n_478), .Y(n_808) );
AND2x2_ASAP7_75t_L g809 ( .A(n_697), .B(n_446), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_646), .B(n_692), .Y(n_810) );
AND2x4_ASAP7_75t_L g811 ( .A(n_743), .B(n_734), .Y(n_811) );
AOI21xp33_ASAP7_75t_L g812 ( .A1(n_693), .A2(n_649), .B(n_628), .Y(n_812) );
AOI21x1_ASAP7_75t_L g813 ( .A1(n_644), .A2(n_629), .B(n_642), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_646), .B(n_692), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_703), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_650), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_697), .B(n_446), .Y(n_817) );
BUFx2_ASAP7_75t_L g818 ( .A(n_689), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_703), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g820 ( .A1(n_697), .A2(n_550), .B1(n_695), .B2(n_692), .Y(n_820) );
OAI21xp5_ASAP7_75t_L g821 ( .A1(n_646), .A2(n_544), .B(n_542), .Y(n_821) );
NOR2xp33_ASAP7_75t_SL g822 ( .A(n_697), .B(n_688), .Y(n_822) );
BUFx3_ASAP7_75t_L g823 ( .A(n_696), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_646), .B(n_692), .Y(n_824) );
BUFx2_ASAP7_75t_SL g825 ( .A(n_689), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_646), .B(n_692), .Y(n_826) );
AND2x4_ASAP7_75t_L g827 ( .A(n_743), .B(n_734), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_703), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g829 ( .A(n_684), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_693), .A2(n_745), .B(n_544), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_697), .A2(n_539), .B1(n_460), .B2(n_563), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_703), .Y(n_832) );
INVxp67_ASAP7_75t_L g833 ( .A(n_707), .Y(n_833) );
AND2x4_ASAP7_75t_L g834 ( .A(n_743), .B(n_734), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_703), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_646), .B(n_692), .Y(n_836) );
AOI21x1_ASAP7_75t_L g837 ( .A1(n_644), .A2(n_629), .B(n_642), .Y(n_837) );
BUFx3_ASAP7_75t_L g838 ( .A(n_696), .Y(n_838) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_693), .A2(n_745), .B(n_544), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_697), .B(n_552), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_697), .B(n_446), .Y(n_841) );
BUFx8_ASAP7_75t_L g842 ( .A(n_700), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_697), .B(n_446), .Y(n_843) );
NOR2xp33_ASAP7_75t_SL g844 ( .A(n_697), .B(n_688), .Y(n_844) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_707), .A2(n_563), .B1(n_406), .B2(n_489), .C1(n_530), .C2(n_520), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_646), .B(n_692), .Y(n_846) );
AND2x4_ASAP7_75t_L g847 ( .A(n_752), .B(n_811), .Y(n_847) );
OR2x2_ASAP7_75t_L g848 ( .A(n_820), .B(n_809), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_817), .B(n_841), .Y(n_849) );
INVx8_ASAP7_75t_L g850 ( .A(n_811), .Y(n_850) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_822), .Y(n_851) );
INVx1_ASAP7_75t_L g852 ( .A(n_788), .Y(n_852) );
OA21x2_ASAP7_75t_L g853 ( .A1(n_801), .A2(n_798), .B(n_800), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_845), .B(n_843), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_750), .B(n_810), .Y(n_855) );
OR2x2_ASAP7_75t_L g856 ( .A(n_820), .B(n_840), .Y(n_856) );
INVx3_ASAP7_75t_SL g857 ( .A(n_761), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_783), .Y(n_858) );
BUFx4f_ASAP7_75t_SL g859 ( .A(n_829), .Y(n_859) );
AO21x2_ASAP7_75t_L g860 ( .A1(n_800), .A2(n_797), .B(n_839), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g861 ( .A1(n_831), .A2(n_770), .B1(n_767), .B2(n_771), .C(n_782), .Y(n_861) );
AOI222xp33_ASAP7_75t_L g862 ( .A1(n_773), .A2(n_833), .B1(n_808), .B2(n_749), .C1(n_846), .C2(n_826), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_783), .Y(n_863) );
AO21x2_ASAP7_75t_L g864 ( .A1(n_797), .A2(n_830), .B(n_802), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_748), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_845), .B(n_750), .Y(n_866) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_822), .Y(n_867) );
AND2x4_ASAP7_75t_L g868 ( .A(n_752), .B(n_827), .Y(n_868) );
AND2x2_ASAP7_75t_L g869 ( .A(n_810), .B(n_814), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_751), .Y(n_870) );
AND2x2_ASAP7_75t_L g871 ( .A(n_814), .B(n_824), .Y(n_871) );
AND2x4_ASAP7_75t_L g872 ( .A(n_827), .B(n_834), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_844), .A2(n_770), .B1(n_805), .B2(n_772), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_815), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_775), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_844), .A2(n_779), .B1(n_760), .B2(n_764), .Y(n_876) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_816), .Y(n_877) );
HB1xp67_ASAP7_75t_L g878 ( .A(n_755), .Y(n_878) );
OR2x2_ASAP7_75t_L g879 ( .A(n_824), .B(n_826), .Y(n_879) );
INVx2_ASAP7_75t_SL g880 ( .A(n_806), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_765), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_819), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_836), .B(n_846), .Y(n_883) );
OA21x2_ASAP7_75t_L g884 ( .A1(n_803), .A2(n_796), .B(n_762), .Y(n_884) );
INVx1_ASAP7_75t_L g885 ( .A(n_828), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_832), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_842), .Y(n_887) );
AND2x4_ASAP7_75t_L g888 ( .A(n_834), .B(n_792), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_835), .Y(n_889) );
INVx4_ASAP7_75t_L g890 ( .A(n_761), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_836), .Y(n_891) );
BUFx3_ASAP7_75t_L g892 ( .A(n_806), .Y(n_892) );
OR2x2_ASAP7_75t_L g893 ( .A(n_776), .B(n_758), .Y(n_893) );
AO21x2_ASAP7_75t_L g894 ( .A1(n_812), .A2(n_794), .B(n_837), .Y(n_894) );
AO21x2_ASAP7_75t_L g895 ( .A1(n_813), .A2(n_821), .B(n_807), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_776), .B(n_758), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_754), .B(n_759), .Y(n_897) );
INVx1_ASAP7_75t_L g898 ( .A(n_799), .Y(n_898) );
INVx2_ASAP7_75t_SL g899 ( .A(n_761), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_799), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_799), .Y(n_901) );
OA21x2_ASAP7_75t_L g902 ( .A1(n_766), .A2(n_821), .B(n_807), .Y(n_902) );
INVx2_ASAP7_75t_L g903 ( .A(n_790), .Y(n_903) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_842), .Y(n_904) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_779), .A2(n_825), .B1(n_793), .B2(n_818), .Y(n_905) );
INVx2_ASAP7_75t_L g906 ( .A(n_790), .Y(n_906) );
AOI21xp5_ASAP7_75t_SL g907 ( .A1(n_786), .A2(n_804), .B(n_763), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_784), .A2(n_795), .B1(n_781), .B2(n_766), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_777), .B(n_769), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_785), .B(n_780), .Y(n_910) );
AO21x2_ASAP7_75t_L g911 ( .A1(n_787), .A2(n_789), .B(n_804), .Y(n_911) );
BUFx2_ASAP7_75t_L g912 ( .A(n_791), .Y(n_912) );
BUFx2_ASAP7_75t_SL g913 ( .A(n_757), .Y(n_913) );
OAI211xp5_ASAP7_75t_L g914 ( .A1(n_774), .A2(n_768), .B(n_756), .C(n_823), .Y(n_914) );
OR2x2_ASAP7_75t_L g915 ( .A(n_753), .B(n_778), .Y(n_915) );
AND2x2_ASAP7_75t_L g916 ( .A(n_753), .B(n_778), .Y(n_916) );
BUFx3_ASAP7_75t_L g917 ( .A(n_838), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_753), .B(n_778), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g919 ( .A1(n_845), .A2(n_697), .B1(n_539), .B2(n_689), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_788), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_845), .B(n_563), .Y(n_921) );
AND2x2_ASAP7_75t_L g922 ( .A(n_809), .B(n_697), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_811), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_852), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_855), .B(n_869), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_855), .B(n_869), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_871), .B(n_898), .Y(n_927) );
AND2x4_ASAP7_75t_L g928 ( .A(n_898), .B(n_900), .Y(n_928) );
OR2x2_ASAP7_75t_L g929 ( .A(n_848), .B(n_856), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_871), .B(n_900), .Y(n_930) );
HB1xp67_ASAP7_75t_L g931 ( .A(n_877), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_901), .B(n_849), .Y(n_932) );
OR2x2_ASAP7_75t_L g933 ( .A(n_848), .B(n_856), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_881), .Y(n_934) );
NOR2x1p5_ASAP7_75t_L g935 ( .A(n_851), .B(n_867), .Y(n_935) );
INVxp67_ASAP7_75t_L g936 ( .A(n_912), .Y(n_936) );
AND2x2_ASAP7_75t_L g937 ( .A(n_901), .B(n_849), .Y(n_937) );
BUFx2_ASAP7_75t_L g938 ( .A(n_912), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_920), .Y(n_939) );
OR2x2_ASAP7_75t_L g940 ( .A(n_879), .B(n_883), .Y(n_940) );
AND2x2_ASAP7_75t_L g941 ( .A(n_916), .B(n_918), .Y(n_941) );
BUFx3_ASAP7_75t_L g942 ( .A(n_850), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_865), .Y(n_943) );
INVxp67_ASAP7_75t_L g944 ( .A(n_913), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_878), .Y(n_945) );
BUFx4f_ASAP7_75t_SL g946 ( .A(n_857), .Y(n_946) );
INVx1_ASAP7_75t_SL g947 ( .A(n_893), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_916), .B(n_918), .Y(n_948) );
NAND2xp5_ASAP7_75t_SL g949 ( .A(n_890), .B(n_862), .Y(n_949) );
INVx4_ASAP7_75t_L g950 ( .A(n_850), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_865), .Y(n_951) );
NOR2x1_ASAP7_75t_L g952 ( .A(n_890), .B(n_914), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_870), .Y(n_953) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_893), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_870), .Y(n_955) );
INVx2_ASAP7_75t_SL g956 ( .A(n_892), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_891), .B(n_879), .Y(n_957) );
INVxp67_ASAP7_75t_SL g958 ( .A(n_896), .Y(n_958) );
OR2x2_ASAP7_75t_L g959 ( .A(n_883), .B(n_896), .Y(n_959) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_919), .B(n_866), .Y(n_960) );
AND2x4_ASAP7_75t_L g961 ( .A(n_911), .B(n_915), .Y(n_961) );
NOR3xp33_ASAP7_75t_SL g962 ( .A(n_921), .B(n_881), .C(n_861), .Y(n_962) );
INVx5_ASAP7_75t_L g963 ( .A(n_890), .Y(n_963) );
AND2x2_ASAP7_75t_L g964 ( .A(n_902), .B(n_903), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_891), .B(n_902), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_902), .B(n_903), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g967 ( .A(n_859), .Y(n_967) );
AND2x2_ASAP7_75t_L g968 ( .A(n_906), .B(n_910), .Y(n_968) );
AND2x4_ASAP7_75t_L g969 ( .A(n_911), .B(n_915), .Y(n_969) );
INVx1_ASAP7_75t_L g970 ( .A(n_874), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_910), .B(n_863), .Y(n_971) );
AND2x2_ASAP7_75t_L g972 ( .A(n_882), .B(n_886), .Y(n_972) );
INVx2_ASAP7_75t_L g973 ( .A(n_924), .Y(n_973) );
BUFx2_ASAP7_75t_L g974 ( .A(n_944), .Y(n_974) );
OR2x2_ASAP7_75t_L g975 ( .A(n_947), .B(n_922), .Y(n_975) );
AND2x4_ASAP7_75t_SL g976 ( .A(n_950), .B(n_872), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_947), .B(n_885), .Y(n_977) );
AND2x2_ASAP7_75t_L g978 ( .A(n_941), .B(n_864), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_941), .B(n_864), .Y(n_979) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_967), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_958), .B(n_885), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_972), .Y(n_982) );
INVx4_ASAP7_75t_L g983 ( .A(n_963), .Y(n_983) );
NOR2xp33_ASAP7_75t_L g984 ( .A(n_960), .B(n_854), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_972), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_943), .Y(n_986) );
AND2x2_ASAP7_75t_SL g987 ( .A(n_938), .B(n_950), .Y(n_987) );
AND2x4_ASAP7_75t_L g988 ( .A(n_928), .B(n_911), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_925), .B(n_882), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_925), .B(n_926), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_926), .B(n_889), .Y(n_991) );
AND2x2_ASAP7_75t_L g992 ( .A(n_948), .B(n_864), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_943), .Y(n_993) );
OR2x2_ASAP7_75t_L g994 ( .A(n_940), .B(n_922), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_948), .B(n_895), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_954), .B(n_886), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_927), .B(n_889), .Y(n_997) );
AND2x2_ASAP7_75t_L g998 ( .A(n_930), .B(n_895), .Y(n_998) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_940), .B(n_858), .Y(n_999) );
AND2x2_ASAP7_75t_L g1000 ( .A(n_932), .B(n_895), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_932), .B(n_853), .Y(n_1001) );
NAND2xp5_ASAP7_75t_SL g1002 ( .A(n_952), .B(n_873), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_951), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_951), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_953), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_928), .B(n_860), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_953), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_955), .Y(n_1008) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_937), .B(n_853), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1010 ( .A(n_937), .B(n_853), .Y(n_1010) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_959), .B(n_897), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_952), .A2(n_907), .B(n_894), .Y(n_1012) );
NAND4xp25_ASAP7_75t_L g1013 ( .A(n_949), .B(n_905), .C(n_876), .D(n_908), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_955), .Y(n_1014) );
OR2x2_ASAP7_75t_L g1015 ( .A(n_945), .B(n_875), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_964), .B(n_853), .Y(n_1016) );
AND2x4_ASAP7_75t_L g1017 ( .A(n_928), .B(n_860), .Y(n_1017) );
NOR2xp33_ASAP7_75t_R g1018 ( .A(n_946), .B(n_857), .Y(n_1018) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_931), .B(n_875), .Y(n_1019) );
NOR3xp33_ASAP7_75t_L g1020 ( .A(n_956), .B(n_899), .C(n_904), .Y(n_1020) );
NOR2x1_ASAP7_75t_L g1021 ( .A(n_950), .B(n_913), .Y(n_1021) );
AND2x2_ASAP7_75t_SL g1022 ( .A(n_950), .B(n_887), .Y(n_1022) );
AND2x2_ASAP7_75t_L g1023 ( .A(n_964), .B(n_884), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_966), .B(n_884), .Y(n_1024) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_957), .B(n_899), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_966), .B(n_884), .Y(n_1026) );
OR2x2_ASAP7_75t_L g1027 ( .A(n_929), .B(n_917), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_990), .B(n_929), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_978), .B(n_961), .Y(n_1029) );
INVx2_ASAP7_75t_L g1030 ( .A(n_973), .Y(n_1030) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_982), .B(n_968), .Y(n_1031) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_985), .B(n_968), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1033 ( .A(n_979), .B(n_961), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_989), .B(n_971), .Y(n_1034) );
NOR2xp33_ASAP7_75t_L g1035 ( .A(n_984), .B(n_917), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_979), .B(n_961), .Y(n_1036) );
INVx1_ASAP7_75t_L g1037 ( .A(n_986), .Y(n_1037) );
OR2x2_ASAP7_75t_L g1038 ( .A(n_992), .B(n_933), .Y(n_1038) );
INVxp67_ASAP7_75t_L g1039 ( .A(n_974), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_993), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1003), .Y(n_1041) );
AND2x2_ASAP7_75t_L g1042 ( .A(n_992), .B(n_961), .Y(n_1042) );
NOR2xp33_ASAP7_75t_L g1043 ( .A(n_984), .B(n_857), .Y(n_1043) );
OR2x2_ASAP7_75t_L g1044 ( .A(n_991), .B(n_933), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_997), .B(n_971), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_981), .B(n_936), .Y(n_1046) );
INVxp67_ASAP7_75t_SL g1047 ( .A(n_1015), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g1048 ( .A1(n_1013), .A2(n_969), .B1(n_942), .B2(n_935), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_998), .B(n_965), .Y(n_1049) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_995), .B(n_969), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_998), .B(n_965), .Y(n_1051) );
INVxp67_ASAP7_75t_SL g1052 ( .A(n_1019), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_995), .B(n_1001), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_994), .B(n_936), .Y(n_1054) );
NAND2xp5_ASAP7_75t_L g1055 ( .A(n_996), .B(n_970), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1004), .Y(n_1056) );
INVx1_ASAP7_75t_SL g1057 ( .A(n_1022), .Y(n_1057) );
OR2x2_ASAP7_75t_L g1058 ( .A(n_1000), .B(n_939), .Y(n_1058) );
INVxp67_ASAP7_75t_L g1059 ( .A(n_1027), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1005), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1001), .B(n_969), .Y(n_1061) );
BUFx2_ASAP7_75t_SL g1062 ( .A(n_983), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_1007), .Y(n_1063) );
NOR2x1p5_ASAP7_75t_L g1064 ( .A(n_983), .B(n_942), .Y(n_1064) );
OR2x2_ASAP7_75t_L g1065 ( .A(n_1000), .B(n_939), .Y(n_1065) );
INVx1_ASAP7_75t_SL g1066 ( .A(n_1022), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1008), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1068 ( .A(n_987), .Y(n_1068) );
INVx1_ASAP7_75t_SL g1069 ( .A(n_976), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_1020), .A2(n_962), .B1(n_942), .B2(n_935), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_1009), .B(n_969), .Y(n_1071) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_1053), .B(n_1016), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_1047), .Y(n_1073) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1030), .Y(n_1074) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1053), .B(n_1016), .Y(n_1075) );
AND2x4_ASAP7_75t_L g1076 ( .A(n_1068), .B(n_988), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_1052), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_1038), .B(n_1009), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_1049), .B(n_1023), .Y(n_1079) );
XNOR2xp5_ASAP7_75t_L g1080 ( .A(n_1064), .B(n_980), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1061), .B(n_1023), .Y(n_1081) );
INVx1_ASAP7_75t_SL g1082 ( .A(n_1069), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_1049), .B(n_1024), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1063), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1063), .Y(n_1085) );
NAND2xp5_ASAP7_75t_L g1086 ( .A(n_1038), .B(n_1010), .Y(n_1086) );
AOI22xp33_ASAP7_75t_L g1087 ( .A1(n_1068), .A2(n_988), .B1(n_1002), .B2(n_987), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1067), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_1067), .Y(n_1089) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_1051), .B(n_1024), .Y(n_1090) );
INVxp67_ASAP7_75t_SL g1091 ( .A(n_1039), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1037), .Y(n_1092) );
INVx2_ASAP7_75t_L g1093 ( .A(n_1030), .Y(n_1093) );
INVx1_ASAP7_75t_SL g1094 ( .A(n_1062), .Y(n_1094) );
NOR2xp33_ASAP7_75t_L g1095 ( .A(n_1035), .B(n_980), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_1028), .B(n_1010), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_1051), .B(n_1026), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1028), .B(n_1026), .Y(n_1098) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1040), .Y(n_1099) );
INVx3_ASAP7_75t_SL g1100 ( .A(n_1057), .Y(n_1100) );
INVxp33_ASAP7_75t_L g1101 ( .A(n_1043), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1058), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1073), .Y(n_1103) );
INVx3_ASAP7_75t_L g1104 ( .A(n_1094), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1077), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_1079), .B(n_1058), .Y(n_1106) );
INVx2_ASAP7_75t_L g1107 ( .A(n_1079), .Y(n_1107) );
NAND2xp5_ASAP7_75t_L g1108 ( .A(n_1102), .B(n_1044), .Y(n_1108) );
OR2x2_ASAP7_75t_L g1109 ( .A(n_1083), .B(n_1065), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1084), .Y(n_1110) );
AOI21xp33_ASAP7_75t_L g1111 ( .A1(n_1101), .A2(n_1002), .B(n_1021), .Y(n_1111) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_1087), .A2(n_1048), .B1(n_1070), .B2(n_1066), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_1085), .Y(n_1113) );
OAI32xp33_ASAP7_75t_L g1114 ( .A1(n_1082), .A2(n_983), .A3(n_1044), .B1(n_1059), .B2(n_1065), .Y(n_1114) );
AOI322xp5_ASAP7_75t_L g1115 ( .A1(n_1091), .A2(n_1054), .A3(n_1029), .B1(n_1036), .B2(n_1042), .C1(n_1033), .C2(n_1050), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1102), .B(n_1029), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1088), .Y(n_1117) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1089), .Y(n_1118) );
NAND2xp5_ASAP7_75t_SL g1119 ( .A(n_1080), .B(n_1018), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1072), .B(n_1033), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1121 ( .A1(n_1101), .A2(n_988), .B1(n_1017), .B2(n_1006), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1092), .Y(n_1122) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_1099), .B(n_1012), .C(n_1046), .Y(n_1123) );
INVx1_ASAP7_75t_L g1124 ( .A(n_1108), .Y(n_1124) );
AOI22xp5_ASAP7_75t_L g1125 ( .A1(n_1112), .A2(n_1100), .B1(n_1076), .B2(n_1080), .Y(n_1125) );
OAI221xp5_ASAP7_75t_SL g1126 ( .A1(n_1115), .A2(n_975), .B1(n_1090), .B2(n_1097), .C(n_1083), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1108), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1103), .B(n_1072), .Y(n_1128) );
NAND2xp5_ASAP7_75t_L g1129 ( .A(n_1105), .B(n_1075), .Y(n_1129) );
AOI211xp5_ASAP7_75t_L g1130 ( .A1(n_1119), .A2(n_1100), .B(n_1095), .C(n_1018), .Y(n_1130) );
HB1xp67_ASAP7_75t_L g1131 ( .A(n_1104), .Y(n_1131) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_1114), .A2(n_1098), .B1(n_1096), .B2(n_1078), .C(n_1086), .Y(n_1132) );
INVxp67_ASAP7_75t_L g1133 ( .A(n_1104), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g1134 ( .A1(n_1111), .A2(n_1076), .B(n_1090), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1116), .Y(n_1135) );
AOI221xp5_ASAP7_75t_L g1136 ( .A1(n_1123), .A2(n_1111), .B1(n_1122), .B2(n_1116), .C(n_1107), .Y(n_1136) );
NOR3xp33_ASAP7_75t_L g1137 ( .A(n_1110), .B(n_956), .C(n_880), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g1138 ( .A1(n_1125), .A2(n_1076), .B1(n_1121), .B2(n_1118), .Y(n_1138) );
OAI221xp5_ASAP7_75t_SL g1139 ( .A1(n_1132), .A2(n_1109), .B1(n_1106), .B2(n_1097), .C(n_1120), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1131), .Y(n_1140) );
AOI222xp33_ASAP7_75t_L g1141 ( .A1(n_1136), .A2(n_1113), .B1(n_1117), .B2(n_1055), .C1(n_1075), .C2(n_1042), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1142 ( .A(n_1126), .B(n_934), .C(n_1056), .Y(n_1142) );
AOI221xp5_ASAP7_75t_SL g1143 ( .A1(n_1134), .A2(n_1133), .B1(n_1130), .B2(n_1124), .C(n_1127), .Y(n_1143) );
XNOR2x1_ASAP7_75t_L g1144 ( .A(n_1135), .B(n_1062), .Y(n_1144) );
OAI21xp33_ASAP7_75t_SL g1145 ( .A1(n_1133), .A2(n_1081), .B(n_1071), .Y(n_1145) );
AOI21xp33_ASAP7_75t_L g1146 ( .A1(n_1128), .A2(n_977), .B(n_880), .Y(n_1146) );
NAND2xp5_ASAP7_75t_SL g1147 ( .A(n_1143), .B(n_1137), .Y(n_1147) );
OAI221xp5_ASAP7_75t_SL g1148 ( .A1(n_1142), .A2(n_1129), .B1(n_1011), .B2(n_1034), .C(n_1045), .Y(n_1148) );
NOR3xp33_ASAP7_75t_L g1149 ( .A(n_1142), .B(n_909), .C(n_1025), .Y(n_1149) );
OAI221xp5_ASAP7_75t_L g1150 ( .A1(n_1139), .A2(n_1041), .B1(n_1060), .B2(n_1031), .C(n_1032), .Y(n_1150) );
NAND3xp33_ASAP7_75t_L g1151 ( .A(n_1141), .B(n_1093), .C(n_1074), .Y(n_1151) );
NOR3xp33_ASAP7_75t_L g1152 ( .A(n_1140), .B(n_892), .C(n_999), .Y(n_1152) );
NAND4xp25_ASAP7_75t_L g1153 ( .A(n_1138), .B(n_923), .C(n_847), .D(n_868), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1152), .B(n_1144), .Y(n_1154) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1151), .Y(n_1155) );
NAND3xp33_ASAP7_75t_L g1156 ( .A(n_1147), .B(n_1145), .C(n_1146), .Y(n_1156) );
NAND3xp33_ASAP7_75t_L g1157 ( .A(n_1148), .B(n_1093), .C(n_1074), .Y(n_1157) );
AND3x4_ASAP7_75t_L g1158 ( .A(n_1149), .B(n_923), .C(n_847), .Y(n_1158) );
NOR3xp33_ASAP7_75t_L g1159 ( .A(n_1156), .B(n_1153), .C(n_1150), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1155), .Y(n_1160) );
INVx3_ASAP7_75t_L g1161 ( .A(n_1154), .Y(n_1161) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1157), .Y(n_1162) );
INVxp67_ASAP7_75t_SL g1163 ( .A(n_1160), .Y(n_1163) );
OA22x2_ASAP7_75t_L g1164 ( .A1(n_1161), .A2(n_1158), .B1(n_976), .B2(n_1081), .Y(n_1164) );
XNOR2xp5_ASAP7_75t_L g1165 ( .A(n_1161), .B(n_847), .Y(n_1165) );
AOI22x1_ASAP7_75t_L g1166 ( .A1(n_1163), .A2(n_1162), .B1(n_1159), .B2(n_868), .Y(n_1166) );
BUFx8_ASAP7_75t_L g1167 ( .A(n_1165), .Y(n_1167) );
HB1xp67_ASAP7_75t_L g1168 ( .A(n_1164), .Y(n_1168) );
AOI222xp33_ASAP7_75t_L g1169 ( .A1(n_1168), .A2(n_1159), .B1(n_970), .B2(n_963), .C1(n_868), .C2(n_888), .Y(n_1169) );
OA21x2_ASAP7_75t_L g1170 ( .A1(n_1166), .A2(n_888), .B(n_1014), .Y(n_1170) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_1169), .A2(n_1167), .B1(n_963), .B2(n_888), .Y(n_1171) );
OAI21xp5_ASAP7_75t_L g1172 ( .A1(n_1170), .A2(n_963), .B(n_907), .Y(n_1172) );
OR2x6_ASAP7_75t_L g1173 ( .A(n_1172), .B(n_1171), .Y(n_1173) );
AOI21xp5_ASAP7_75t_L g1174 ( .A1(n_1173), .A2(n_963), .B(n_850), .Y(n_1174) );
endmodule