module fake_jpeg_31931_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_0),
.B(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_36),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_17),
.B(n_0),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_22),
.Y(n_61)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

BUFx2_ASAP7_75t_SL g54 ( 
.A(n_51),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_54),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_19),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_59),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_33),
.B1(n_34),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_24),
.B1(n_31),
.B2(n_3),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_71),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_25),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_73),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_76),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_24),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_45),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_22),
.B1(n_34),
.B2(n_24),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_28),
.B1(n_20),
.B2(n_27),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_45),
.A2(n_34),
.B1(n_21),
.B2(n_33),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_83),
.B1(n_33),
.B2(n_23),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_84),
.Y(n_103)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_82),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_21),
.B1(n_33),
.B2(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_38),
.B(n_29),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_87),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_46),
.B(n_29),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_88),
.Y(n_127)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_89),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_90),
.B(n_109),
.Y(n_134)
);

OR2x4_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_23),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_98),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_23),
.B(n_20),
.C(n_28),
.Y(n_92)
);

O2A1O1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_92),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_111),
.B1(n_66),
.B2(n_86),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_116),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_30),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_27),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_114),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_55),
.A2(n_16),
.B(n_14),
.C(n_3),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_67),
.B(n_7),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_14),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_70),
.A2(n_1),
.B(n_2),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_115),
.A2(n_6),
.B(n_8),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_83),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_86),
.C(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_117),
.B(n_130),
.Y(n_168)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_76),
.A3(n_62),
.B1(n_85),
.B2(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_132),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_99),
.B(n_2),
.C(n_4),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_120),
.A2(n_113),
.B(n_112),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_125),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_80),
.B1(n_58),
.B2(n_52),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_128),
.B1(n_131),
.B2(n_136),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_68),
.B1(n_69),
.B2(n_53),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_79),
.B1(n_78),
.B2(n_10),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_78),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_79),
.B1(n_8),
.B2(n_10),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_92),
.B(n_115),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_95),
.B(n_11),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_140),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_13),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_91),
.A2(n_106),
.B1(n_104),
.B2(n_102),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_100),
.B1(n_114),
.B2(n_108),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_96),
.C(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_97),
.Y(n_162)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_145),
.B(n_147),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_148),
.B(n_150),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_116),
.B1(n_92),
.B2(n_97),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_162),
.Y(n_173)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_109),
.B(n_88),
.Y(n_155)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_151),
.B1(n_146),
.B2(n_150),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_165),
.Y(n_181)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_103),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_169),
.B(n_131),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_158),
.B(n_121),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_145),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_123),
.B1(n_135),
.B2(n_128),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_164),
.B1(n_155),
.B2(n_147),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_129),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_182),
.C(n_159),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_SL g180 ( 
.A1(n_161),
.A2(n_130),
.A3(n_136),
.B1(n_141),
.B2(n_126),
.C1(n_135),
.C2(n_129),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_169),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_117),
.C(n_126),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_184),
.A2(n_177),
.B(n_170),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_125),
.B1(n_100),
.B2(n_88),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_188),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_105),
.B(n_101),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_187),
.A2(n_155),
.B(n_154),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_90),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_189),
.A2(n_191),
.B(n_200),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_190),
.B(n_193),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_178),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_203),
.C(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_198),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_199),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_170),
.A2(n_164),
.B1(n_155),
.B2(n_165),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_181),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_173),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_188),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_185),
.C(n_179),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_203),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_205),
.C(n_206),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_184),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_183),
.C(n_187),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_195),
.C(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_172),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_221),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_214),
.A2(n_189),
.B(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_211),
.A2(n_184),
.B(n_172),
.Y(n_219)
);

NOR2xp67_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_223),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_205),
.C(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_210),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_196),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_224),
.B1(n_208),
.B2(n_186),
.Y(n_225)
);

AOI321xp33_ASAP7_75t_L g223 ( 
.A1(n_204),
.A2(n_175),
.A3(n_155),
.B1(n_192),
.B2(n_197),
.C(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_215),
.B(n_153),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_230),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_176),
.C(n_148),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_209),
.C(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_229),
.B(n_176),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_213),
.B1(n_164),
.B2(n_198),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_228),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_176),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_235),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_231),
.C(n_227),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.C(n_156),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_233),
.A2(n_230),
.B1(n_231),
.B2(n_149),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_240),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_233),
.B(n_149),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_241),
.Y(n_245)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_239),
.A3(n_238),
.B1(n_156),
.B2(n_122),
.C1(n_101),
.C2(n_143),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_244),
.B(n_242),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_245),
.Y(n_247)
);


endmodule