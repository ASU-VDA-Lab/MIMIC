module fake_jpeg_20459_n_187 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_187);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_187;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_13),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_31),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_25),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_58),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_20),
.B1(n_15),
.B2(n_19),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_37),
.B1(n_35),
.B2(n_24),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_20),
.B1(n_15),
.B2(n_19),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_49),
.A2(n_24),
.B1(n_37),
.B2(n_17),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_53),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_52),
.Y(n_81)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_57),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_66),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_35),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_65),
.A2(n_89),
.B1(n_30),
.B2(n_4),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_29),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_69),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_16),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_79),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_39),
.B1(n_40),
.B2(n_33),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_72),
.A2(n_80),
.B1(n_87),
.B2(n_88),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_21),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_2),
.Y(n_103)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_17),
.B1(n_21),
.B2(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_28),
.B1(n_27),
.B2(n_18),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_48),
.Y(n_90)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_68),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_99),
.C(n_105),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_22),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_102),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_53),
.B(n_27),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_63),
.B(n_81),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_51),
.C(n_47),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_28),
.A3(n_47),
.B1(n_48),
.B2(n_38),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_2),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_65),
.B(n_61),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g130 ( 
.A(n_104),
.B(n_74),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_65),
.B(n_51),
.C(n_30),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_61),
.B1(n_4),
.B2(n_5),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_88),
.B1(n_76),
.B2(n_75),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_112),
.B(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_69),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_119),
.B1(n_93),
.B2(n_108),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_127),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_62),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_116),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_70),
.B1(n_83),
.B2(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

BUFx24_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_83),
.C(n_81),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_100),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_109),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_105),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_96),
.C(n_90),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_139),
.B(n_121),
.Y(n_154)
);

OAI211xp5_ASAP7_75t_SL g134 ( 
.A1(n_124),
.A2(n_111),
.B(n_110),
.C(n_104),
.Y(n_134)
);

AOI222xp33_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_130),
.B1(n_127),
.B2(n_125),
.C1(n_107),
.C2(n_86),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_119),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_102),
.B(n_100),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_122),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_115),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_95),
.B1(n_103),
.B2(n_78),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_123),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_146),
.B(n_151),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_139),
.B1(n_141),
.B2(n_131),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_154),
.B(n_155),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_118),
.C(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_152),
.C(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_142),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_130),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

OAI22x1_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_138),
.B1(n_134),
.B2(n_136),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_163),
.B1(n_135),
.B2(n_133),
.Y(n_167)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_164),
.B(n_4),
.Y(n_171)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_135),
.B(n_139),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_149),
.C(n_141),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_158),
.A2(n_156),
.B(n_125),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_160),
.B(n_6),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_107),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_161),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_82),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_177),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_159),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_176),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_175),
.A2(n_168),
.B1(n_160),
.B2(n_167),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_173),
.B1(n_170),
.B2(n_166),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_181),
.A2(n_182),
.B(n_180),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_178),
.A2(n_173),
.B1(n_169),
.B2(n_11),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_184),
.A3(n_9),
.B1(n_14),
.B2(n_12),
.C1(n_11),
.C2(n_74),
.Y(n_185)
);

NOR2x1_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_180),
.Y(n_184)
);

AOI322xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_176),
.C2(n_159),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_5),
.Y(n_187)
);


endmodule