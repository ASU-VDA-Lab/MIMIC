module fake_ariane_364_n_1326 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1326);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1326;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_868;
wire n_1314;
wire n_884;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_461;
wire n_1121;
wire n_490;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_746;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_776;
wire n_424;
wire n_466;
wire n_1263;
wire n_346;
wire n_552;
wire n_348;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1266;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_1204;
wire n_994;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1148;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_47),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_163),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_83),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_182),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_239),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_93),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_43),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_288),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_2),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_137),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_157),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_325),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_173),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_138),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_62),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_204),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_171),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_87),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_112),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_273),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_214),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_81),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_231),
.B(n_17),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_18),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_118),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_72),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_283),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_289),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_0),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_135),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_269),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_90),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_175),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_217),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_272),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_294),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_30),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_61),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_17),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_196),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_203),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_47),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_140),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_284),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_255),
.Y(n_373)
);

BUFx8_ASAP7_75t_SL g374 ( 
.A(n_89),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_232),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_311),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_81),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_293),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_183),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_267),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_36),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_35),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_304),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_265),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_66),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_67),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_261),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_56),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_111),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_155),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_122),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_99),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_314),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_238),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_117),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_268),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_199),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_190),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_148),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_274),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_30),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_215),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_71),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_9),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_139),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_14),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_67),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_131),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_65),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_109),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_201),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_212),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_64),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_233),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_6),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_143),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_98),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_278),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_129),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_316),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_20),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_295),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_280),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_236),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_193),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_174),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_150),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_263),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_169),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_237),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_252),
.B(n_251),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_210),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_240),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_149),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_68),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_260),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_55),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_38),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_189),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_205),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_89),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_85),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_26),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_202),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_277),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_264),
.Y(n_448)
);

BUFx10_ASAP7_75t_L g449 ( 
.A(n_27),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_51),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_123),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_213),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_317),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_282),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_59),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_164),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_106),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_188),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_74),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_93),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_275),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_78),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_124),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_168),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_243),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_245),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_103),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_70),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_14),
.Y(n_469)
);

BUFx10_ASAP7_75t_L g470 ( 
.A(n_55),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_18),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_286),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_114),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_221),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_326),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_285),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_105),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_144),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_145),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_186),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_107),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_312),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_197),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_309),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_303),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_41),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_64),
.Y(n_487)
);

INVx5_ASAP7_75t_L g488 ( 
.A(n_363),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_377),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_453),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_347),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_440),
.B(n_1),
.Y(n_493)
);

CKINVDCx11_ASAP7_75t_R g494 ( 
.A(n_449),
.Y(n_494)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_363),
.Y(n_495)
);

BUFx12f_ASAP7_75t_L g496 ( 
.A(n_442),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_469),
.Y(n_497)
);

AND2x4_ASAP7_75t_L g498 ( 
.A(n_361),
.B(n_1),
.Y(n_498)
);

INVx5_ASAP7_75t_L g499 ( 
.A(n_442),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_343),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_347),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_469),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_374),
.Y(n_503)
);

OAI22x1_ASAP7_75t_SL g504 ( 
.A1(n_367),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_347),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_343),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_361),
.B(n_3),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_388),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_485),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_469),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_347),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_485),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_370),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_469),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_456),
.B(n_4),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_456),
.B(n_5),
.Y(n_516)
);

AOI22x1_ASAP7_75t_SL g517 ( 
.A1(n_460),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_517)
);

BUFx8_ASAP7_75t_SL g518 ( 
.A(n_353),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_350),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_420),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_335),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_329),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_449),
.B(n_10),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_333),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_336),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_346),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_352),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_400),
.Y(n_528)
);

INVx5_ASAP7_75t_L g529 ( 
.A(n_400),
.Y(n_529)
);

BUFx8_ASAP7_75t_L g530 ( 
.A(n_384),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_468),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_349),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_354),
.Y(n_533)
);

CKINVDCx6p67_ASAP7_75t_R g534 ( 
.A(n_358),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_327),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_338),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_438),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_418),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_328),
.B(n_12),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_383),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_357),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_468),
.Y(n_542)
);

AND2x4_ASAP7_75t_L g543 ( 
.A(n_439),
.B(n_13),
.Y(n_543)
);

INVx6_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_381),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_462),
.B(n_15),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_418),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_360),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_366),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_368),
.B(n_16),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_386),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_368),
.B(n_19),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_382),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_392),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_383),
.B(n_19),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_402),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_387),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_411),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_418),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_401),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_425),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_489),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_491),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_495),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_561),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_518),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_537),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_534),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_522),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_495),
.B(n_428),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_494),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_503),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_549),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_492),
.Y(n_575)
);

NOR2xp67_ASAP7_75t_L g576 ( 
.A(n_488),
.B(n_412),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_496),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_512),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_535),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_536),
.Y(n_582)
);

AO21x2_ASAP7_75t_L g583 ( 
.A1(n_539),
.A2(n_351),
.B(n_337),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_557),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_L g585 ( 
.A(n_488),
.B(n_458),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_544),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_499),
.B(n_448),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_490),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_499),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_509),
.B(n_461),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_509),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_544),
.Y(n_592)
);

BUFx10_ASAP7_75t_L g593 ( 
.A(n_498),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_509),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_529),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_560),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_530),
.Y(n_597)
);

CKINVDCx16_ASAP7_75t_R g598 ( 
.A(n_550),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_530),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_548),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_553),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_492),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_500),
.B(n_463),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_525),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_531),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_526),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_542),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_506),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_521),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_532),
.Y(n_610)
);

NAND3xp33_ASAP7_75t_L g611 ( 
.A(n_565),
.B(n_516),
.C(n_507),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_570),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_571),
.B(n_498),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_582),
.Y(n_614)
);

BUFx8_ASAP7_75t_L g615 ( 
.A(n_601),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_562),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_588),
.B(n_523),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_563),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_587),
.B(n_552),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_590),
.B(n_555),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_593),
.B(n_515),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_603),
.B(n_508),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_583),
.B(n_540),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_580),
.B(n_543),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_583),
.B(n_543),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_564),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_609),
.B(n_546),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_584),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_596),
.B(n_546),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_579),
.B(n_606),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_564),
.B(n_598),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_604),
.B(n_497),
.Y(n_632)
);

OR2x6_ASAP7_75t_L g633 ( 
.A(n_608),
.B(n_493),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_610),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_566),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_575),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_589),
.B(n_591),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_586),
.B(n_504),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_605),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_581),
.B(n_520),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_607),
.B(n_519),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_594),
.B(n_529),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_568),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_602),
.Y(n_644)
);

AO221x1_ASAP7_75t_L g645 ( 
.A1(n_600),
.A2(n_504),
.B1(n_417),
.B2(n_459),
.C(n_455),
.Y(n_645)
);

AOI221xp5_ASAP7_75t_L g646 ( 
.A1(n_573),
.A2(n_471),
.B1(n_487),
.B2(n_467),
.C(n_437),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_595),
.Y(n_648)
);

INVxp33_ASAP7_75t_L g649 ( 
.A(n_576),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_585),
.B(n_502),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_586),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_597),
.B(n_385),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_592),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_599),
.Y(n_654)
);

AOI221xp5_ASAP7_75t_L g655 ( 
.A1(n_574),
.A2(n_533),
.B1(n_541),
.B2(n_527),
.C(n_526),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_577),
.B(n_578),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_592),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_569),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_567),
.B(n_510),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_595),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_603),
.B(n_519),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_571),
.B(n_527),
.Y(n_663)
);

BUFx6f_ASAP7_75t_SL g664 ( 
.A(n_564),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_587),
.B(n_538),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_571),
.B(n_533),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_603),
.B(n_541),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_562),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_621),
.A2(n_620),
.B(n_630),
.Y(n_670)
);

BUFx12f_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_628),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_663),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_667),
.B(n_332),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_616),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_628),
.B(n_545),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_651),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_618),
.Y(n_678)
);

CKINVDCx11_ASAP7_75t_R g679 ( 
.A(n_660),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_611),
.A2(n_405),
.B1(n_409),
.B2(n_408),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_619),
.B(n_376),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_614),
.B(n_551),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_617),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_639),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_611),
.A2(n_344),
.B1(n_359),
.B2(n_356),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_632),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_632),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_612),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_668),
.B(n_430),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_L g690 ( 
.A(n_631),
.B(n_551),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_624),
.B(n_554),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_629),
.B(n_625),
.Y(n_692)
);

HB1xp67_ASAP7_75t_L g693 ( 
.A(n_657),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_626),
.B(n_415),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_622),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_653),
.Y(n_696)
);

INVx5_ASAP7_75t_L g697 ( 
.A(n_624),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_634),
.B(n_419),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_640),
.A2(n_365),
.B1(n_444),
.B2(n_406),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_665),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_643),
.B(n_423),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_662),
.B(n_556),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_615),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_624),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_630),
.B(n_556),
.Y(n_705)
);

AND2x4_ASAP7_75t_SL g706 ( 
.A(n_633),
.B(n_558),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_633),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_627),
.B(n_558),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_647),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_660),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_664),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_623),
.B(n_443),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_655),
.B(n_445),
.Y(n_713)
);

NOR2x2_ASAP7_75t_L g714 ( 
.A(n_638),
.B(n_517),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_646),
.A2(n_450),
.B1(n_401),
.B2(n_334),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_669),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_637),
.A2(n_372),
.B1(n_373),
.B2(n_371),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_648),
.B(n_661),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_635),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_659),
.B(n_654),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_664),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_652),
.B(n_477),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_660),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_658),
.B(n_486),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_666),
.B(n_330),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_649),
.B(n_331),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_636),
.Y(n_727)
);

INVxp67_ASAP7_75t_L g728 ( 
.A(n_656),
.Y(n_728)
);

INVxp33_ASAP7_75t_L g729 ( 
.A(n_650),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_644),
.A2(n_399),
.B(n_403),
.C(n_375),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_642),
.A2(n_413),
.B1(n_416),
.B2(n_404),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_638),
.B(n_433),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_638),
.B(n_421),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_645),
.A2(n_432),
.B1(n_434),
.B2(n_431),
.Y(n_734)
);

INVx8_ASAP7_75t_L g735 ( 
.A(n_664),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_632),
.Y(n_736)
);

BUFx12f_ASAP7_75t_L g737 ( 
.A(n_615),
.Y(n_737)
);

AO21x2_ASAP7_75t_L g738 ( 
.A1(n_623),
.A2(n_447),
.B(n_436),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_641),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_641),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_632),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_663),
.B(n_339),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_641),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_632),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_632),
.Y(n_745)
);

CKINVDCx6p67_ASAP7_75t_R g746 ( 
.A(n_664),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_647),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_632),
.Y(n_748)
);

BUFx6f_ASAP7_75t_L g749 ( 
.A(n_647),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_613),
.B(n_473),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_641),
.B(n_514),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_663),
.B(n_340),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_614),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_611),
.A2(n_475),
.B1(n_476),
.B2(n_474),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_632),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_632),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_611),
.A2(n_484),
.B1(n_481),
.B2(n_410),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_639),
.B(n_20),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_616),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_615),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_663),
.B(n_341),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_663),
.B(n_342),
.Y(n_762)
);

NAND3xp33_ASAP7_75t_SL g763 ( 
.A(n_674),
.B(n_348),
.C(n_345),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_697),
.B(n_753),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_719),
.Y(n_765)
);

BUFx8_ASAP7_75t_L g766 ( 
.A(n_671),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_670),
.A2(n_362),
.B(n_355),
.Y(n_767)
);

INVxp33_ASAP7_75t_L g768 ( 
.A(n_682),
.Y(n_768)
);

O2A1O1Ixp5_ASAP7_75t_L g769 ( 
.A1(n_750),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_R g770 ( 
.A(n_677),
.B(n_364),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_697),
.B(n_22),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_692),
.B(n_369),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_716),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_684),
.Y(n_774)
);

INVxp33_ASAP7_75t_L g775 ( 
.A(n_682),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_742),
.B(n_378),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_752),
.B(n_379),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_761),
.B(n_380),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_740),
.B(n_695),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_678),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_685),
.A2(n_390),
.B(n_391),
.C(n_389),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_705),
.A2(n_394),
.B(n_393),
.Y(n_782)
);

CKINVDCx11_ASAP7_75t_R g783 ( 
.A(n_737),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_729),
.B(n_683),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_746),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_743),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_762),
.A2(n_396),
.B(n_397),
.C(n_395),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_672),
.B(n_398),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_700),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_706),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_691),
.B(n_689),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_707),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_680),
.A2(n_754),
.B(n_708),
.C(n_713),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_725),
.A2(n_414),
.B(n_407),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_747),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_691),
.Y(n_796)
);

AO21x2_ASAP7_75t_L g797 ( 
.A1(n_738),
.A2(n_480),
.B(n_425),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_760),
.Y(n_798)
);

AO21x1_ASAP7_75t_L g799 ( 
.A1(n_757),
.A2(n_712),
.B(n_681),
.Y(n_799)
);

OAI22x1_ASAP7_75t_L g800 ( 
.A1(n_733),
.A2(n_424),
.B1(n_426),
.B2(n_422),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_686),
.A2(n_429),
.B(n_427),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_687),
.A2(n_441),
.B(n_435),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_735),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_736),
.B(n_446),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_741),
.B(n_744),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_679),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_745),
.A2(n_452),
.B(n_451),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_748),
.A2(n_457),
.B(n_454),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_672),
.A2(n_465),
.B1(n_466),
.B2(n_464),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_755),
.A2(n_478),
.B(n_472),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_697),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_756),
.B(n_479),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_759),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_698),
.A2(n_482),
.B(n_483),
.C(n_480),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_720),
.A2(n_483),
.B1(n_505),
.B2(n_501),
.Y(n_815)
);

BUFx4f_ASAP7_75t_L g816 ( 
.A(n_735),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_672),
.B(n_710),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_718),
.A2(n_483),
.B(n_501),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_676),
.B(n_24),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_676),
.B(n_25),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_747),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_739),
.B(n_501),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_751),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_717),
.B(n_26),
.C(n_28),
.Y(n_824)
);

BUFx2_ASAP7_75t_L g825 ( 
.A(n_693),
.Y(n_825)
);

NOR2xp67_ASAP7_75t_L g826 ( 
.A(n_711),
.B(n_721),
.Y(n_826)
);

AND2x6_ASAP7_75t_L g827 ( 
.A(n_747),
.B(n_505),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_702),
.B(n_28),
.Y(n_828)
);

BUFx12f_ASAP7_75t_L g829 ( 
.A(n_703),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_749),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_704),
.B(n_511),
.Y(n_831)
);

OAI22x1_ASAP7_75t_L g832 ( 
.A1(n_734),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_749),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_728),
.B(n_29),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_694),
.A2(n_547),
.B(n_528),
.Y(n_835)
);

O2A1O1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_758),
.A2(n_34),
.B(n_31),
.C(n_33),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_696),
.B(n_722),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_715),
.A2(n_561),
.B1(n_547),
.B2(n_559),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_749),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_727),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_722),
.A2(n_547),
.B1(n_559),
.B2(n_528),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_724),
.B(n_33),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_726),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_730),
.A2(n_41),
.B(n_39),
.C(n_40),
.Y(n_844)
);

AND2x6_ASAP7_75t_SL g845 ( 
.A(n_732),
.B(n_40),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_723),
.B(n_42),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_709),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_690),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_724),
.B(n_44),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_699),
.B(n_731),
.Y(n_850)
);

XOR2xp5_ASAP7_75t_L g851 ( 
.A(n_714),
.B(n_108),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_673),
.A2(n_48),
.B1(n_45),
.B2(n_46),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_688),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_673),
.B(n_46),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_673),
.B(n_48),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_753),
.Y(n_856)
);

NOR3xp33_ASAP7_75t_SL g857 ( 
.A(n_701),
.B(n_49),
.C(n_50),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_672),
.B(n_49),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_672),
.B(n_50),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_688),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_670),
.A2(n_113),
.B(n_110),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_673),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_753),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_673),
.B(n_52),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_670),
.A2(n_116),
.B(n_115),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_695),
.B(n_53),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_691),
.B(n_119),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_688),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_673),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_673),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_697),
.B(n_63),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_673),
.B(n_63),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_688),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_675),
.Y(n_874)
);

BUFx6f_ASAP7_75t_L g875 ( 
.A(n_747),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_753),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_673),
.A2(n_68),
.B1(n_65),
.B2(n_66),
.Y(n_877)
);

NAND3xp33_ASAP7_75t_L g878 ( 
.A(n_673),
.B(n_69),
.C(n_70),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_670),
.A2(n_121),
.B(n_120),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_677),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_672),
.B(n_69),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_672),
.B(n_71),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_673),
.B(n_73),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_688),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_695),
.B(n_75),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_750),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_886)
);

BUFx12f_ASAP7_75t_L g887 ( 
.A(n_679),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_750),
.A2(n_82),
.B(n_79),
.C(n_80),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_750),
.A2(n_84),
.B(n_80),
.C(n_83),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_753),
.Y(n_890)
);

NOR2xp67_ASAP7_75t_SL g891 ( 
.A(n_672),
.B(n_84),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_750),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_783),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_796),
.Y(n_894)
);

BUFx3_ASAP7_75t_L g895 ( 
.A(n_856),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_825),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_768),
.B(n_88),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_816),
.Y(n_898)
);

AO21x2_ASAP7_75t_L g899 ( 
.A1(n_797),
.A2(n_126),
.B(n_125),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_775),
.B(n_90),
.Y(n_900)
);

BUFx3_ASAP7_75t_L g901 ( 
.A(n_890),
.Y(n_901)
);

AO21x2_ASAP7_75t_L g902 ( 
.A1(n_799),
.A2(n_128),
.B(n_127),
.Y(n_902)
);

CKINVDCx6p67_ASAP7_75t_R g903 ( 
.A(n_887),
.Y(n_903)
);

BUFx2_ASAP7_75t_L g904 ( 
.A(n_774),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_803),
.Y(n_905)
);

INVx4_ASAP7_75t_L g906 ( 
.A(n_764),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_764),
.B(n_91),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_853),
.Y(n_908)
);

NAND2x1p5_ASAP7_75t_L g909 ( 
.A(n_863),
.B(n_130),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_805),
.A2(n_91),
.B(n_92),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_765),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_779),
.B(n_92),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_880),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_829),
.B(n_94),
.Y(n_914)
);

AOI22x1_ASAP7_75t_L g915 ( 
.A1(n_861),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_792),
.Y(n_916)
);

AND2x4_ASAP7_75t_L g917 ( 
.A(n_791),
.B(n_95),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_96),
.Y(n_918)
);

AOI22x1_ASAP7_75t_L g919 ( 
.A1(n_865),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_919)
);

BUFx2_ASAP7_75t_SL g920 ( 
.A(n_867),
.Y(n_920)
);

BUFx12f_ASAP7_75t_L g921 ( 
.A(n_766),
.Y(n_921)
);

OA21x2_ASAP7_75t_L g922 ( 
.A1(n_818),
.A2(n_133),
.B(n_132),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_860),
.Y(n_923)
);

NAND2x1p5_ASAP7_75t_L g924 ( 
.A(n_790),
.B(n_134),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_806),
.B(n_136),
.Y(n_925)
);

INVx2_ASAP7_75t_SL g926 ( 
.A(n_785),
.Y(n_926)
);

INVx5_ASAP7_75t_L g927 ( 
.A(n_867),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_811),
.B(n_97),
.Y(n_928)
);

BUFx2_ASAP7_75t_SL g929 ( 
.A(n_867),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_868),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_873),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_770),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_772),
.B(n_823),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_837),
.A2(n_102),
.B1(n_100),
.B2(n_101),
.Y(n_934)
);

INVx5_ASAP7_75t_L g935 ( 
.A(n_867),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_884),
.Y(n_936)
);

BUFx2_ASAP7_75t_SL g937 ( 
.A(n_826),
.Y(n_937)
);

CKINVDCx11_ASAP7_75t_R g938 ( 
.A(n_845),
.Y(n_938)
);

AOI22x1_ASAP7_75t_L g939 ( 
.A1(n_879),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_795),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_793),
.A2(n_104),
.B(n_105),
.Y(n_941)
);

BUFx2_ASAP7_75t_SL g942 ( 
.A(n_771),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_795),
.Y(n_943)
);

BUFx4f_ASAP7_75t_SL g944 ( 
.A(n_766),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_830),
.B(n_141),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_828),
.A2(n_104),
.B(n_142),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_814),
.A2(n_146),
.B(n_147),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_798),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_784),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_817),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_840),
.Y(n_951)
);

AO21x2_ASAP7_75t_L g952 ( 
.A1(n_767),
.A2(n_151),
.B(n_152),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_833),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_833),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_871),
.B(n_153),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_835),
.A2(n_154),
.B(n_156),
.Y(n_956)
);

AO21x2_ASAP7_75t_L g957 ( 
.A1(n_776),
.A2(n_158),
.B(n_159),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_833),
.Y(n_958)
);

AO21x2_ASAP7_75t_L g959 ( 
.A1(n_777),
.A2(n_160),
.B(n_161),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_876),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_773),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_875),
.Y(n_962)
);

OR2x6_ASAP7_75t_L g963 ( 
.A(n_849),
.B(n_162),
.Y(n_963)
);

AO21x2_ASAP7_75t_L g964 ( 
.A1(n_778),
.A2(n_165),
.B(n_166),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_786),
.B(n_167),
.Y(n_965)
);

BUFx2_ASAP7_75t_SL g966 ( 
.A(n_827),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_813),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_780),
.Y(n_968)
);

AO21x2_ASAP7_75t_L g969 ( 
.A1(n_787),
.A2(n_170),
.B(n_172),
.Y(n_969)
);

INVx5_ASAP7_75t_L g970 ( 
.A(n_827),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_875),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_789),
.Y(n_972)
);

BUFx3_ASAP7_75t_L g973 ( 
.A(n_875),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_821),
.Y(n_974)
);

AOI21x1_ASAP7_75t_L g975 ( 
.A1(n_822),
.A2(n_176),
.B(n_177),
.Y(n_975)
);

INVx8_ASAP7_75t_L g976 ( 
.A(n_827),
.Y(n_976)
);

BUFx3_ASAP7_75t_L g977 ( 
.A(n_839),
.Y(n_977)
);

BUFx4f_ASAP7_75t_SL g978 ( 
.A(n_866),
.Y(n_978)
);

OR2x6_ASAP7_75t_L g979 ( 
.A(n_819),
.B(n_178),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_820),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_885),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_854),
.A2(n_179),
.B(n_180),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_842),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_821),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_831),
.A2(n_181),
.B(n_184),
.Y(n_985)
);

AO21x2_ASAP7_75t_L g986 ( 
.A1(n_782),
.A2(n_185),
.B(n_187),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_874),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_848),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_850),
.A2(n_824),
.B1(n_832),
.B2(n_855),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_847),
.Y(n_990)
);

BUFx12f_ASAP7_75t_L g991 ( 
.A(n_848),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_769),
.Y(n_992)
);

BUFx2_ASAP7_75t_SL g993 ( 
.A(n_858),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_834),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_846),
.Y(n_995)
);

NAND2x1p5_ASAP7_75t_L g996 ( 
.A(n_788),
.B(n_191),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_859),
.B(n_192),
.Y(n_997)
);

BUFx2_ASAP7_75t_R g998 ( 
.A(n_881),
.Y(n_998)
);

OA21x2_ASAP7_75t_L g999 ( 
.A1(n_815),
.A2(n_194),
.B(n_195),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_864),
.A2(n_198),
.B(n_200),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_872),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_882),
.B(n_206),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_851),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_891),
.Y(n_1004)
);

AO21x2_ASAP7_75t_L g1005 ( 
.A1(n_763),
.A2(n_207),
.B(n_208),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_883),
.A2(n_209),
.B(n_211),
.Y(n_1006)
);

AO21x2_ASAP7_75t_L g1007 ( 
.A1(n_794),
.A2(n_216),
.B(n_218),
.Y(n_1007)
);

AOI22x1_ASAP7_75t_L g1008 ( 
.A1(n_801),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_857),
.Y(n_1009)
);

BUFx2_ASAP7_75t_R g1010 ( 
.A(n_804),
.Y(n_1010)
);

OA21x2_ASAP7_75t_L g1011 ( 
.A1(n_812),
.A2(n_223),
.B(n_224),
.Y(n_1011)
);

AOI22x1_ASAP7_75t_L g1012 ( 
.A1(n_802),
.A2(n_810),
.B1(n_807),
.B2(n_808),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_843),
.A2(n_225),
.B(n_226),
.Y(n_1013)
);

BUFx3_ASAP7_75t_L g1014 ( 
.A(n_800),
.Y(n_1014)
);

BUFx2_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_844),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_878),
.Y(n_1017)
);

BUFx12f_ASAP7_75t_L g1018 ( 
.A(n_852),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_841),
.B(n_227),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_888),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_SL g1021 ( 
.A(n_862),
.Y(n_1021)
);

OA21x2_ASAP7_75t_L g1022 ( 
.A1(n_992),
.A2(n_892),
.B(n_889),
.Y(n_1022)
);

OA21x2_ASAP7_75t_L g1023 ( 
.A1(n_992),
.A2(n_781),
.B(n_877),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_944),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_972),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_1021),
.A2(n_989),
.B1(n_1018),
.B2(n_912),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_908),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_923),
.Y(n_1028)
);

AO21x2_ASAP7_75t_L g1029 ( 
.A1(n_941),
.A2(n_836),
.B(n_870),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_976),
.Y(n_1030)
);

CKINVDCx11_ASAP7_75t_R g1031 ( 
.A(n_921),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_894),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1015),
.A2(n_869),
.B1(n_838),
.B2(n_809),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_893),
.Y(n_1034)
);

BUFx2_ASAP7_75t_R g1035 ( 
.A(n_949),
.Y(n_1035)
);

HB1xp67_ASAP7_75t_L g1036 ( 
.A(n_896),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_980),
.B(n_324),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_917),
.B(n_228),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_1020),
.A2(n_229),
.B1(n_230),
.B2(n_234),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_931),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_911),
.B(n_235),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_936),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_SL g1043 ( 
.A(n_910),
.B(n_241),
.C(n_242),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_976),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_895),
.Y(n_1045)
);

CKINVDCx11_ASAP7_75t_R g1046 ( 
.A(n_903),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_SL g1047 ( 
.A1(n_1014),
.A2(n_244),
.B1(n_246),
.B2(n_247),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_978),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_1048)
);

AOI22xp33_ASAP7_75t_L g1049 ( 
.A1(n_1019),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_898),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_904),
.Y(n_1051)
);

CKINVDCx8_ASAP7_75t_R g1052 ( 
.A(n_932),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_SL g1053 ( 
.A1(n_918),
.A2(n_1020),
.B1(n_1003),
.B2(n_1009),
.Y(n_1053)
);

OAI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_918),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_901),
.Y(n_1055)
);

NAND2x1p5_ASAP7_75t_L g1056 ( 
.A(n_970),
.B(n_262),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_981),
.A2(n_994),
.B1(n_968),
.B2(n_987),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_933),
.A2(n_270),
.B1(n_271),
.B2(n_276),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_930),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_917),
.B(n_279),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_951),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_960),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_SL g1063 ( 
.A(n_898),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_916),
.B(n_281),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_942),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_951),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_906),
.B(n_287),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_967),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_961),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_905),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_990),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_988),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_988),
.Y(n_1073)
);

CKINVDCx11_ASAP7_75t_R g1074 ( 
.A(n_938),
.Y(n_1074)
);

BUFx4f_ASAP7_75t_SL g1075 ( 
.A(n_991),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_920),
.A2(n_291),
.B1(n_292),
.B2(n_296),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_SL g1077 ( 
.A1(n_920),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_906),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_988),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_948),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_995),
.A2(n_300),
.B1(n_301),
.B2(n_302),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_942),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_950),
.B(n_323),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_955),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_955),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_963),
.Y(n_1086)
);

BUFx4f_ASAP7_75t_SL g1087 ( 
.A(n_926),
.Y(n_1087)
);

INVxp67_ASAP7_75t_SL g1088 ( 
.A(n_1016),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_913),
.B(n_305),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_977),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_963),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_946),
.B(n_306),
.C(n_307),
.Y(n_1092)
);

CKINVDCx11_ASAP7_75t_R g1093 ( 
.A(n_914),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_907),
.B(n_322),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_973),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_927),
.B(n_310),
.Y(n_1096)
);

OAI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_979),
.A2(n_914),
.B1(n_1016),
.B2(n_1001),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_928),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_897),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_900),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_927),
.B(n_321),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_979),
.B(n_315),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_1010),
.B(n_320),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_971),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_971),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_965),
.B(n_318),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_940),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_983),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_993),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_935),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_1036),
.Y(n_1111)
);

NAND2xp33_ASAP7_75t_SL g1112 ( 
.A(n_1062),
.B(n_1017),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_1024),
.B(n_983),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1051),
.B(n_998),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1045),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_1036),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_1065),
.B(n_935),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1031),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_SL g1119 ( 
.A(n_1026),
.B(n_934),
.C(n_925),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_1052),
.Y(n_1120)
);

CKINVDCx9p33_ASAP7_75t_R g1121 ( 
.A(n_1078),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1106),
.A2(n_1000),
.B(n_982),
.C(n_1006),
.Y(n_1122)
);

NOR3xp33_ASAP7_75t_SL g1123 ( 
.A(n_1034),
.B(n_937),
.C(n_1017),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1032),
.B(n_958),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1032),
.B(n_953),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_R g1126 ( 
.A(n_1070),
.B(n_958),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1029),
.A2(n_929),
.B1(n_915),
.B2(n_919),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1075),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1053),
.B(n_943),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_R g1130 ( 
.A(n_1063),
.B(n_984),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1068),
.Y(n_1131)
);

INVxp67_ASAP7_75t_L g1132 ( 
.A(n_1090),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_1046),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1050),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_1088),
.A2(n_1004),
.B1(n_919),
.B2(n_915),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1099),
.B(n_1100),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1027),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_R g1138 ( 
.A(n_1087),
.B(n_974),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_R g1139 ( 
.A(n_1093),
.B(n_974),
.Y(n_1139)
);

XNOR2xp5_ASAP7_75t_L g1140 ( 
.A(n_1108),
.B(n_1103),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1028),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_1080),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_1050),
.B(n_984),
.Y(n_1143)
);

AO32x2_ASAP7_75t_L g1144 ( 
.A1(n_1033),
.A2(n_954),
.A3(n_962),
.B1(n_939),
.B2(n_902),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_R g1145 ( 
.A(n_1074),
.B(n_1004),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1055),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1029),
.A2(n_939),
.B1(n_1012),
.B2(n_924),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1033),
.A2(n_1013),
.B(n_1002),
.Y(n_1148)
);

NAND2xp33_ASAP7_75t_R g1149 ( 
.A(n_1096),
.B(n_1011),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1094),
.B(n_954),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1054),
.A2(n_1004),
.B(n_1012),
.C(n_909),
.Y(n_1151)
);

NOR3xp33_ASAP7_75t_SL g1152 ( 
.A(n_1097),
.B(n_1091),
.C(n_1086),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_R g1153 ( 
.A(n_1096),
.B(n_999),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1098),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1109),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1030),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_1067),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1040),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_1049),
.A2(n_997),
.B1(n_996),
.B2(n_1008),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1037),
.B(n_1038),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1042),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_1035),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1071),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_SL g1164 ( 
.A(n_1084),
.B(n_969),
.C(n_1005),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1025),
.A2(n_899),
.A3(n_957),
.B(n_959),
.Y(n_1165)
);

NAND3xp33_ASAP7_75t_SL g1166 ( 
.A(n_1109),
.B(n_945),
.C(n_964),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1035),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_SL g1168 ( 
.A(n_1085),
.B(n_1007),
.C(n_986),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1060),
.B(n_966),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1095),
.B(n_966),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1104),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1066),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_1043),
.B(n_952),
.C(n_947),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_1064),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1072),
.Y(n_1175)
);

CKINVDCx16_ASAP7_75t_R g1176 ( 
.A(n_1102),
.Y(n_1176)
);

OAI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1058),
.A2(n_975),
.B1(n_922),
.B2(n_956),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1059),
.Y(n_1178)
);

NAND2xp33_ASAP7_75t_R g1179 ( 
.A(n_1101),
.B(n_922),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1073),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1079),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1061),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1069),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1044),
.B(n_985),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1092),
.A2(n_1043),
.B(n_1066),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1163),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1116),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1119),
.A2(n_1047),
.B1(n_1092),
.B2(n_1057),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1178),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_1172),
.B(n_1022),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1182),
.B(n_1023),
.Y(n_1191)
);

INVxp67_ASAP7_75t_L g1192 ( 
.A(n_1136),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1183),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1134),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1134),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1111),
.B(n_1022),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1137),
.B(n_1107),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1141),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1124),
.B(n_1082),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1134),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1158),
.B(n_1041),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1161),
.Y(n_1202)
);

OR2x2_ASAP7_75t_L g1203 ( 
.A(n_1155),
.B(n_1089),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1125),
.B(n_1105),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1184),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1131),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_1113),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1144),
.B(n_1076),
.Y(n_1208)
);

BUFx2_ASAP7_75t_L g1209 ( 
.A(n_1121),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1144),
.B(n_1077),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1154),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1176),
.A2(n_1076),
.B1(n_1077),
.B2(n_1048),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1144),
.B(n_1058),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1160),
.B(n_1039),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1129),
.B(n_1039),
.Y(n_1215)
);

OR2x6_ASAP7_75t_L g1216 ( 
.A(n_1157),
.B(n_1056),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1174),
.B(n_1110),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1152),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1169),
.B(n_1081),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_1149),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1170),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1186),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1186),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1187),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1192),
.B(n_1142),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1201),
.B(n_1171),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1198),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1212),
.A2(n_1122),
.B1(n_1127),
.B2(n_1147),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1198),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1205),
.B(n_1148),
.Y(n_1230)
);

NAND3xp33_ASAP7_75t_L g1231 ( 
.A(n_1188),
.B(n_1168),
.C(n_1185),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1211),
.B(n_1166),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_1207),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1217),
.B(n_1132),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1205),
.B(n_1164),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1217),
.B(n_1146),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1211),
.B(n_1115),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1190),
.B(n_1114),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1196),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1220),
.B(n_1117),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1208),
.B(n_1150),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1208),
.B(n_1135),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1210),
.B(n_1173),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1210),
.B(n_1165),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1209),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1189),
.B(n_1126),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1213),
.B(n_1191),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1240),
.B(n_1193),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1222),
.Y(n_1249)
);

NOR4xp25_ASAP7_75t_SL g1250 ( 
.A(n_1233),
.B(n_1209),
.C(n_1179),
.D(n_1153),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1239),
.B(n_1196),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1247),
.B(n_1190),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1223),
.Y(n_1253)
);

NOR2x1_ASAP7_75t_L g1254 ( 
.A(n_1237),
.B(n_1216),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1224),
.B(n_1204),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1245),
.B(n_1214),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1240),
.B(n_1193),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1241),
.B(n_1202),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1227),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1247),
.B(n_1199),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1238),
.B(n_1221),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1233),
.B(n_1207),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1243),
.B(n_1219),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1243),
.B(n_1191),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1229),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1242),
.B(n_1197),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_1237),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1238),
.B(n_1219),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1249),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1251),
.B(n_1232),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1263),
.B(n_1230),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1268),
.B(n_1230),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1253),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1251),
.B(n_1232),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_1248),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1259),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1264),
.A2(n_1228),
.B1(n_1231),
.B2(n_1213),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1265),
.Y(n_1278)
);

AOI32xp33_ASAP7_75t_L g1279 ( 
.A1(n_1264),
.A2(n_1242),
.A3(n_1215),
.B1(n_1218),
.B2(n_1244),
.Y(n_1279)
);

O2A1O1Ixp5_ASAP7_75t_L g1280 ( 
.A1(n_1255),
.A2(n_1246),
.B(n_1235),
.C(n_1226),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1252),
.B(n_1234),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1254),
.B(n_1235),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1261),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1257),
.A2(n_1215),
.B1(n_1244),
.B2(n_1112),
.Y(n_1284)
);

OAI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1277),
.A2(n_1266),
.B1(n_1258),
.B2(n_1260),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1279),
.A2(n_1262),
.B(n_1118),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1269),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1283),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1275),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1271),
.Y(n_1290)
);

AO22x2_ASAP7_75t_L g1291 ( 
.A1(n_1270),
.A2(n_1225),
.B1(n_1267),
.B2(n_1206),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1284),
.A2(n_1267),
.B1(n_1250),
.B2(n_1256),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1286),
.A2(n_1270),
.B1(n_1274),
.B2(n_1281),
.Y(n_1293)
);

O2A1O1Ixp33_ASAP7_75t_L g1294 ( 
.A1(n_1285),
.A2(n_1280),
.B(n_1274),
.C(n_1151),
.Y(n_1294)
);

NAND2x1_ASAP7_75t_L g1295 ( 
.A(n_1290),
.B(n_1272),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1287),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1288),
.B(n_1133),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_SL g1298 ( 
.A(n_1294),
.B(n_1292),
.C(n_1282),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1296),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1295),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1293),
.B(n_1273),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1297),
.Y(n_1302)
);

NOR4xp75_ASAP7_75t_L g1303 ( 
.A(n_1293),
.B(n_1290),
.C(n_1236),
.D(n_1120),
.Y(n_1303)
);

BUFx4_ASAP7_75t_R g1304 ( 
.A(n_1299),
.Y(n_1304)
);

NOR3xp33_ASAP7_75t_L g1305 ( 
.A(n_1298),
.B(n_1162),
.C(n_1167),
.Y(n_1305)
);

NOR3xp33_ASAP7_75t_SL g1306 ( 
.A(n_1301),
.B(n_1140),
.C(n_1145),
.Y(n_1306)
);

OAI211xp5_ASAP7_75t_L g1307 ( 
.A1(n_1305),
.A2(n_1301),
.B(n_1300),
.C(n_1302),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1306),
.B(n_1291),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1307),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1309),
.B(n_1308),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_SL g1311 ( 
.A1(n_1310),
.A2(n_1128),
.B1(n_1304),
.B2(n_1303),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1310),
.Y(n_1312)
);

AO22x2_ASAP7_75t_L g1313 ( 
.A1(n_1312),
.A2(n_1289),
.B1(n_1278),
.B2(n_1276),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1311),
.Y(n_1314)
);

OAI31xp33_ASAP7_75t_L g1315 ( 
.A1(n_1314),
.A2(n_1291),
.A3(n_1159),
.B(n_1177),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1313),
.B(n_1194),
.Y(n_1316)
);

NOR2x1_ASAP7_75t_L g1317 ( 
.A(n_1316),
.B(n_1083),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1315),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1318),
.A2(n_1282),
.B1(n_1123),
.B2(n_1181),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1317),
.A2(n_1195),
.B1(n_1200),
.B2(n_1194),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1319),
.B(n_1139),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1320),
.B(n_1138),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1321),
.A2(n_1175),
.B1(n_1180),
.B2(n_1156),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1322),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1324),
.B(n_1203),
.Y(n_1325)
);

AOI211xp5_ASAP7_75t_L g1326 ( 
.A1(n_1325),
.A2(n_1323),
.B(n_1143),
.C(n_1130),
.Y(n_1326)
);


endmodule