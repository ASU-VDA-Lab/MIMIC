module fake_jpeg_20718_n_108 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_108);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_108;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_106;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_28),
.Y(n_31)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_33),
.Y(n_42)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_23),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_31),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_31),
.B(n_29),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_18),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_50),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_26),
.B1(n_29),
.B2(n_24),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_48),
.A2(n_24),
.B1(n_25),
.B2(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_14),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_65),
.Y(n_68)
);

BUFx24_ASAP7_75t_SL g56 ( 
.A(n_49),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_56),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_31),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_17),
.C(n_22),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_46),
.B1(n_38),
.B2(n_18),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_49),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_61),
.B(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_70),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_39),
.B(n_50),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_76),
.Y(n_78)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_75),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_82),
.B1(n_84),
.B2(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_58),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_21),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_83),
.A2(n_20),
.B(n_17),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_54),
.B1(n_40),
.B2(n_21),
.Y(n_84)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_72),
.CI(n_68),
.CON(n_86),
.SN(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_91),
.C(n_84),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_81),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_76),
.B(n_71),
.Y(n_90)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_13),
.B(n_16),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_68),
.C(n_16),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_91),
.C(n_88),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_78),
.B1(n_77),
.B2(n_85),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_93),
.B(n_94),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_95),
.A2(n_90),
.B(n_20),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_100),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_95),
.B(n_15),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_86),
.A3(n_15),
.B1(n_12),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_98),
.B(n_94),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_101),
.Y(n_106)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_102),
.A2(n_104),
.A3(n_8),
.B1(n_10),
.B2(n_4),
.C1(n_2),
.C2(n_3),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_12),
.C(n_6),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_103),
.Y(n_107)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_106),
.B1(n_104),
.B2(n_4),
.C(n_3),
.Y(n_108)
);


endmodule