module real_jpeg_21045_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_184;
wire n_48;
wire n_56;
wire n_164;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_0),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_53),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_72),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_2),
.A2(n_28),
.B1(n_30),
.B2(n_72),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_72),
.Y(n_224)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_4),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_4),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_4),
.A2(n_28),
.B1(n_30),
.B2(n_38),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_5),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_5),
.A2(n_52),
.B(n_119),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_5),
.A2(n_65),
.B1(n_71),
.B2(n_117),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_5),
.B(n_74),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_5),
.A2(n_36),
.B(n_40),
.C(n_179),
.D(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_5),
.B(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_60),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_5),
.A2(n_26),
.B(n_194),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_54),
.B(n_55),
.C(n_128),
.D(n_226),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_5),
.B(n_54),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_6),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_46),
.Y(n_87)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_7),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_7),
.A2(n_122),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_7),
.A2(n_168),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_7),
.A2(n_169),
.B(n_209),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_65),
.B1(n_71),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_52),
.B1(n_54),
.B2(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_76),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_76),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_65),
.B1(n_71),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_11),
.A2(n_52),
.B1(n_54),
.B2(n_96),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_96),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_11),
.A2(n_28),
.B1(n_30),
.B2(n_96),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_31),
.B1(n_36),
.B2(n_37),
.Y(n_82)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_14),
.A2(n_52),
.B1(n_54),
.B2(n_67),
.Y(n_69)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_131),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_129),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_104),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_77),
.B2(n_78),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_48),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_25),
.B(n_34),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_26),
.A2(n_27),
.B(n_32),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_26),
.A2(n_29),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_26),
.A2(n_87),
.B1(n_88),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_26),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_26),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_26),
.B(n_196),
.Y(n_209)
);

NAND2x1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_28),
.A2(n_42),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_30),
.B(n_41),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_30),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_35),
.A2(n_39),
.B1(n_47),
.B2(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_36),
.A2(n_37),
.B1(n_56),
.B2(n_57),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_36),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_37),
.B(n_57),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_39),
.A2(n_45),
.B1(n_47),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_39),
.A2(n_47),
.B1(n_191),
.B2(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_39),
.A2(n_224),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_40),
.B(n_143),
.Y(n_142)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_47),
.A2(n_92),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_47),
.B(n_144),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_47),
.A2(n_142),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_47),
.B(n_117),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_62),
.B2(n_63),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_60),
.B2(n_61),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_51),
.Y(n_99)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_56),
.B(n_59),
.C(n_60),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_55),
.Y(n_126)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_59),
.Y(n_232)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_70),
.B(n_73),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_69),
.B1(n_70),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B(n_68),
.C(n_69),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_67),
.B(n_117),
.C(n_118),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_95),
.B(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_81),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_93),
.C(n_97),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_86),
.B(n_91),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_88),
.A2(n_201),
.B(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_88),
.B(n_117),
.Y(n_214)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_89),
.B(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_100),
.B(n_101),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_103),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_100),
.A2(n_125),
.B1(n_126),
.B2(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_100),
.A2(n_101),
.B(n_150),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.C(n_108),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_107),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_108),
.A2(n_109),
.B1(n_152),
.B2(n_153),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_123),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_111),
.B1(n_123),
.B2(n_124),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_146),
.B(n_147),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_171),
.Y(n_131)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_154),
.B(n_170),
.Y(n_133)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_151),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_139),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.C(n_148),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_140),
.A2(n_141),
.B1(n_148),
.B2(n_149),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_155),
.B(n_157),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_158),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_160),
.A2(n_162),
.B1(n_163),
.B2(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_160),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_164),
.A2(n_165),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_166),
.B(n_167),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_253),
.C(n_254),
.Y(n_171)
);

AOI21x1_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_247),
.B(n_252),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_236),
.B(n_246),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_218),
.B(n_235),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_197),
.B(n_217),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_185),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_177),
.B(n_185),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_179),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_180),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_205),
.B(n_216),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_203),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_215),
.Y(n_205)
);

NOR2xp67_ASAP7_75t_R g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_207),
.B(n_210),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_219),
.B(n_220),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_229),
.B2(n_234),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_223),
.Y(n_228)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_228),
.C(n_234),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_229),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_237),
.B(n_238),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_243),
.C(n_244),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_240),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);


endmodule