module fake_jpeg_30173_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

CKINVDCx16_ASAP7_75t_R g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx5_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_5),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_21),
.B1(n_12),
.B2(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

AND2x6_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_19),
.A2(n_11),
.B1(n_13),
.B2(n_3),
.Y(n_25)
);

AOI21xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_10),
.B(n_14),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_9),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_21),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B1(n_18),
.B2(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

AND2x6_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_34),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_17),
.C(n_19),
.Y(n_39)
);

A2O1A1O1Ixp25_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_33),
.B(n_35),
.C(n_29),
.D(n_24),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_39),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_43),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_37),
.C(n_38),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_33),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_33),
.B(n_1),
.Y(n_47)
);

AOI321xp33_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_6),
.A3(n_30),
.B1(n_34),
.B2(n_15),
.C(n_16),
.Y(n_49)
);

AOI221xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_4),
.B1(n_15),
.B2(n_16),
.C(n_47),
.Y(n_50)
);


endmodule