module fake_aes_841_n_14 (n_1, n_2, n_0, n_14);
input n_1;
input n_2;
input n_0;
output n_14;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
NAND2xp5_ASAP7_75t_L g4 ( .A(n_1), .B(n_2), .Y(n_4) );
INVx3_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
OAI22x1_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_1), .B1(n_2), .B2(n_0), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_3), .B(n_0), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
OR2x6_ASAP7_75t_L g10 ( .A(n_9), .B(n_7), .Y(n_10) );
AOI322xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_4), .A3(n_5), .B1(n_8), .B2(n_7), .C1(n_0), .C2(n_1), .Y(n_11) );
NAND3xp33_ASAP7_75t_L g12 ( .A(n_11), .B(n_10), .C(n_5), .Y(n_12) );
NAND3xp33_ASAP7_75t_L g13 ( .A(n_12), .B(n_10), .C(n_2), .Y(n_13) );
NAND3x1_ASAP7_75t_L g14 ( .A(n_13), .B(n_4), .C(n_11), .Y(n_14) );
endmodule