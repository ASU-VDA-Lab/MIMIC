module fake_jpeg_8470_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_SL g6 ( 
.A(n_0),
.B(n_1),
.Y(n_6)
);

HAxp5_ASAP7_75t_SL g7 ( 
.A(n_5),
.B(n_4),
.CON(n_7),
.SN(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_1),
.B(n_0),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_3),
.B(n_2),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_11),
.B(n_12),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_22),
.Y(n_26)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_7),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_13),
.B1(n_21),
.B2(n_22),
.Y(n_23)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_6),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_25),
.C(n_16),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_14),
.A2(n_13),
.B1(n_18),
.B2(n_17),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_20),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.C(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_36),
.B(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_35),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);


endmodule