module fake_jpeg_28547_n_417 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_417);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_417;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_12),
.B(n_11),
.C(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_5),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

AND2x4_ASAP7_75t_SL g50 ( 
.A(n_20),
.B(n_42),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_20),
.B(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_56),
.B(n_57),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_58),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_0),
.CON(n_60),
.SN(n_60)
);

OAI21xp33_ASAP7_75t_L g117 ( 
.A1(n_60),
.A2(n_32),
.B(n_31),
.Y(n_117)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_14),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_70),
.Y(n_102)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_34),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_14),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_71),
.B(n_41),
.Y(n_105)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_72),
.B(n_73),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_19),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_34),
.B(n_12),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_78),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_42),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_35),
.B(n_0),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

INVx4_ASAP7_75t_SL g81 ( 
.A(n_37),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_86),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_31),
.B(n_1),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_85),
.Y(n_109)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_43),
.B1(n_33),
.B2(n_26),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_89),
.A2(n_110),
.B1(n_1),
.B2(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_99),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_22),
.B1(n_17),
.B2(n_33),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_96),
.A2(n_98),
.B1(n_107),
.B2(n_128),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_50),
.A2(n_22),
.B1(n_17),
.B2(n_33),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_29),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_47),
.A2(n_17),
.B1(n_22),
.B2(n_41),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_104),
.A2(n_18),
.B1(n_86),
.B2(n_69),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_105),
.B(n_131),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_50),
.A2(n_66),
.B1(n_79),
.B2(n_62),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_33),
.B1(n_17),
.B2(n_22),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_16),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_126),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_58),
.B(n_75),
.C(n_18),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_68),
.B(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_18),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_45),
.B(n_39),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_40),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_127),
.B(n_130),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_46),
.A2(n_40),
.B1(n_39),
.B2(n_23),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_23),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_54),
.B(n_16),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_58),
.C(n_37),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_135),
.B(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_137),
.B(n_140),
.Y(n_184)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_121),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_82),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_164),
.C(n_109),
.Y(n_196)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_92),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_74),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_153),
.Y(n_189)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_87),
.B(n_18),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_93),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_18),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_103),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_154),
.B(n_163),
.Y(n_195)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_155),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_88),
.B(n_59),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_88),
.B(n_67),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_118),
.Y(n_158)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_159),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_92),
.A2(n_51),
.B1(n_49),
.B2(n_48),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_123),
.B1(n_119),
.B2(n_108),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_107),
.B1(n_98),
.B2(n_96),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_162),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_91),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_111),
.B(n_85),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_111),
.B1(n_115),
.B2(n_99),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_2),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_167),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_116),
.B(n_3),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_168),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_3),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_176),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_173),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_95),
.B(n_3),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_129),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_179),
.A2(n_184),
.B(n_189),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_196),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_182),
.A2(n_202),
.B1(n_139),
.B2(n_136),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_93),
.B(n_125),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_198),
.B(n_120),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_132),
.B1(n_97),
.B2(n_119),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_203),
.B1(n_206),
.B2(n_143),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_192),
.A2(n_144),
.B1(n_139),
.B2(n_173),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_135),
.A2(n_120),
.B1(n_129),
.B2(n_106),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_109),
.B(n_100),
.Y(n_198)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_154),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_169),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_100),
.B1(n_97),
.B2(n_123),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_156),
.A2(n_132),
.B1(n_108),
.B2(n_120),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_157),
.A2(n_152),
.B1(n_150),
.B2(n_143),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_152),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_225),
.Y(n_251)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_217),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_150),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_218),
.B(n_207),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_221),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_220),
.A2(n_223),
.B1(n_241),
.B2(n_192),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_222),
.B(n_224),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_164),
.B1(n_160),
.B2(n_140),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_148),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_226),
.B(n_227),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_234),
.B1(n_236),
.B2(n_240),
.Y(n_250)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx13_ASAP7_75t_L g230 ( 
.A(n_188),
.Y(n_230)
);

BUFx4f_ASAP7_75t_SL g261 ( 
.A(n_230),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_149),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_247),
.C(n_188),
.Y(n_265)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_137),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_180),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_235),
.A2(n_180),
.B(n_201),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_196),
.A2(n_174),
.B1(n_146),
.B2(n_147),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_163),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_239),
.B(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_204),
.A2(n_142),
.B1(n_158),
.B2(n_144),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_187),
.A2(n_155),
.B1(n_134),
.B2(n_138),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_159),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_185),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_191),
.Y(n_269)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_193),
.Y(n_246)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_168),
.C(n_162),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_264),
.Y(n_281)
);

AOI32xp33_ASAP7_75t_L g253 ( 
.A1(n_216),
.A2(n_198),
.A3(n_214),
.B1(n_203),
.B2(n_201),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_253),
.A2(n_274),
.B(n_276),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_265),
.C(n_268),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_219),
.B(n_193),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_221),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_245),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_234),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_240),
.Y(n_291)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_230),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_267),
.B(n_232),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_210),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_272),
.A2(n_248),
.B1(n_244),
.B2(n_243),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_216),
.A2(n_178),
.B1(n_186),
.B2(n_208),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_228),
.A2(n_178),
.B1(n_191),
.B2(n_210),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_241),
.B1(n_223),
.B2(n_220),
.Y(n_283)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_229),
.Y(n_279)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_280),
.B(n_291),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_283),
.A2(n_286),
.B1(n_272),
.B2(n_259),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_251),
.B(n_225),
.Y(n_284)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g285 ( 
.A(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_285),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_266),
.A2(n_233),
.B1(n_235),
.B2(n_247),
.Y(n_286)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_257),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_293),
.B(n_298),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_254),
.B(n_218),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_300),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_268),
.B(n_248),
.C(n_236),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_238),
.C(n_237),
.Y(n_322)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_251),
.B(n_215),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_262),
.B(n_246),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_311)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_258),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_258),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_304),
.A2(n_250),
.B1(n_264),
.B2(n_278),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_270),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_306),
.A2(n_224),
.B1(n_227),
.B2(n_209),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_322),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_309),
.B(n_310),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_283),
.A2(n_271),
.B1(n_250),
.B2(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_277),
.B1(n_263),
.B2(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_304),
.A2(n_274),
.B1(n_275),
.B2(n_279),
.Y(n_315)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_315),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_299),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_316),
.B(n_281),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_275),
.B1(n_273),
.B2(n_260),
.Y(n_319)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_288),
.A2(n_273),
.B1(n_265),
.B2(n_255),
.Y(n_321)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_323),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_280),
.A2(n_256),
.B1(n_178),
.B2(n_217),
.Y(n_326)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_326),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_281),
.A2(n_209),
.B1(n_186),
.B2(n_208),
.Y(n_327)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_327),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_261),
.B1(n_199),
.B2(n_212),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_330),
.B(n_261),
.Y(n_335)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_333),
.B(n_334),
.Y(n_356)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_318),
.A2(n_284),
.B(n_298),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_335),
.B(n_321),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_317),
.B(n_289),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_341),
.B(n_342),
.Y(n_358)
);

O2A1O1Ixp33_ASAP7_75t_L g342 ( 
.A1(n_314),
.A2(n_282),
.B(n_306),
.C(n_290),
.Y(n_342)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_328),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_343),
.B(n_347),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_329),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_294),
.C(n_282),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_348),
.B(n_303),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_350),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_348),
.B(n_313),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_365),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_353),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g353 ( 
.A(n_345),
.B(n_310),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_332),
.A2(n_319),
.B1(n_312),
.B2(n_318),
.Y(n_354)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_354),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_345),
.B(n_322),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_355),
.B(n_363),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_334),
.B(n_329),
.CI(n_315),
.CON(n_357),
.SN(n_357)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_332),
.A2(n_308),
.B1(n_309),
.B2(n_326),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_361),
.A2(n_346),
.B1(n_338),
.B2(n_336),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_308),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_327),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_335),
.Y(n_374)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_366),
.B(n_367),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_330),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_360),
.A2(n_336),
.B(n_320),
.Y(n_368)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_370),
.A2(n_364),
.B1(n_363),
.B2(n_362),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_358),
.B(n_324),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_374),
.Y(n_388)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_356),
.A2(n_337),
.B(n_338),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_373),
.A2(n_324),
.B(n_325),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_337),
.C(n_344),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_377),
.B(n_379),
.C(n_352),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_353),
.B(n_346),
.C(n_340),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_357),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_383),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_377),
.B(n_372),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_384),
.B(n_391),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_378),
.A2(n_361),
.B1(n_340),
.B2(n_349),
.Y(n_385)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_385),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_370),
.A2(n_359),
.B(n_349),
.Y(n_386)
);

AOI21x1_ASAP7_75t_L g399 ( 
.A1(n_386),
.A2(n_373),
.B(n_375),
.Y(n_399)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_376),
.Y(n_387)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_392),
.Y(n_398)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_390),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_380),
.B(n_325),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_343),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_384),
.B(n_380),
.C(n_375),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_397),
.B(n_399),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_381),
.A2(n_297),
.B1(n_302),
.B2(n_301),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_401),
.B(n_385),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_403),
.B(n_407),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_393),
.A2(n_388),
.B(n_386),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_404),
.A2(n_400),
.B(n_287),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_397),
.B(n_390),
.C(n_305),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_405),
.B(n_406),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_293),
.C(n_292),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_287),
.C(n_212),
.Y(n_407)
);

NAND4xp25_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_401),
.C(n_396),
.D(n_394),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_408),
.A2(n_120),
.B(n_176),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_410),
.A2(n_141),
.B(n_151),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_412),
.A2(n_413),
.B1(n_409),
.B2(n_411),
.Y(n_414)
);

OAI321xp33_ASAP7_75t_L g415 ( 
.A1(n_414),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_415),
.B(n_4),
.Y(n_416)
);

AOI321xp33_ASAP7_75t_L g417 ( 
.A1(n_416),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_9),
.C(n_285),
.Y(n_417)
);


endmodule