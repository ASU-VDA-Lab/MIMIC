module real_jpeg_3988_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_0),
.B(n_82),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_0),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_0),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_0),
.B(n_287),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_0),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_0),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_0),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_1),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_1),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_1),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_1),
.B(n_93),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_1),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_1),
.B(n_339),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_1),
.B(n_407),
.Y(n_406)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_2),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_2),
.Y(n_308)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_2),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_2),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_3),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_3),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_3),
.B(n_38),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_3),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_3),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_3),
.B(n_308),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_3),
.B(n_412),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_82),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_4),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_4),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_4),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_4),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_4),
.B(n_264),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_4),
.B(n_404),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_5),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_5),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_5),
.Y(n_185)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_5),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_6),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_6),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_6),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_6),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_6),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g222 ( 
.A(n_6),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_7),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_7),
.B(n_32),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_7),
.B(n_116),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_7),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_7),
.B(n_253),
.Y(n_414)
);

INVxp33_ASAP7_75t_L g495 ( 
.A(n_8),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_9),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_9),
.Y(n_200)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_10),
.Y(n_492)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_11),
.Y(n_281)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_13),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_14),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_14),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_14),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_14),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_14),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_14),
.B(n_69),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_14),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_14),
.B(n_401),
.Y(n_400)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_16),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_16),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_16),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_16),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_16),
.B(n_38),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_16),
.B(n_377),
.Y(n_376)
);

AND2x4_ASAP7_75t_SL g393 ( 
.A(n_16),
.B(n_394),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_17),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_17),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_17),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_17),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_17),
.B(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_19),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_19),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_19),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_19),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_19),
.B(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_490),
.B(n_493),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_187),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_186),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_146),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_25),
.B(n_146),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_110),
.B2(n_145),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_78),
.C(n_95),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_28),
.B(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_46),
.C(n_59),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_29),
.A2(n_30),
.B1(n_46),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_37),
.C(n_40),
.Y(n_119)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_38),
.Y(n_268)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_39),
.Y(n_402)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_44),
.Y(n_205)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_44),
.Y(n_348)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_45),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g374 ( 
.A(n_45),
.Y(n_374)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_46),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.C(n_56),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_47),
.B(n_56),
.Y(n_166)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_51),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_54),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_55),
.Y(n_288)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_59),
.B(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_66),
.C(n_72),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_62),
.Y(n_228)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_63),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_63),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_63),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_72),
.B2(n_77),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_65),
.A2(n_66),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_114),
.C(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_70),
.Y(n_311)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_71),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_72),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_98),
.C(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_72),
.A2(n_77),
.B1(n_98),
.B2(n_99),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_76),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_95),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_79),
.B(n_84),
.C(n_94),
.Y(n_129)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_94),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_88),
.Y(n_380)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_107),
.C(n_109),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_96),
.A2(n_97),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_157),
.C(n_162),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_98),
.A2(n_99),
.B1(n_162),
.B2(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_101),
.Y(n_223)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_101),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_102),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_106),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_107),
.A2(n_109),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_107),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_173),
.C(n_181),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_107),
.A2(n_170),
.B1(n_181),
.B2(n_182),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.C(n_119),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_115),
.B1(n_138),
.B2(n_139),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_119),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_130),
.B2(n_144),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_142),
.B2(n_143),
.Y(n_130)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_141),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_133),
.Y(n_141)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_147),
.B(n_149),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_151),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_167),
.C(n_172),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_152),
.A2(n_153),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.C(n_165),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_154),
.B(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_156),
.B(n_165),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_167),
.B(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_174),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_180),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_180),
.Y(n_195)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

AO21x1_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_483),
.B(n_488),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_290),
.B(n_482),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_236),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_191),
.B(n_236),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_229),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_192),
.B(n_230),
.C(n_233),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_211),
.C(n_213),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_193),
.B(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.C(n_208),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_194),
.B(n_468),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_196),
.A2(n_197),
.B1(n_208),
.B2(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.C(n_206),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_198),
.B(n_206),
.Y(n_458)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_199),
.Y(n_395)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_201),
.B(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_205),
.Y(n_332)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_205),
.Y(n_407)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_208),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_213),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_224),
.C(n_226),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_214),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.C(n_222),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_215),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_222),
.Y(n_248)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_221),
.Y(n_323)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_221),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_224),
.B(n_226),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_240),
.C(n_243),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_238),
.B(n_241),
.Y(n_478)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_243),
.B(n_478),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_269),
.C(n_272),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_245),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.C(n_258),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_246),
.A2(n_247),
.B1(n_449),
.B2(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_249),
.A2(n_250),
.B(n_254),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_249),
.B(n_258),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_266),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_426)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_266),
.B(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_267),
.B(n_288),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_272),
.Y(n_472)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_286),
.C(n_289),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_274),
.B(n_460),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.C(n_282),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_275),
.B(n_438),
.Y(n_437)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_278),
.A2(n_282),
.B1(n_283),
.B2(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_278),
.Y(n_439)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_286),
.B(n_289),
.Y(n_460)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_476),
.B(n_481),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_463),
.B(n_475),
.Y(n_291)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_445),
.B(n_462),
.Y(n_292)
);

OAI21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_419),
.B(n_444),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_384),
.B(n_418),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_354),
.B(n_383),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_334),
.B(n_353),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_317),
.B(n_333),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_312),
.B(n_316),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_309),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_306),
.Y(n_318)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_319),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_326),
.B2(n_327),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_329),
.C(n_330),
.Y(n_352)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_352),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_352),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_344),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_343),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_343),
.C(n_356),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_341),
.Y(n_359)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_344),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_369),
.C(n_370),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx8_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_357),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_367),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_368),
.C(n_371),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_359),
.B(n_361),
.C(n_362),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_365),
.B2(n_366),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_363),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_366),
.Y(n_388)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_371),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_372),
.B(n_379),
.C(n_381),
.Y(n_416)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_375)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_376),
.Y(n_381)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g382 ( 
.A(n_379),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_417),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_417),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_397),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_396),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_387),
.B(n_396),
.C(n_443),
.Y(n_442)
);

XNOR2x1_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_388),
.B(n_433),
.C(n_434),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_390),
.Y(n_433)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_393),
.Y(n_434)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_408),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_398),
.B(n_410),
.C(n_415),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_406),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_400),
.B(n_403),
.C(n_406),
.Y(n_430)
);

INVx6_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_409),
.A2(n_410),
.B1(n_415),
.B2(n_416),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_414),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_411),
.B(n_414),
.Y(n_429)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_442),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_442),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_431),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_422),
.B(n_423),
.C(n_431),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_427),
.B2(n_428),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_454),
.C(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_429),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_436),
.C(n_441),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_440),
.B2(n_441),
.Y(n_435)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_437),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_461),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_446),
.B(n_461),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_452),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_451),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_448),
.B(n_451),
.C(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_452),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_457),
.C(n_459),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_473),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_464),
.B(n_473),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_466),
.Y(n_464)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_465),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_470),
.C(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_479),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_477),
.B(n_479),
.Y(n_481)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_485),
.B(n_487),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_485),
.B(n_487),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx4f_ASAP7_75t_SL g490 ( 
.A(n_491),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_491),
.Y(n_494)
);

INVx13_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);


endmodule