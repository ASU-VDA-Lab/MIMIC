module fake_netlist_6_988_n_2200 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_661, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_671, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_673, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_669, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_667, n_71, n_74, n_229, n_542, n_644, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_658, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_656, n_96, n_8, n_666, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_653, n_112, n_172, n_648, n_657, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_668, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_662, n_89, n_374, n_659, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_650, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_654, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_652, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_674, n_571, n_268, n_271, n_404, n_651, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_665, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_672, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_655, n_13, n_670, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_110, n_151, n_412, n_640, n_81, n_660, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_663, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_664, n_171, n_192, n_57, n_169, n_51, n_649, n_283, n_2200);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_661;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_671;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_673;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_669;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_667;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_658;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_656;
input n_96;
input n_8;
input n_666;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_653;
input n_112;
input n_172;
input n_648;
input n_657;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_668;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_662;
input n_89;
input n_374;
input n_659;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_650;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_654;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_652;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_674;
input n_571;
input n_268;
input n_271;
input n_404;
input n_651;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_665;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_672;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_655;
input n_13;
input n_670;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_660;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_663;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_664;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2200;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_1380;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_830;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_907;
wire n_1446;
wire n_1815;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_699;
wire n_1986;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_1970;
wire n_2101;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_1064;
wire n_1396;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_697;
wire n_687;
wire n_890;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_851;
wire n_682;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_2069;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_683;
wire n_811;
wire n_1207;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_1993;
wire n_1427;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_995;
wire n_1159;
wire n_1092;
wire n_1060;
wire n_1951;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_775;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_956;
wire n_960;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_1905;
wire n_2016;
wire n_793;
wire n_1593;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_1254;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_1270;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_1667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_1057;
wire n_991;
wire n_1657;
wire n_1126;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2037;
wire n_782;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_1406;
wire n_1332;
wire n_962;
wire n_1041;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_1222;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1640;
wire n_804;
wire n_1846;
wire n_806;
wire n_959;
wire n_879;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_1292;
wire n_1373;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_1716;
wire n_1256;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_924;
wire n_1582;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_1218;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_985;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_1170;
wire n_1629;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2116;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_305),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_143),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_403),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_490),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_276),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_590),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_594),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_478),
.Y(n_683)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_529),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_294),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_436),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_583),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_170),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_524),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_54),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_320),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_575),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_577),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_43),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_586),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_645),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_551),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_488),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_481),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_104),
.Y(n_700)
);

CKINVDCx16_ASAP7_75t_R g701 ( 
.A(n_563),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_510),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_640),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_633),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_319),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_623),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_570),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_189),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_207),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_611),
.Y(n_710)
);

INVx1_ASAP7_75t_SL g711 ( 
.A(n_542),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_607),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_151),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_275),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_360),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_379),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_302),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_409),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_477),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_157),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_27),
.Y(n_721)
);

INVxp67_ASAP7_75t_SL g722 ( 
.A(n_326),
.Y(n_722)
);

INVxp67_ASAP7_75t_L g723 ( 
.A(n_589),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_184),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_247),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_343),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_238),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_651),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_155),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_521),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_672),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_573),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_25),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_246),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_404),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_104),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_608),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_648),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_578),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_12),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_271),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_206),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_613),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_641),
.Y(n_744)
);

BUFx10_ASAP7_75t_L g745 ( 
.A(n_654),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_517),
.Y(n_746)
);

BUFx10_ASAP7_75t_L g747 ( 
.A(n_597),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_549),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_584),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_598),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_23),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_505),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_169),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_46),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_606),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_643),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_615),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_261),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_216),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_486),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_601),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_530),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_614),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_132),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_91),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_512),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_566),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_536),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_288),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_445),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_555),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_66),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_247),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_642),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_12),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_494),
.Y(n_776)
);

BUFx10_ASAP7_75t_L g777 ( 
.A(n_571),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_634),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_649),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_502),
.Y(n_780)
);

CKINVDCx16_ASAP7_75t_R g781 ( 
.A(n_393),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_622),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_595),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_509),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_125),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_284),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_593),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_30),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_511),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_121),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_91),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_628),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_503),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_335),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_576),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_658),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_495),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_610),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_355),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_86),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_451),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_637),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_620),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_561),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_507),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_574),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_346),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_652),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_553),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_653),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_582),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_647),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_621),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_267),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_513),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_70),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_496),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_506),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_527),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_461),
.Y(n_820)
);

BUFx2_ASAP7_75t_SL g821 ( 
.A(n_197),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_635),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_531),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_493),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_8),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_600),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_369),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_657),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_483),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_587),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_548),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_559),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_330),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_285),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_599),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_159),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_619),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_194),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_562),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_655),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_605),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_2),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_499),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_500),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_630),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_222),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_656),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_239),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_44),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_567),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_489),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_646),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_564),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_588),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_508),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_534),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_73),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_639),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_552),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_617),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_165),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_475),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_565),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_419),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_612),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_609),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_64),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_556),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_408),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_467),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_516),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_554),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_250),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_596),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_233),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_665),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_592),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_280),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_580),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_227),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_616),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_270),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_540),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_81),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_558),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_312),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_172),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_631),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_301),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_214),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_662),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_208),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_378),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_400),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_56),
.Y(n_895)
);

INVxp67_ASAP7_75t_L g896 ( 
.A(n_119),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_298),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_7),
.Y(n_898)
);

BUFx10_ASAP7_75t_L g899 ( 
.A(n_585),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_174),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_533),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_632),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_121),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_81),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_458),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_568),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_331),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_358),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_5),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_364),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_602),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_603),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_625),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_37),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_154),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_66),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_541),
.Y(n_917)
);

BUFx2_ASAP7_75t_L g918 ( 
.A(n_638),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_550),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_636),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_417),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_629),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_205),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_572),
.Y(n_924)
);

CKINVDCx16_ASAP7_75t_R g925 ( 
.A(n_624),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_669),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_313),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_547),
.Y(n_928)
);

CKINVDCx20_ASAP7_75t_R g929 ( 
.A(n_535),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_579),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_581),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_604),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_230),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_34),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_53),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_557),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_28),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_591),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_504),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_119),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_627),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_60),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_618),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_569),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_560),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_676),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_821),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_675),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_678),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_725),
.Y(n_950)
);

INVxp67_ASAP7_75t_SL g951 ( 
.A(n_776),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_684),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_725),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_682),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_683),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_725),
.Y(n_956)
);

INVxp67_ASAP7_75t_SL g957 ( 
.A(n_815),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_708),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_688),
.Y(n_959)
);

CKINVDCx20_ASAP7_75t_R g960 ( 
.A(n_696),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_679),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_714),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_720),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_721),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_712),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_727),
.Y(n_966)
);

CKINVDCx20_ASAP7_75t_R g967 ( 
.A(n_717),
.Y(n_967)
);

HB1xp67_ASAP7_75t_L g968 ( 
.A(n_733),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_734),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_742),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_751),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_692),
.Y(n_972)
);

BUFx2_ASAP7_75t_SL g973 ( 
.A(n_728),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_693),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_953),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_950),
.Y(n_976)
);

INVx3_ASAP7_75t_L g977 ( 
.A(n_956),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_961),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_959),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_962),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_951),
.B(n_908),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_963),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_958),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_957),
.B(n_918),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_964),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_966),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_970),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_947),
.B(n_948),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_954),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_971),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_955),
.B(n_677),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_946),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_972),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_974),
.B(n_701),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_946),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_968),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_968),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_969),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_949),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_973),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_952),
.Y(n_1001)
);

OA21x2_ASAP7_75t_L g1002 ( 
.A1(n_960),
.A2(n_681),
.B(n_680),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_965),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_988),
.B(n_732),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_994),
.B(n_718),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_976),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_993),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_976),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_986),
.Y(n_1010)
);

INVx3_ASAP7_75t_L g1011 ( 
.A(n_987),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_995),
.B(n_838),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_1003),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_981),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_991),
.B(n_738),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_987),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_984),
.B(n_738),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_977),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_978),
.Y(n_1019)
);

INVx4_ASAP7_75t_SL g1020 ( 
.A(n_1003),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_1000),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_992),
.B(n_769),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_996),
.B(n_967),
.Y(n_1023)
);

INVx4_ASAP7_75t_L g1024 ( 
.A(n_983),
.Y(n_1024)
);

AND2x6_ASAP7_75t_L g1025 ( 
.A(n_998),
.B(n_881),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_975),
.B(n_978),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_982),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_979),
.B(n_781),
.Y(n_1028)
);

INVx8_ASAP7_75t_L g1029 ( 
.A(n_1001),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_997),
.B(n_755),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_999),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_980),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_1002),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_990),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_1002),
.A2(n_754),
.B1(n_764),
.B2(n_759),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_990),
.B(n_925),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_985),
.Y(n_1037)
);

INVx5_ASAP7_75t_L g1038 ( 
.A(n_975),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_995),
.B(n_880),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_986),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_976),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_988),
.B(n_881),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_989),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_979),
.B(n_699),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_981),
.A2(n_916),
.B1(n_740),
.B2(n_791),
.Y(n_1045)
);

CKINVDCx16_ASAP7_75t_R g1046 ( 
.A(n_1013),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_1016),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1027),
.Y(n_1048)
);

AO22x2_ASAP7_75t_L g1049 ( 
.A1(n_1031),
.A2(n_940),
.B1(n_937),
.B2(n_775),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1019),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1044),
.B(n_753),
.Y(n_1051)
);

AO22x2_ASAP7_75t_L g1052 ( 
.A1(n_1012),
.A2(n_909),
.B1(n_836),
.B2(n_842),
.Y(n_1052)
);

AO22x2_ASAP7_75t_L g1053 ( 
.A1(n_1023),
.A2(n_903),
.B1(n_887),
.B2(n_825),
.Y(n_1053)
);

INVxp67_ASAP7_75t_L g1054 ( 
.A(n_1028),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1032),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_1022),
.B(n_773),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1042),
.B(n_722),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1020),
.B(n_857),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1034),
.Y(n_1059)
);

BUFx8_ASAP7_75t_L g1060 ( 
.A(n_1007),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1010),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1040),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1004),
.B(n_761),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1014),
.A2(n_835),
.B1(n_853),
.B2(n_817),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1026),
.Y(n_1065)
);

OAI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1045),
.A2(n_896),
.B1(n_884),
.B2(n_890),
.C(n_875),
.Y(n_1066)
);

AO22x2_ASAP7_75t_L g1067 ( 
.A1(n_1030),
.A2(n_933),
.B1(n_923),
.B2(n_892),
.Y(n_1067)
);

AND2x2_ASAP7_75t_SL g1068 ( 
.A(n_1039),
.B(n_867),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1037),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1014),
.Y(n_1070)
);

OAI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1017),
.A2(n_934),
.B1(n_914),
.B2(n_898),
.C(n_723),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1006),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_1016),
.Y(n_1073)
);

AO22x2_ASAP7_75t_L g1074 ( 
.A1(n_1005),
.A2(n_833),
.B1(n_744),
.B2(n_711),
.Y(n_1074)
);

AO22x2_ASAP7_75t_L g1075 ( 
.A1(n_1036),
.A2(n_703),
.B1(n_691),
.B2(n_702),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1018),
.Y(n_1076)
);

NAND2x1_ASAP7_75t_L g1077 ( 
.A(n_1011),
.B(n_685),
.Y(n_1077)
);

AO22x2_ASAP7_75t_L g1078 ( 
.A1(n_1035),
.A2(n_1015),
.B1(n_735),
.B2(n_737),
.Y(n_1078)
);

OAI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_1021),
.A2(n_819),
.B1(n_866),
.B2(n_774),
.C(n_749),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1009),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1041),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1024),
.B(n_856),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_1041),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1038),
.Y(n_1084)
);

AOI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1025),
.A2(n_869),
.B1(n_897),
.B2(n_868),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_1029),
.Y(n_1086)
);

AO22x2_ASAP7_75t_L g1087 ( 
.A1(n_1043),
.A2(n_762),
.B1(n_768),
.B2(n_686),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_1029),
.B(n_942),
.C(n_935),
.Y(n_1088)
);

INVxp67_ASAP7_75t_L g1089 ( 
.A(n_1025),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_1038),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_1025),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1042),
.B(n_770),
.Y(n_1092)
);

AO22x2_ASAP7_75t_L g1093 ( 
.A1(n_1031),
.A2(n_780),
.B1(n_786),
.B2(n_782),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1019),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1019),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1019),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1019),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1019),
.Y(n_1098)
);

AO22x2_ASAP7_75t_L g1099 ( 
.A1(n_1031),
.A2(n_801),
.B1(n_808),
.B2(n_805),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1033),
.A2(n_929),
.B1(n_697),
.B2(n_704),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_1044),
.A2(n_689),
.B1(n_747),
.B2(n_745),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1019),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1019),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1013),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1042),
.B(n_811),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1016),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_1044),
.B(n_690),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1019),
.Y(n_1108)
);

INVx1_ASAP7_75t_SL g1109 ( 
.A(n_1031),
.Y(n_1109)
);

AO22x2_ASAP7_75t_L g1110 ( 
.A1(n_1031),
.A2(n_820),
.B1(n_832),
.B2(n_812),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_1022),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1019),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1027),
.Y(n_1113)
);

INVx2_ASAP7_75t_SL g1114 ( 
.A(n_1033),
.Y(n_1114)
);

AO22x2_ASAP7_75t_L g1115 ( 
.A1(n_1031),
.A2(n_841),
.B1(n_847),
.B2(n_837),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1042),
.B(n_854),
.Y(n_1116)
);

AO22x2_ASAP7_75t_L g1117 ( 
.A1(n_1031),
.A2(n_862),
.B1(n_863),
.B2(n_859),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1013),
.Y(n_1118)
);

AO22x2_ASAP7_75t_L g1119 ( 
.A1(n_1031),
.A2(n_874),
.B1(n_876),
.B2(n_872),
.Y(n_1119)
);

NAND2x1p5_ASAP7_75t_L g1120 ( 
.A(n_1008),
.B(n_803),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1045),
.A2(n_913),
.B1(n_889),
.B2(n_901),
.C(n_885),
.Y(n_1121)
);

OA22x2_ASAP7_75t_L g1122 ( 
.A1(n_1014),
.A2(n_694),
.B1(n_709),
.B2(n_700),
.Y(n_1122)
);

NAND2x1p5_ASAP7_75t_L g1123 ( 
.A(n_1008),
.B(n_911),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1042),
.B(n_917),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1016),
.Y(n_1125)
);

AO22x2_ASAP7_75t_L g1126 ( 
.A1(n_1031),
.A2(n_928),
.B1(n_930),
.B2(n_922),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_1044),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_1044),
.B(n_713),
.Y(n_1128)
);

OAI221xp5_ASAP7_75t_L g1129 ( 
.A1(n_1045),
.A2(n_939),
.B1(n_941),
.B2(n_724),
.C(n_741),
.Y(n_1129)
);

AO22x2_ASAP7_75t_L g1130 ( 
.A1(n_1031),
.A2(n_698),
.B1(n_822),
.B2(n_726),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1022),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1019),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1033),
.A2(n_705),
.B1(n_706),
.B2(n_695),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1042),
.B(n_687),
.Y(n_1134)
);

OAI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_1045),
.A2(n_736),
.B1(n_765),
.B2(n_758),
.C(n_729),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1019),
.Y(n_1136)
);

NAND2xp33_ASAP7_75t_SL g1137 ( 
.A(n_1086),
.B(n_707),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1127),
.B(n_710),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1065),
.B(n_716),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1128),
.B(n_719),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1107),
.B(n_1057),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1063),
.B(n_730),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1068),
.B(n_731),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1054),
.B(n_739),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1114),
.B(n_743),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1114),
.B(n_1100),
.Y(n_1146)
);

NAND2xp33_ASAP7_75t_SL g1147 ( 
.A(n_1131),
.B(n_746),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_1109),
.B(n_748),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1133),
.B(n_750),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1050),
.B(n_752),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_SL g1151 ( 
.A(n_1111),
.B(n_756),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1069),
.B(n_840),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_1085),
.B(n_757),
.Y(n_1153)
);

NAND2xp33_ASAP7_75t_SL g1154 ( 
.A(n_1082),
.B(n_760),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1064),
.B(n_1051),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_1061),
.B(n_905),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1062),
.B(n_763),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1070),
.B(n_766),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1136),
.B(n_767),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1055),
.B(n_771),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1059),
.B(n_943),
.Y(n_1161)
);

AND2x4_ASAP7_75t_L g1162 ( 
.A(n_1076),
.B(n_281),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1094),
.B(n_778),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1095),
.B(n_282),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1096),
.B(n_783),
.Y(n_1165)
);

NAND2xp33_ASAP7_75t_SL g1166 ( 
.A(n_1104),
.B(n_784),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_SL g1167 ( 
.A(n_1097),
.B(n_789),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1098),
.B(n_792),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1102),
.B(n_793),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_SL g1170 ( 
.A(n_1118),
.B(n_795),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1056),
.B(n_772),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1103),
.B(n_796),
.Y(n_1172)
);

NAND2xp33_ASAP7_75t_SL g1173 ( 
.A(n_1084),
.B(n_797),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1108),
.B(n_1112),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_1132),
.B(n_798),
.Y(n_1175)
);

NAND2xp33_ASAP7_75t_SL g1176 ( 
.A(n_1090),
.B(n_804),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_1048),
.B(n_806),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_1113),
.B(n_807),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1092),
.B(n_809),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1089),
.B(n_810),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1091),
.B(n_813),
.Y(n_1181)
);

NAND2xp33_ASAP7_75t_SL g1182 ( 
.A(n_1105),
.B(n_1124),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1116),
.B(n_818),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1046),
.B(n_824),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1134),
.B(n_826),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1052),
.B(n_785),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1101),
.B(n_827),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1072),
.B(n_828),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_SL g1189 ( 
.A(n_1081),
.B(n_829),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_SL g1190 ( 
.A(n_1123),
.B(n_830),
.Y(n_1190)
);

NAND2xp33_ASAP7_75t_SL g1191 ( 
.A(n_1073),
.B(n_831),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1075),
.B(n_834),
.Y(n_1192)
);

NAND2xp33_ASAP7_75t_SL g1193 ( 
.A(n_1106),
.B(n_843),
.Y(n_1193)
);

NAND2xp33_ASAP7_75t_SL g1194 ( 
.A(n_1125),
.B(n_844),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1120),
.B(n_845),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_1058),
.B(n_850),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1047),
.B(n_851),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1122),
.B(n_852),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1080),
.B(n_283),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1083),
.B(n_855),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1060),
.B(n_858),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1067),
.B(n_860),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1078),
.B(n_864),
.Y(n_1203)
);

NAND2xp33_ASAP7_75t_SL g1204 ( 
.A(n_1077),
.B(n_865),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1074),
.B(n_870),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1129),
.B(n_871),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1088),
.B(n_877),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1130),
.B(n_883),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1093),
.B(n_886),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1053),
.B(n_888),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1135),
.B(n_891),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1099),
.B(n_893),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1110),
.B(n_894),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1115),
.B(n_902),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1087),
.B(n_286),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1117),
.B(n_906),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1119),
.B(n_907),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1126),
.B(n_910),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1121),
.B(n_912),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1049),
.B(n_919),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1066),
.B(n_920),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1079),
.B(n_921),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_SL g1223 ( 
.A(n_1071),
.B(n_924),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_1127),
.B(n_926),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1086),
.B(n_927),
.Y(n_1225)
);

NAND2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1086),
.B(n_931),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_1127),
.B(n_932),
.Y(n_1227)
);

NAND2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1086),
.B(n_936),
.Y(n_1228)
);

NAND2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1086),
.B(n_938),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1086),
.B(n_944),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1065),
.B(n_945),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1127),
.B(n_689),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1065),
.B(n_685),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1127),
.B(n_745),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1127),
.B(n_747),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1065),
.B(n_685),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_SL g1237 ( 
.A(n_1127),
.B(n_777),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1127),
.B(n_777),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1065),
.B(n_715),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_SL g1240 ( 
.A(n_1127),
.B(n_787),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1127),
.B(n_787),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1065),
.B(n_715),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1127),
.B(n_794),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1127),
.B(n_794),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1127),
.B(n_899),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1127),
.B(n_899),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_SL g1247 ( 
.A(n_1127),
.B(n_779),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1127),
.B(n_779),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1127),
.B(n_779),
.Y(n_1249)
);

NAND2xp33_ASAP7_75t_SL g1250 ( 
.A(n_1086),
.B(n_788),
.Y(n_1250)
);

NAND2xp33_ASAP7_75t_SL g1251 ( 
.A(n_1086),
.B(n_790),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_SL g1252 ( 
.A(n_1127),
.B(n_799),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1127),
.B(n_799),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1127),
.B(n_799),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1127),
.B(n_802),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1127),
.B(n_802),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1127),
.B(n_802),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1065),
.B(n_823),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1127),
.B(n_823),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1065),
.B(n_823),
.Y(n_1260)
);

NAND2xp33_ASAP7_75t_SL g1261 ( 
.A(n_1086),
.B(n_800),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1127),
.B(n_839),
.Y(n_1262)
);

NAND2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1086),
.B(n_814),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1065),
.B(n_879),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1127),
.B(n_879),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1065),
.B(n_816),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_SL g1267 ( 
.A(n_1127),
.B(n_846),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1127),
.B(n_848),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1127),
.B(n_849),
.Y(n_1269)
);

NAND2xp33_ASAP7_75t_SL g1270 ( 
.A(n_1086),
.B(n_861),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1086),
.B(n_873),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1127),
.B(n_878),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1233),
.A2(n_289),
.B(n_287),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1236),
.A2(n_291),
.B(n_290),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1141),
.B(n_882),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1231),
.B(n_895),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_SL g1277 ( 
.A1(n_1239),
.A2(n_293),
.B(n_292),
.Y(n_1277)
);

NOR2x1_ASAP7_75t_R g1278 ( 
.A(n_1215),
.B(n_1201),
.Y(n_1278)
);

NOR2x1_ASAP7_75t_SL g1279 ( 
.A(n_1146),
.B(n_295),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1242),
.A2(n_297),
.B(n_296),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1155),
.B(n_900),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_L g1282 ( 
.A(n_1266),
.B(n_299),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1164),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1258),
.A2(n_303),
.B(n_300),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1152),
.B(n_304),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1174),
.B(n_904),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1162),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1179),
.B(n_915),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1260),
.A2(n_307),
.B(n_306),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1152),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1182),
.A2(n_1139),
.B(n_1185),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1199),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1264),
.A2(n_667),
.A3(n_668),
.B(n_666),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1150),
.A2(n_309),
.B(n_308),
.Y(n_1294)
);

HB1xp67_ASAP7_75t_L g1295 ( 
.A(n_1156),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1161),
.A2(n_311),
.B(n_310),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1180),
.A2(n_315),
.B(n_314),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1142),
.A2(n_317),
.A3(n_318),
.B(n_316),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1171),
.B(n_0),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1162),
.Y(n_1300)
);

O2A1O1Ixp5_ASAP7_75t_L g1301 ( 
.A1(n_1140),
.A2(n_660),
.B(n_661),
.C(n_659),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_SL g1302 ( 
.A1(n_1215),
.A2(n_322),
.B(n_321),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1181),
.A2(n_324),
.B(n_323),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1159),
.A2(n_1165),
.B(n_1160),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1156),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1199),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1163),
.B(n_0),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1188),
.A2(n_327),
.B(n_325),
.Y(n_1308)
);

INVx5_ASAP7_75t_L g1309 ( 
.A(n_1186),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1145),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1177),
.A2(n_329),
.B(n_328),
.Y(n_1311)
);

BUFx4_ASAP7_75t_SL g1312 ( 
.A(n_1250),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1178),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1192),
.A2(n_333),
.A3(n_334),
.B(n_332),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1138),
.B(n_1),
.Y(n_1315)
);

NOR2x1_ASAP7_75t_SL g1316 ( 
.A(n_1167),
.B(n_336),
.Y(n_1316)
);

AOI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1168),
.A2(n_338),
.B(n_337),
.Y(n_1317)
);

NAND2x1_ASAP7_75t_L g1318 ( 
.A(n_1203),
.B(n_339),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1224),
.B(n_2),
.Y(n_1319)
);

OAI22x1_ASAP7_75t_L g1320 ( 
.A1(n_1187),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1169),
.A2(n_341),
.B(n_340),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1172),
.A2(n_1175),
.B(n_1157),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1144),
.Y(n_1323)
);

OR2x2_ASAP7_75t_L g1324 ( 
.A(n_1267),
.B(n_1268),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1269),
.B(n_3),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1221),
.Y(n_1326)
);

AO21x2_ASAP7_75t_L g1327 ( 
.A1(n_1183),
.A2(n_344),
.B(n_342),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1158),
.A2(n_347),
.B(n_345),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1205),
.A2(n_7),
.B1(n_4),
.B2(n_6),
.C(n_8),
.Y(n_1329)
);

OA21x2_ASAP7_75t_L g1330 ( 
.A1(n_1247),
.A2(n_349),
.B(n_348),
.Y(n_1330)
);

AND2x6_ASAP7_75t_L g1331 ( 
.A(n_1202),
.B(n_10),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1209),
.A2(n_670),
.A3(n_671),
.B(n_664),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1211),
.A2(n_351),
.B(n_350),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1190),
.A2(n_353),
.B(n_352),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1206),
.A2(n_356),
.B(n_354),
.Y(n_1335)
);

INVx5_ASAP7_75t_L g1336 ( 
.A(n_1251),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1218),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1272),
.B(n_9),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1208),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1227),
.B(n_9),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1154),
.A2(n_1249),
.A3(n_1252),
.B(n_1248),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1195),
.A2(n_1198),
.B(n_1197),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1253),
.A2(n_359),
.B(n_357),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1143),
.B(n_10),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1254),
.A2(n_362),
.B(n_361),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1255),
.A2(n_365),
.B(n_363),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1149),
.A2(n_367),
.B(n_366),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1256),
.A2(n_370),
.B(n_368),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1257),
.A2(n_674),
.A3(n_372),
.B(n_373),
.Y(n_1349)
);

NOR2x1_ASAP7_75t_SL g1350 ( 
.A(n_1259),
.B(n_371),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1153),
.A2(n_375),
.B1(n_376),
.B2(n_374),
.Y(n_1351)
);

NOR4xp25_ASAP7_75t_L g1352 ( 
.A(n_1220),
.B(n_14),
.C(n_11),
.D(n_13),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1148),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1166),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1262),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1184),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1200),
.A2(n_380),
.B(n_377),
.Y(n_1357)
);

AOI221xp5_ASAP7_75t_L g1358 ( 
.A1(n_1212),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.C(n_17),
.Y(n_1358)
);

AOI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1265),
.A2(n_382),
.B(n_381),
.Y(n_1359)
);

BUFx8_ASAP7_75t_L g1360 ( 
.A(n_1261),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1232),
.B(n_383),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1213),
.B(n_15),
.Y(n_1362)
);

CKINVDCx20_ASAP7_75t_R g1363 ( 
.A(n_1170),
.Y(n_1363)
);

AOI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1207),
.A2(n_385),
.B(n_384),
.Y(n_1364)
);

AND2x6_ASAP7_75t_L g1365 ( 
.A(n_1210),
.B(n_1214),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1234),
.Y(n_1366)
);

AND2x4_ASAP7_75t_L g1367 ( 
.A(n_1196),
.B(n_1235),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1219),
.A2(n_387),
.B(n_386),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1222),
.A2(n_389),
.B(n_388),
.Y(n_1369)
);

BUFx5_ASAP7_75t_L g1370 ( 
.A(n_1173),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1216),
.A2(n_1217),
.B(n_1237),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1238),
.A2(n_391),
.B(n_390),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1326),
.A2(n_1241),
.B(n_1240),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1275),
.B(n_1243),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1281),
.A2(n_1223),
.B1(n_1245),
.B2(n_1244),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1305),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1292),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1287),
.B(n_1246),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1369),
.A2(n_1176),
.B(n_1189),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1286),
.B(n_1151),
.Y(n_1380)
);

OAI222xp33_ASAP7_75t_L g1381 ( 
.A1(n_1325),
.A2(n_18),
.B1(n_20),
.B2(n_16),
.C1(n_17),
.C2(n_19),
.Y(n_1381)
);

INVxp33_ASAP7_75t_L g1382 ( 
.A(n_1278),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1360),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1276),
.B(n_1147),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1288),
.B(n_1263),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1295),
.Y(n_1386)
);

INVxp67_ASAP7_75t_SL g1387 ( 
.A(n_1283),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1291),
.A2(n_1193),
.B(n_1191),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1279),
.A2(n_1204),
.A3(n_1194),
.B(n_1137),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1294),
.A2(n_1226),
.B(n_1225),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1307),
.A2(n_1229),
.B(n_1228),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1324),
.B(n_1270),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1309),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1296),
.A2(n_1230),
.B(n_1271),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1336),
.Y(n_1395)
);

OR2x6_ASAP7_75t_L g1396 ( 
.A(n_1302),
.B(n_392),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1300),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1303),
.A2(n_395),
.B(n_394),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1273),
.A2(n_397),
.B(n_396),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1274),
.A2(n_399),
.B(n_398),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1313),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1336),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1280),
.A2(n_1289),
.B(n_1284),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1355),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1308),
.A2(n_402),
.B(n_401),
.Y(n_1406)
);

INVx3_ASAP7_75t_SL g1407 ( 
.A(n_1363),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1299),
.B(n_18),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1311),
.A2(n_406),
.B(n_405),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1290),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1334),
.A2(n_410),
.B(n_407),
.Y(n_1411)
);

INVxp67_ASAP7_75t_SL g1412 ( 
.A(n_1323),
.Y(n_1412)
);

HB1xp67_ASAP7_75t_L g1413 ( 
.A(n_1339),
.Y(n_1413)
);

NAND2x1p5_ASAP7_75t_L g1414 ( 
.A(n_1354),
.B(n_414),
.Y(n_1414)
);

A2O1A1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1304),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_1415)
);

CKINVDCx6p67_ASAP7_75t_R g1416 ( 
.A(n_1320),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1364),
.A2(n_412),
.B(n_411),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1285),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1322),
.A2(n_415),
.B(n_413),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1353),
.B(n_416),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_L g1421 ( 
.A(n_1356),
.B(n_21),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1344),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1333),
.A2(n_420),
.B(n_418),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1310),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1342),
.A2(n_422),
.B(n_421),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1317),
.Y(n_1426)
);

OA21x2_ASAP7_75t_L g1427 ( 
.A1(n_1335),
.A2(n_424),
.B(n_423),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1362),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1366),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1359),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1368),
.A2(n_426),
.B(n_425),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1315),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1301),
.A2(n_428),
.B(n_427),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1319),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1337),
.B(n_22),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1367),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1343),
.A2(n_430),
.B(n_429),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1340),
.Y(n_1438)
);

INVx3_ASAP7_75t_L g1439 ( 
.A(n_1371),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1345),
.A2(n_432),
.B(n_431),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1358),
.A2(n_1329),
.B1(n_1338),
.B2(n_1365),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1372),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1365),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1346),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1331),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1348),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1318),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1282),
.A2(n_434),
.B(n_433),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1341),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1312),
.Y(n_1450)
);

OA21x2_ASAP7_75t_L g1451 ( 
.A1(n_1347),
.A2(n_1297),
.B(n_1277),
.Y(n_1451)
);

NAND2x1p5_ASAP7_75t_L g1452 ( 
.A(n_1361),
.B(n_437),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1331),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1316),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1350),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_SL g1456 ( 
.A(n_1327),
.B(n_35),
.Y(n_1456)
);

NOR2xp67_ASAP7_75t_SL g1457 ( 
.A(n_1328),
.B(n_36),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1349),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1321),
.A2(n_438),
.B(n_435),
.Y(n_1459)
);

AOI21xp33_ASAP7_75t_L g1460 ( 
.A1(n_1351),
.A2(n_37),
.B(n_38),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1330),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1349),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_SL g1463 ( 
.A(n_1370),
.B(n_439),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1357),
.A2(n_441),
.B(n_440),
.Y(n_1464)
);

CKINVDCx14_ASAP7_75t_R g1465 ( 
.A(n_1370),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1298),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1293),
.A2(n_443),
.B(n_442),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1352),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1314),
.Y(n_1469)
);

OAI222xp33_ASAP7_75t_L g1470 ( 
.A1(n_1332),
.A2(n_41),
.B1(n_43),
.B2(n_39),
.C1(n_40),
.C2(n_42),
.Y(n_1470)
);

AOI22x1_ASAP7_75t_L g1471 ( 
.A1(n_1314),
.A2(n_446),
.B1(n_447),
.B2(n_444),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1293),
.A2(n_44),
.B1(n_41),
.B2(n_42),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1306),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1369),
.A2(n_449),
.B(n_448),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1306),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1306),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1369),
.A2(n_452),
.B(n_450),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1306),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1369),
.A2(n_454),
.B(n_453),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1369),
.A2(n_456),
.B(n_455),
.Y(n_1480)
);

CKINVDCx8_ASAP7_75t_R g1481 ( 
.A(n_1336),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1412),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1424),
.Y(n_1483)
);

OA21x2_ASAP7_75t_L g1484 ( 
.A1(n_1466),
.A2(n_459),
.B(n_457),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1449),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1393),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1404),
.A2(n_462),
.B(n_460),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1401),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1405),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1408),
.B(n_45),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1441),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1376),
.Y(n_1492)
);

OAI211xp5_ASAP7_75t_L g1493 ( 
.A1(n_1443),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1425),
.A2(n_464),
.B(n_463),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1403),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1476),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1474),
.A2(n_466),
.B(n_465),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1374),
.B(n_468),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1395),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1436),
.A2(n_57),
.B1(n_65),
.B2(n_49),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1429),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1473),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1475),
.Y(n_1503)
);

AO21x2_ASAP7_75t_L g1504 ( 
.A1(n_1458),
.A2(n_470),
.B(n_469),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1438),
.B(n_50),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1478),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1397),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1462),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1428),
.B(n_50),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1410),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_472),
.B(n_471),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1432),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1418),
.B(n_473),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1434),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1439),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1479),
.A2(n_476),
.B(n_474),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1402),
.B(n_479),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1385),
.B(n_51),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1426),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1435),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1460),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1442),
.A2(n_482),
.B(n_480),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1430),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1392),
.B(n_54),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1387),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1455),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1454),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1480),
.A2(n_1400),
.B(n_1399),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1469),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1416),
.B(n_55),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1417),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1469),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1386),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1406),
.A2(n_485),
.B(n_484),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1467),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1444),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1446),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1461),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1421),
.B(n_55),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1481),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1375),
.B(n_56),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1464),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1413),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1447),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1468),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1471),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1384),
.B(n_57),
.Y(n_1547)
);

XOR2xp5_ASAP7_75t_L g1548 ( 
.A(n_1501),
.B(n_1450),
.Y(n_1548)
);

NAND2xp33_ASAP7_75t_R g1549 ( 
.A(n_1517),
.B(n_1378),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1545),
.B(n_1407),
.Y(n_1550)
);

XNOR2xp5_ASAP7_75t_L g1551 ( 
.A(n_1486),
.B(n_1382),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1499),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_R g1553 ( 
.A(n_1540),
.B(n_1465),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1520),
.B(n_1380),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_1543),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1533),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1508),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1373),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1498),
.B(n_1391),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_R g1560 ( 
.A(n_1495),
.B(n_1383),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1525),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1513),
.B(n_1377),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_1530),
.Y(n_1563)
);

OR2x6_ASAP7_75t_L g1564 ( 
.A(n_1517),
.B(n_1396),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_SL g1565 ( 
.A(n_1518),
.B(n_1414),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1539),
.B(n_1445),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1509),
.B(n_1453),
.Y(n_1567)
);

NAND2xp33_ASAP7_75t_R g1568 ( 
.A(n_1524),
.B(n_1420),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1508),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1507),
.Y(n_1570)
);

XOR2xp5_ASAP7_75t_L g1571 ( 
.A(n_1547),
.B(n_1452),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_R g1572 ( 
.A(n_1545),
.B(n_1377),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1514),
.B(n_1422),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1510),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1513),
.B(n_1396),
.Y(n_1575)
);

INVx8_ASAP7_75t_L g1576 ( 
.A(n_1505),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1502),
.Y(n_1577)
);

XNOR2xp5_ASAP7_75t_L g1578 ( 
.A(n_1490),
.B(n_1472),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1503),
.B(n_1415),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1544),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1483),
.B(n_1447),
.Y(n_1581)
);

AND2x4_ASAP7_75t_L g1582 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1492),
.B(n_1389),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1582),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1550),
.B(n_1526),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1556),
.B(n_1527),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1558),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1569),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1561),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1574),
.B(n_1496),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1583),
.B(n_1529),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1577),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_SL g1594 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1570),
.B(n_1482),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1555),
.B(n_1506),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1564),
.B(n_1529),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1581),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1579),
.Y(n_1599)
);

NOR3xp33_ASAP7_75t_SL g1600 ( 
.A(n_1559),
.B(n_1381),
.C(n_1493),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1565),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1571),
.B(n_1566),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1575),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1519),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1562),
.B(n_1515),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1580),
.B(n_1515),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1485),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1576),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1551),
.B(n_1500),
.Y(n_1610)
);

INVx2_ASAP7_75t_SL g1611 ( 
.A(n_1552),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1578),
.B(n_1523),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1572),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1564),
.B(n_1532),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1553),
.Y(n_1615)
);

NOR3xp33_ASAP7_75t_SL g1616 ( 
.A(n_1549),
.B(n_1470),
.C(n_1491),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1563),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1548),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1560),
.Y(n_1619)
);

BUFx2_ASAP7_75t_L g1620 ( 
.A(n_1568),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1582),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1552),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1602),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1620),
.B(n_1485),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1588),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1589),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1604),
.B(n_1536),
.Y(n_1627)
);

NOR3xp33_ASAP7_75t_SL g1628 ( 
.A(n_1594),
.B(n_1456),
.C(n_1448),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1604),
.B(n_1536),
.Y(n_1629)
);

OAI221xp5_ASAP7_75t_L g1630 ( 
.A1(n_1600),
.A2(n_1521),
.B1(n_1457),
.B2(n_1419),
.C(n_1431),
.Y(n_1630)
);

OR2x2_ASAP7_75t_SL g1631 ( 
.A(n_1613),
.B(n_1484),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_SL g1632 ( 
.A(n_1619),
.B(n_1538),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1593),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1609),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1602),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1587),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1616),
.B(n_1546),
.C(n_1535),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1603),
.B(n_1537),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1595),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1601),
.B(n_1546),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1599),
.B(n_1601),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1591),
.Y(n_1642)
);

AOI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1610),
.A2(n_1451),
.B1(n_1427),
.B2(n_1423),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1608),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1590),
.B(n_1504),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1585),
.B(n_1522),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1586),
.Y(n_1648)
);

INVxp33_ASAP7_75t_L g1649 ( 
.A(n_1618),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1584),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1612),
.A2(n_1484),
.B1(n_1531),
.B2(n_1459),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1621),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1615),
.A2(n_1388),
.B1(n_1394),
.B2(n_1390),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1596),
.B(n_1487),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1605),
.B(n_1528),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1597),
.Y(n_1656)
);

AOI21xp33_ASAP7_75t_L g1657 ( 
.A1(n_1598),
.A2(n_1379),
.B(n_1497),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1597),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1614),
.A2(n_1433),
.B1(n_1494),
.B2(n_1511),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1614),
.A2(n_1534),
.B1(n_1516),
.B2(n_1398),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1592),
.B(n_1411),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1607),
.B(n_1463),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1606),
.Y(n_1663)
);

OAI211xp5_ASAP7_75t_SL g1664 ( 
.A1(n_1619),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1611),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1622),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1617),
.A2(n_1409),
.B(n_1437),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1592),
.B(n_1440),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1620),
.B(n_1389),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1620),
.B(n_58),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1620),
.B(n_59),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1590),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1588),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1611),
.Y(n_1674)
);

NAND4xp25_ASAP7_75t_L g1675 ( 
.A(n_1594),
.B(n_63),
.C(n_61),
.D(n_62),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1602),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1587),
.B(n_61),
.Y(n_1677)
);

BUFx3_ASAP7_75t_L g1678 ( 
.A(n_1590),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1587),
.B(n_62),
.Y(n_1679)
);

INVx1_ASAP7_75t_SL g1680 ( 
.A(n_1590),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1588),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1620),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1620),
.B(n_67),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1635),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1625),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1626),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1656),
.B(n_67),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1658),
.B(n_1663),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1639),
.B(n_68),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1645),
.B(n_68),
.Y(n_1690)
);

INVx1_ASAP7_75t_SL g1691 ( 
.A(n_1680),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1636),
.B(n_69),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1673),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1675),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1644),
.B(n_71),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1681),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1623),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1676),
.Y(n_1698)
);

AOI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1664),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.C(n_76),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1642),
.B(n_74),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1672),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1650),
.B(n_75),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1638),
.B(n_76),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1641),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1652),
.B(n_77),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1633),
.Y(n_1706)
);

AND2x4_ASAP7_75t_SL g1707 ( 
.A(n_1674),
.B(n_644),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1648),
.B(n_77),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1627),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1624),
.B(n_78),
.Y(n_1710)
);

OR2x2_ASAP7_75t_L g1711 ( 
.A(n_1655),
.B(n_78),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1677),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1678),
.B(n_1634),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1640),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1679),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1649),
.B(n_1674),
.Y(n_1716)
);

NAND2xp67_ASAP7_75t_L g1717 ( 
.A(n_1671),
.B(n_79),
.Y(n_1717)
);

OR2x6_ASAP7_75t_L g1718 ( 
.A(n_1674),
.B(n_79),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1669),
.B(n_80),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1632),
.B(n_80),
.Y(n_1720)
);

OAI332xp33_ASAP7_75t_L g1721 ( 
.A1(n_1670),
.A2(n_108),
.A3(n_90),
.B1(n_125),
.B2(n_116),
.B3(n_132),
.C1(n_99),
.C2(n_82),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1646),
.B(n_82),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1629),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1665),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1647),
.B(n_83),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1666),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1654),
.B(n_83),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1683),
.B(n_84),
.Y(n_1728)
);

AND2x4_ASAP7_75t_L g1729 ( 
.A(n_1662),
.B(n_84),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1661),
.B(n_1668),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1631),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1637),
.B(n_85),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1668),
.B(n_1653),
.Y(n_1733)
);

AOI21xp33_ASAP7_75t_L g1734 ( 
.A1(n_1630),
.A2(n_85),
.B(n_86),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1651),
.B(n_87),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1643),
.B(n_87),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1628),
.B(n_88),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1682),
.A2(n_90),
.B1(n_88),
.B2(n_89),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1667),
.B(n_1657),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1659),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1660),
.B(n_89),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1635),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1680),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1639),
.B(n_92),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1635),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1656),
.B(n_93),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1635),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1656),
.B(n_93),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1635),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1639),
.B(n_94),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1639),
.B(n_94),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1656),
.B(n_95),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1623),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1635),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1656),
.B(n_96),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1656),
.B(n_96),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1656),
.B(n_97),
.Y(n_1757)
);

AND2x4_ASAP7_75t_SL g1758 ( 
.A(n_1674),
.B(n_650),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1639),
.B(n_97),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1684),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1714),
.B(n_98),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1712),
.B(n_98),
.Y(n_1762)
);

AO221x2_ASAP7_75t_L g1763 ( 
.A1(n_1731),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.C(n_102),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1701),
.Y(n_1764)
);

BUFx2_ASAP7_75t_L g1765 ( 
.A(n_1753),
.Y(n_1765)
);

AO221x2_ASAP7_75t_L g1766 ( 
.A1(n_1719),
.A2(n_102),
.B1(n_105),
.B2(n_101),
.C(n_103),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1713),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1742),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1688),
.B(n_100),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1691),
.Y(n_1770)
);

INVxp67_ASAP7_75t_L g1771 ( 
.A(n_1725),
.Y(n_1771)
);

INVxp67_ASAP7_75t_SL g1772 ( 
.A(n_1698),
.Y(n_1772)
);

NAND2xp33_ASAP7_75t_SL g1773 ( 
.A(n_1720),
.B(n_106),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_SL g1774 ( 
.A(n_1732),
.B(n_107),
.Y(n_1774)
);

INVxp33_ASAP7_75t_SL g1775 ( 
.A(n_1743),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1715),
.B(n_108),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1740),
.B(n_109),
.Y(n_1777)
);

NAND2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1687),
.B(n_110),
.Y(n_1778)
);

NOR2x1_ASAP7_75t_L g1779 ( 
.A(n_1716),
.B(n_110),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1718),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_SL g1781 ( 
.A1(n_1718),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1726),
.Y(n_1782)
);

AO221x2_ASAP7_75t_L g1783 ( 
.A1(n_1721),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.C(n_114),
.Y(n_1783)
);

AO221x2_ASAP7_75t_L g1784 ( 
.A1(n_1728),
.A2(n_116),
.B1(n_114),
.B2(n_115),
.C(n_117),
.Y(n_1784)
);

CKINVDCx20_ASAP7_75t_R g1785 ( 
.A(n_1707),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1697),
.B(n_115),
.Y(n_1786)
);

INVx1_ASAP7_75t_SL g1787 ( 
.A(n_1689),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1724),
.B(n_117),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1730),
.B(n_118),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1704),
.B(n_118),
.Y(n_1790)
);

AO221x2_ASAP7_75t_L g1791 ( 
.A1(n_1744),
.A2(n_1759),
.B1(n_1750),
.B2(n_1737),
.C(n_1736),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1699),
.A2(n_123),
.B1(n_120),
.B2(n_122),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1711),
.B(n_122),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_L g1794 ( 
.A1(n_1694),
.A2(n_127),
.B1(n_124),
.B2(n_126),
.C(n_128),
.Y(n_1794)
);

AO221x2_ASAP7_75t_L g1795 ( 
.A1(n_1703),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.C(n_130),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1717),
.B(n_129),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1745),
.B(n_131),
.Y(n_1797)
);

NAND2xp33_ASAP7_75t_SL g1798 ( 
.A(n_1746),
.B(n_133),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1747),
.B(n_134),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1749),
.B(n_134),
.Y(n_1800)
);

NAND2xp33_ASAP7_75t_SL g1801 ( 
.A(n_1748),
.B(n_135),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1754),
.B(n_136),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1739),
.B(n_136),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1709),
.B(n_137),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1685),
.B(n_137),
.Y(n_1805)
);

NOR2xp33_ASAP7_75t_L g1806 ( 
.A(n_1751),
.B(n_138),
.Y(n_1806)
);

AO221x2_ASAP7_75t_L g1807 ( 
.A1(n_1692),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.C(n_141),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1686),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1729),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1727),
.B(n_140),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_L g1811 ( 
.A(n_1693),
.B(n_141),
.Y(n_1811)
);

NOR2x1_ASAP7_75t_L g1812 ( 
.A(n_1735),
.B(n_142),
.Y(n_1812)
);

AO221x2_ASAP7_75t_L g1813 ( 
.A1(n_1696),
.A2(n_1723),
.B1(n_1706),
.B2(n_1741),
.C(n_1722),
.Y(n_1813)
);

NOR2xp33_ASAP7_75t_L g1814 ( 
.A(n_1752),
.B(n_142),
.Y(n_1814)
);

AOI22xp5_ASAP7_75t_L g1815 ( 
.A1(n_1733),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_1815)
);

CKINVDCx8_ASAP7_75t_R g1816 ( 
.A(n_1690),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1755),
.B(n_144),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1756),
.Y(n_1818)
);

AO221x2_ASAP7_75t_L g1819 ( 
.A1(n_1757),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.C(n_148),
.Y(n_1819)
);

NAND2xp33_ASAP7_75t_SL g1820 ( 
.A(n_1710),
.B(n_146),
.Y(n_1820)
);

AO221x2_ASAP7_75t_L g1821 ( 
.A1(n_1708),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_152),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1695),
.Y(n_1822)
);

OAI221xp5_ASAP7_75t_L g1823 ( 
.A1(n_1738),
.A2(n_1700),
.B1(n_1705),
.B2(n_1702),
.C(n_1758),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1705),
.Y(n_1824)
);

OAI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1734),
.A2(n_152),
.B1(n_149),
.B2(n_150),
.C(n_153),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1699),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1714),
.B(n_158),
.Y(n_1827)
);

AOI21xp33_ASAP7_75t_L g1828 ( 
.A1(n_1739),
.A2(n_160),
.B(n_161),
.Y(n_1828)
);

AO221x2_ASAP7_75t_L g1829 ( 
.A1(n_1731),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1714),
.B(n_162),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1714),
.B(n_166),
.Y(n_1831)
);

CKINVDCx20_ASAP7_75t_R g1832 ( 
.A(n_1701),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1684),
.Y(n_1833)
);

NAND2x1_ASAP7_75t_L g1834 ( 
.A(n_1731),
.B(n_167),
.Y(n_1834)
);

INVxp67_ASAP7_75t_L g1835 ( 
.A(n_1725),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1712),
.B(n_168),
.Y(n_1836)
);

OAI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1735),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1712),
.B(n_171),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1714),
.B(n_172),
.Y(n_1839)
);

NOR2x1_ASAP7_75t_L g1840 ( 
.A(n_1701),
.B(n_173),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1714),
.B(n_173),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1714),
.B(n_175),
.Y(n_1842)
);

NAND2xp33_ASAP7_75t_SL g1843 ( 
.A(n_1720),
.B(n_176),
.Y(n_1843)
);

AOI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1699),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1770),
.Y(n_1845)
);

NOR2x1_ASAP7_75t_L g1846 ( 
.A(n_1811),
.B(n_177),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1791),
.B(n_178),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1791),
.B(n_179),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1771),
.B(n_180),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1782),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1760),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1783),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1835),
.B(n_181),
.Y(n_1853)
);

INVx1_ASAP7_75t_SL g1854 ( 
.A(n_1775),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1779),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1768),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1832),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1765),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1833),
.Y(n_1859)
);

HB1xp67_ASAP7_75t_L g1860 ( 
.A(n_1808),
.Y(n_1860)
);

INVxp67_ASAP7_75t_L g1861 ( 
.A(n_1840),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1787),
.B(n_183),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1780),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1824),
.Y(n_1864)
);

AND3x2_ASAP7_75t_L g1865 ( 
.A(n_1796),
.B(n_184),
.C(n_185),
.Y(n_1865)
);

INVx3_ASAP7_75t_L g1866 ( 
.A(n_1764),
.Y(n_1866)
);

INVx1_ASAP7_75t_SL g1867 ( 
.A(n_1818),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1772),
.B(n_185),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1777),
.B(n_186),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1822),
.B(n_186),
.Y(n_1870)
);

AND2x2_ASAP7_75t_L g1871 ( 
.A(n_1789),
.B(n_1804),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1761),
.B(n_187),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1790),
.B(n_188),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1786),
.B(n_188),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1816),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_SL g1876 ( 
.A(n_1815),
.B(n_190),
.C(n_191),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1827),
.B(n_192),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1830),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1831),
.Y(n_1879)
);

OR2x6_ASAP7_75t_L g1880 ( 
.A(n_1812),
.B(n_193),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1788),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1839),
.B(n_194),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1841),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1842),
.B(n_195),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1809),
.Y(n_1885)
);

INVx3_ASAP7_75t_L g1886 ( 
.A(n_1763),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1797),
.B(n_195),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1799),
.B(n_196),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1800),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1802),
.Y(n_1890)
);

INVx1_ASAP7_75t_SL g1891 ( 
.A(n_1785),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1805),
.B(n_198),
.Y(n_1892)
);

NOR2x1_ASAP7_75t_L g1893 ( 
.A(n_1762),
.B(n_1776),
.Y(n_1893)
);

INVx1_ASAP7_75t_SL g1894 ( 
.A(n_1778),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1798),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1793),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1803),
.B(n_198),
.Y(n_1897)
);

NOR2x1_ASAP7_75t_L g1898 ( 
.A(n_1806),
.B(n_199),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1836),
.B(n_199),
.Y(n_1899)
);

HB1xp67_ASAP7_75t_L g1900 ( 
.A(n_1763),
.Y(n_1900)
);

INVxp67_ASAP7_75t_L g1901 ( 
.A(n_1801),
.Y(n_1901)
);

BUFx3_ASAP7_75t_L g1902 ( 
.A(n_1814),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1838),
.B(n_200),
.Y(n_1903)
);

NOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1817),
.B(n_1810),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1829),
.B(n_200),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_L g1906 ( 
.A(n_1783),
.B(n_201),
.C(n_202),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1829),
.B(n_201),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1807),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1821),
.B(n_202),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1807),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1784),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1823),
.B(n_1784),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1819),
.B(n_203),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1766),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1795),
.B(n_203),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1820),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1828),
.B(n_204),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1773),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1826),
.B(n_204),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1843),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1837),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1794),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1844),
.B(n_205),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1825),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1760),
.Y(n_1925)
);

NOR2xp33_ASAP7_75t_L g1926 ( 
.A(n_1775),
.B(n_209),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1813),
.B(n_210),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1767),
.B(n_210),
.Y(n_1928)
);

INVx2_ASAP7_75t_SL g1929 ( 
.A(n_1770),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1791),
.B(n_211),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1760),
.Y(n_1931)
);

INVx2_ASAP7_75t_SL g1932 ( 
.A(n_1770),
.Y(n_1932)
);

AOI22xp33_ASAP7_75t_L g1933 ( 
.A1(n_1783),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1775),
.B(n_212),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1783),
.A2(n_213),
.B(n_215),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1771),
.B(n_215),
.Y(n_1936)
);

OAI21xp33_ASAP7_75t_L g1937 ( 
.A1(n_1792),
.A2(n_216),
.B(n_217),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1771),
.B(n_217),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1760),
.Y(n_1939)
);

NAND3xp33_ASAP7_75t_L g1940 ( 
.A(n_1783),
.B(n_218),
.C(n_219),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1782),
.Y(n_1941)
);

OAI221xp5_ASAP7_75t_L g1942 ( 
.A1(n_1774),
.A2(n_220),
.B1(n_218),
.B2(n_219),
.C(n_221),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1760),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1813),
.B(n_220),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1775),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1760),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1775),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1813),
.B(n_223),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1775),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1771),
.B(n_224),
.Y(n_1950)
);

AOI222xp33_ASAP7_75t_L g1951 ( 
.A1(n_1781),
.A2(n_226),
.B1(n_228),
.B2(n_224),
.C1(n_225),
.C2(n_227),
.Y(n_1951)
);

INVx1_ASAP7_75t_SL g1952 ( 
.A(n_1775),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1791),
.B(n_225),
.Y(n_1953)
);

INVx1_ASAP7_75t_SL g1954 ( 
.A(n_1775),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1782),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1760),
.Y(n_1956)
);

BUFx2_ASAP7_75t_L g1957 ( 
.A(n_1765),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1760),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1791),
.B(n_229),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1760),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_SL g1961 ( 
.A(n_1834),
.B(n_229),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1771),
.B(n_230),
.Y(n_1962)
);

INVx5_ASAP7_75t_L g1963 ( 
.A(n_1769),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1771),
.B(n_231),
.Y(n_1964)
);

INVx1_ASAP7_75t_SL g1965 ( 
.A(n_1775),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1760),
.Y(n_1966)
);

HB1xp67_ASAP7_75t_L g1967 ( 
.A(n_1765),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1771),
.B(n_231),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1791),
.B(n_232),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1771),
.B(n_232),
.Y(n_1970)
);

OAI221xp5_ASAP7_75t_L g1971 ( 
.A1(n_1774),
.A2(n_236),
.B1(n_234),
.B2(n_235),
.C(n_237),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1860),
.Y(n_1972)
);

NAND3xp33_ASAP7_75t_L g1973 ( 
.A(n_1906),
.B(n_235),
.C(n_236),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1858),
.B(n_237),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1851),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1866),
.B(n_238),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1900),
.B(n_239),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1864),
.B(n_240),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1940),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1886),
.B(n_242),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1855),
.B(n_243),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1856),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1859),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1925),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1967),
.B(n_1957),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1931),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1939),
.Y(n_1987)
);

NAND2x1_ASAP7_75t_L g1988 ( 
.A(n_1845),
.B(n_243),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1852),
.A2(n_246),
.B1(n_244),
.B2(n_245),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1875),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1929),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1846),
.Y(n_1992)
);

NOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1927),
.B(n_245),
.Y(n_1993)
);

AOI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1922),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_1994)
);

OAI21xp5_ASAP7_75t_L g1995 ( 
.A1(n_1935),
.A2(n_248),
.B(n_249),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1943),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1946),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1924),
.A2(n_251),
.B(n_252),
.Y(n_1998)
);

OAI322xp33_ASAP7_75t_L g1999 ( 
.A1(n_1912),
.A2(n_251),
.A3(n_252),
.B1(n_253),
.B2(n_254),
.C1(n_255),
.C2(n_256),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1956),
.Y(n_2000)
);

OAI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1933),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1958),
.Y(n_2002)
);

NOR4xp25_ASAP7_75t_SL g2003 ( 
.A(n_1961),
.B(n_258),
.C(n_256),
.D(n_257),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1960),
.Y(n_2004)
);

OAI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1944),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_2005)
);

XOR2xp5_ASAP7_75t_L g2006 ( 
.A(n_1904),
.B(n_260),
.Y(n_2006)
);

AO22x1_ASAP7_75t_L g2007 ( 
.A1(n_1908),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1861),
.A2(n_262),
.B(n_263),
.Y(n_2008)
);

AOI22xp5_ASAP7_75t_L g2009 ( 
.A1(n_1921),
.A2(n_266),
.B1(n_264),
.B2(n_265),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1850),
.B(n_265),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1910),
.B(n_266),
.Y(n_2011)
);

AOI222xp33_ASAP7_75t_L g2012 ( 
.A1(n_1937),
.A2(n_269),
.B1(n_271),
.B2(n_267),
.C1(n_268),
.C2(n_270),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1847),
.B(n_268),
.Y(n_2013)
);

AOI21xp5_ASAP7_75t_L g2014 ( 
.A1(n_1848),
.A2(n_269),
.B(n_272),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1911),
.A2(n_274),
.B1(n_272),
.B2(n_273),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1966),
.Y(n_2016)
);

AOI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1951),
.A2(n_273),
.B(n_274),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1941),
.B(n_275),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1854),
.Y(n_2019)
);

OAI21xp5_ASAP7_75t_SL g2020 ( 
.A1(n_1876),
.A2(n_276),
.B(n_277),
.Y(n_2020)
);

AOI222xp33_ASAP7_75t_L g2021 ( 
.A1(n_1914),
.A2(n_279),
.B1(n_278),
.B2(n_277),
.C1(n_280),
.C2(n_673),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1955),
.B(n_278),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1896),
.Y(n_2023)
);

OAI31xp33_ASAP7_75t_L g2024 ( 
.A1(n_1894),
.A2(n_279),
.A3(n_491),
.B(n_487),
.Y(n_2024)
);

INVx1_ASAP7_75t_SL g2025 ( 
.A(n_1945),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1947),
.B(n_492),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1930),
.B(n_1953),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1959),
.B(n_663),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_L g2029 ( 
.A(n_1969),
.B(n_497),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1932),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1881),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1878),
.Y(n_2032)
);

AND2x4_ASAP7_75t_SL g2033 ( 
.A(n_1880),
.B(n_498),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1879),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1963),
.Y(n_2035)
);

NAND2x1p5_ASAP7_75t_L g2036 ( 
.A(n_1963),
.B(n_501),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1883),
.Y(n_2037)
);

INVxp67_ASAP7_75t_SL g2038 ( 
.A(n_1901),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1963),
.B(n_514),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1889),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1890),
.Y(n_2041)
);

AOI32xp33_ASAP7_75t_L g2042 ( 
.A1(n_1905),
.A2(n_519),
.A3(n_515),
.B1(n_518),
.B2(n_520),
.Y(n_2042)
);

AOI21xp5_ASAP7_75t_L g2043 ( 
.A1(n_1923),
.A2(n_522),
.B(n_523),
.Y(n_2043)
);

NAND3xp33_ASAP7_75t_SL g2044 ( 
.A(n_1895),
.B(n_525),
.C(n_526),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1868),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1862),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1853),
.Y(n_2047)
);

OAI21xp5_ASAP7_75t_L g2048 ( 
.A1(n_1948),
.A2(n_528),
.B(n_532),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1936),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1938),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1893),
.B(n_537),
.Y(n_2051)
);

OAI21xp33_ASAP7_75t_SL g2052 ( 
.A1(n_1949),
.A2(n_538),
.B(n_539),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1950),
.Y(n_2053)
);

OAI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1898),
.A2(n_1920),
.B(n_1907),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1962),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_L g2056 ( 
.A1(n_1915),
.A2(n_545),
.B1(n_543),
.B2(n_544),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1916),
.A2(n_1954),
.B1(n_1965),
.B2(n_1952),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1885),
.B(n_546),
.Y(n_2058)
);

INVxp67_ASAP7_75t_SL g2059 ( 
.A(n_1902),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1992),
.B(n_1918),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_2035),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_2019),
.B(n_1863),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1975),
.Y(n_2063)
);

HB1xp67_ASAP7_75t_L g2064 ( 
.A(n_1985),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2025),
.B(n_1865),
.Y(n_2065)
);

INVx1_ASAP7_75t_SL g2066 ( 
.A(n_1988),
.Y(n_2066)
);

OR2x2_ASAP7_75t_L g2067 ( 
.A(n_2038),
.B(n_1884),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1982),
.Y(n_2068)
);

INVx2_ASAP7_75t_SL g2069 ( 
.A(n_1976),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_2057),
.B(n_1867),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_1973),
.A2(n_1995),
.B1(n_2027),
.B2(n_2020),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1983),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1984),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2059),
.B(n_1913),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_1993),
.B(n_1909),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1986),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_SL g2077 ( 
.A(n_1990),
.B(n_1891),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1991),
.B(n_1871),
.Y(n_2078)
);

INVxp67_ASAP7_75t_L g2079 ( 
.A(n_2054),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_2033),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1987),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_2014),
.B(n_1880),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1996),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2030),
.B(n_1857),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2047),
.B(n_1877),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2049),
.B(n_2050),
.Y(n_2086)
);

INVx1_ASAP7_75t_SL g2087 ( 
.A(n_2006),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1997),
.Y(n_2088)
);

NOR2x1p5_ASAP7_75t_SL g2089 ( 
.A(n_1972),
.B(n_1874),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_2000),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2053),
.B(n_1869),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2055),
.B(n_1882),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2002),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_1977),
.B(n_1849),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2004),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2046),
.B(n_1887),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1979),
.A2(n_1934),
.B1(n_1919),
.B2(n_1897),
.Y(n_2097)
);

INVx1_ASAP7_75t_SL g2098 ( 
.A(n_2039),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2045),
.B(n_1872),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2016),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_L g2101 ( 
.A(n_2013),
.B(n_1892),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2009),
.B(n_1888),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2040),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2005),
.B(n_1964),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_2036),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2015),
.A2(n_1942),
.B1(n_1971),
.B2(n_1926),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2041),
.B(n_1870),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2031),
.B(n_1968),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_2017),
.A2(n_1899),
.B1(n_1917),
.B2(n_1903),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2032),
.Y(n_2110)
);

AND2x4_ASAP7_75t_SL g2111 ( 
.A(n_2058),
.B(n_1928),
.Y(n_2111)
);

NAND2x1_ASAP7_75t_L g2112 ( 
.A(n_2023),
.B(n_2034),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1998),
.B(n_1970),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2010),
.B(n_1873),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2037),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2018),
.B(n_2022),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_2052),
.B(n_2024),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1974),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2064),
.Y(n_2119)
);

BUFx4f_ASAP7_75t_SL g2120 ( 
.A(n_2080),
.Y(n_2120)
);

CKINVDCx5p33_ASAP7_75t_R g2121 ( 
.A(n_2062),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2086),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2061),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_2075),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2118),
.Y(n_2125)
);

INVx3_ASAP7_75t_L g2126 ( 
.A(n_2111),
.Y(n_2126)
);

INVx5_ASAP7_75t_L g2127 ( 
.A(n_2105),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2063),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2068),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2087),
.B(n_2007),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_2072),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2073),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2066),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2070),
.B(n_2065),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_2112),
.Y(n_2135)
);

BUFx2_ASAP7_75t_L g2136 ( 
.A(n_2084),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2078),
.Y(n_2137)
);

INVxp33_ASAP7_75t_SL g2138 ( 
.A(n_2060),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2076),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2074),
.Y(n_2140)
);

INVx5_ASAP7_75t_L g2141 ( 
.A(n_2069),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2081),
.Y(n_2142)
);

INVxp33_ASAP7_75t_L g2143 ( 
.A(n_2077),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2116),
.Y(n_2144)
);

INVx2_ASAP7_75t_SL g2145 ( 
.A(n_2114),
.Y(n_2145)
);

CKINVDCx5p33_ASAP7_75t_R g2146 ( 
.A(n_2098),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2083),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2088),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2090),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_2093),
.Y(n_2150)
);

NAND3xp33_ASAP7_75t_L g2151 ( 
.A(n_2134),
.B(n_2079),
.C(n_2021),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2141),
.Y(n_2152)
);

O2A1O1Ixp33_ASAP7_75t_L g2153 ( 
.A1(n_2130),
.A2(n_2071),
.B(n_2082),
.C(n_2117),
.Y(n_2153)
);

NAND3xp33_ASAP7_75t_L g2154 ( 
.A(n_2127),
.B(n_2012),
.C(n_2008),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_SL g2155 ( 
.A(n_2121),
.B(n_2067),
.Y(n_2155)
);

AO21x1_ASAP7_75t_L g2156 ( 
.A1(n_2135),
.A2(n_1980),
.B(n_2011),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2119),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_2120),
.B(n_2102),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_2136),
.B(n_2089),
.Y(n_2159)
);

INVx2_ASAP7_75t_SL g2160 ( 
.A(n_2141),
.Y(n_2160)
);

AOI221xp5_ASAP7_75t_L g2161 ( 
.A1(n_2143),
.A2(n_2106),
.B1(n_1999),
.B2(n_2094),
.C(n_2110),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2126),
.B(n_2085),
.Y(n_2162)
);

NAND3xp33_ASAP7_75t_L g2163 ( 
.A(n_2127),
.B(n_2003),
.C(n_1994),
.Y(n_2163)
);

NAND4xp75_ASAP7_75t_L g2164 ( 
.A(n_2123),
.B(n_2048),
.C(n_2056),
.D(n_2043),
.Y(n_2164)
);

OAI211xp5_ASAP7_75t_SL g2165 ( 
.A1(n_2124),
.A2(n_2109),
.B(n_2097),
.C(n_2113),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2138),
.B(n_2104),
.Y(n_2166)
);

NAND3xp33_ASAP7_75t_SL g2167 ( 
.A(n_2146),
.B(n_2097),
.C(n_2042),
.Y(n_2167)
);

NOR3x1_ASAP7_75t_L g2168 ( 
.A(n_2145),
.B(n_2096),
.C(n_2091),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2160),
.B(n_2133),
.Y(n_2169)
);

NAND3xp33_ASAP7_75t_SL g2170 ( 
.A(n_2154),
.B(n_2140),
.C(n_2125),
.Y(n_2170)
);

NAND4xp25_ASAP7_75t_L g2171 ( 
.A(n_2151),
.B(n_2144),
.C(n_2137),
.D(n_2122),
.Y(n_2171)
);

NAND4xp25_ASAP7_75t_L g2172 ( 
.A(n_2153),
.B(n_2101),
.C(n_2129),
.D(n_2128),
.Y(n_2172)
);

AOI221xp5_ASAP7_75t_L g2173 ( 
.A1(n_2165),
.A2(n_2132),
.B1(n_2142),
.B2(n_2139),
.C(n_2131),
.Y(n_2173)
);

CKINVDCx20_ASAP7_75t_R g2174 ( 
.A(n_2158),
.Y(n_2174)
);

OAI221xp5_ASAP7_75t_L g2175 ( 
.A1(n_2163),
.A2(n_2161),
.B1(n_2159),
.B2(n_2155),
.C(n_2167),
.Y(n_2175)
);

AOI222xp33_ASAP7_75t_L g2176 ( 
.A1(n_2166),
.A2(n_2001),
.B1(n_1989),
.B2(n_2148),
.C1(n_2147),
.C2(n_2149),
.Y(n_2176)
);

BUFx2_ASAP7_75t_L g2177 ( 
.A(n_2152),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2177),
.Y(n_2178)
);

INVx3_ASAP7_75t_L g2179 ( 
.A(n_2169),
.Y(n_2179)
);

NAND2x1p5_ASAP7_75t_L g2180 ( 
.A(n_2174),
.B(n_2162),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_2171),
.B(n_2157),
.Y(n_2181)
);

NAND4xp75_ASAP7_75t_L g2182 ( 
.A(n_2173),
.B(n_2156),
.C(n_2168),
.D(n_2150),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2170),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2172),
.B(n_2099),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_SL g2185 ( 
.A(n_2175),
.B(n_2044),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2178),
.B(n_2176),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2180),
.B(n_2107),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_R g2188 ( 
.A(n_2179),
.B(n_1981),
.Y(n_2188)
);

NAND2xp33_ASAP7_75t_SL g2189 ( 
.A(n_2183),
.B(n_2092),
.Y(n_2189)
);

NAND2xp33_ASAP7_75t_SL g2190 ( 
.A(n_2184),
.B(n_1978),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_2187),
.B(n_2182),
.Y(n_2191)
);

NOR3xp33_ASAP7_75t_L g2192 ( 
.A(n_2186),
.B(n_2181),
.C(n_2029),
.Y(n_2192)
);

AOI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2191),
.A2(n_2190),
.B(n_2185),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2193),
.Y(n_2194)
);

OAI22xp5_ASAP7_75t_SL g2195 ( 
.A1(n_2194),
.A2(n_2189),
.B1(n_2192),
.B2(n_2188),
.Y(n_2195)
);

OR2x6_ASAP7_75t_L g2196 ( 
.A(n_2195),
.B(n_2108),
.Y(n_2196)
);

XOR2xp5_ASAP7_75t_L g2197 ( 
.A(n_2196),
.B(n_2164),
.Y(n_2197)
);

INVx4_ASAP7_75t_L g2198 ( 
.A(n_2197),
.Y(n_2198)
);

AOI221xp5_ASAP7_75t_L g2199 ( 
.A1(n_2198),
.A2(n_2095),
.B1(n_2100),
.B2(n_2115),
.C(n_2103),
.Y(n_2199)
);

AOI211xp5_ASAP7_75t_L g2200 ( 
.A1(n_2199),
.A2(n_2028),
.B(n_2026),
.C(n_2051),
.Y(n_2200)
);


endmodule