module fake_netlist_5_567_n_991 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_991);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_991;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_916;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_956;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_245;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_915;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_951;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_932;
wire n_417;
wire n_946;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_968;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_509;
wire n_568;
wire n_936;
wire n_373;
wire n_820;
wire n_947;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_905;
wire n_906;
wire n_406;
wire n_519;
wire n_470;
wire n_919;
wire n_782;
wire n_908;
wire n_325;
wire n_449;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_240;
wire n_942;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_920;
wire n_894;
wire n_271;
wire n_934;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_654;
wire n_370;
wire n_976;
wire n_234;
wire n_343;
wire n_379;
wire n_428;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_961;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_696;
wire n_255;
wire n_522;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_926;
wire n_344;
wire n_287;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_670;
wire n_486;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_974;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_903;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_966;
wire n_987;
wire n_253;
wire n_261;
wire n_289;
wire n_963;
wire n_745;
wire n_954;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_970;
wire n_911;
wire n_557;
wire n_354;
wire n_575;
wire n_607;
wire n_647;
wire n_480;
wire n_237;
wire n_425;
wire n_710;
wire n_407;
wire n_513;
wire n_707;
wire n_679;
wire n_527;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_656;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_937;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_536;
wire n_531;
wire n_935;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_960;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_904;
wire n_985;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_925;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_173),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_106),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_122),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_86),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_85),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_28),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_50),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_181),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_71),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_45),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_62),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_26),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_144),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_4),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_42),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_18),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_25),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_67),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_69),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_14),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_32),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_100),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_104),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_64),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_23),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_0),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_157),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_12),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g232 ( 
.A(n_110),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_97),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_59),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_4),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_21),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_52),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_148),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_105),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_163),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_135),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_137),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_125),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_51),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_190),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_30),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_79),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_121),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_150),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_94),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_32),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_24),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_162),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_156),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_119),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_49),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_151),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_149),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_27),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_66),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_108),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_23),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_61),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_113),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_155),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_48),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_81),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_172),
.Y(n_275)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_240),
.Y(n_276)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_195),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_260),
.B(n_0),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_228),
.B(n_1),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_232),
.Y(n_281)
);

CKINVDCx6p67_ASAP7_75t_R g282 ( 
.A(n_245),
.Y(n_282)
);

BUFx12f_ASAP7_75t_L g283 ( 
.A(n_194),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_206),
.B(n_222),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_240),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_223),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_206),
.B(n_2),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g289 ( 
.A(n_222),
.B(n_2),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_224),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_196),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_232),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

AND2x4_ASAP7_75t_L g294 ( 
.A(n_262),
.B(n_193),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_262),
.B(n_3),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_232),
.B(n_3),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_199),
.B(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_232),
.B(n_205),
.Y(n_299)
);

BUFx8_ASAP7_75t_L g300 ( 
.A(n_262),
.Y(n_300)
);

BUFx12f_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_232),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_207),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_218),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_232),
.B(n_5),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_250),
.B(n_6),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_209),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_210),
.B(n_6),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_212),
.B(n_192),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_213),
.B(n_7),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_219),
.B(n_7),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_197),
.Y(n_313)
);

AND2x4_ASAP7_75t_L g314 ( 
.A(n_226),
.B(n_191),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_234),
.B(n_41),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_238),
.B(n_8),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_8),
.Y(n_317)
);

AND2x4_ASAP7_75t_L g318 ( 
.A(n_247),
.B(n_43),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_198),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_255),
.B(n_9),
.Y(n_320)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_220),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_231),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_248),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_261),
.B(n_189),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_272),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_201),
.Y(n_327)
);

AND2x6_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_44),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_295),
.A2(n_235),
.B1(n_268),
.B2(n_236),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_274),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_280),
.A2(n_256),
.B1(n_202),
.B2(n_271),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_282),
.A2(n_237),
.B1(n_249),
.B2(n_265),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_288),
.A2(n_214),
.B1(n_203),
.B2(n_204),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_278),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_280),
.A2(n_254),
.B1(n_273),
.B2(n_271),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_254),
.B1(n_273),
.B2(n_270),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_244),
.B1(n_270),
.B2(n_200),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_208),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_309),
.A2(n_256),
.B1(n_244),
.B2(n_227),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_211),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_291),
.B(n_289),
.Y(n_343)
);

OR2x6_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_215),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_312),
.A2(n_275),
.B1(n_267),
.B2(n_266),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_278),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_263),
.B1(n_259),
.B2(n_258),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_305),
.B(n_217),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_297),
.A2(n_257),
.B1(n_253),
.B2(n_252),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_221),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_278),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_323),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_279),
.A2(n_251),
.B1(n_246),
.B2(n_243),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_L g356 ( 
.A1(n_316),
.A2(n_241),
.B1(n_239),
.B2(n_233),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_289),
.A2(n_307),
.B1(n_320),
.B2(n_317),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_321),
.A2(n_230),
.B1(n_225),
.B2(n_11),
.Y(n_358)
);

OAI22xp33_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_359)
);

CKINVDCx6p67_ASAP7_75t_R g360 ( 
.A(n_277),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_323),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_293),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_325),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_307),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_364)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_306),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_320),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_327),
.B(n_46),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_294),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_326),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_299),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_22),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_22),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_294),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g374 ( 
.A1(n_294),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_293),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_310),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_376)
);

AO22x2_ASAP7_75t_L g377 ( 
.A1(n_294),
.A2(n_324),
.B1(n_318),
.B2(n_315),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_301),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_301),
.A2(n_310),
.B1(n_314),
.B2(n_315),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_47),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_310),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_286),
.B(n_35),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_314),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_293),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_348),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_341),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g387 ( 
.A(n_354),
.Y(n_387)
);

OR2x6_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_374),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_346),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_336),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_369),
.B(n_331),
.Y(n_392)
);

OR2x6_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_283),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_283),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_363),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_360),
.B(n_283),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_319),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_319),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_349),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_335),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_353),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_375),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_384),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_L g410 ( 
.A(n_337),
.B(n_319),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_345),
.B(n_313),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_338),
.B(n_314),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_352),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_332),
.B(n_315),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_343),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g421 ( 
.A(n_372),
.B(n_37),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_380),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_345),
.B(n_286),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_357),
.B(n_315),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_357),
.B(n_347),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_374),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_383),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_R g429 ( 
.A(n_344),
.B(n_318),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_356),
.B(n_325),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_383),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_333),
.B(n_313),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_351),
.B(n_318),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_355),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_344),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_330),
.B(n_313),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_373),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_378),
.B(n_319),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_340),
.B(n_318),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_358),
.B(n_290),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_290),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_364),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_334),
.B(n_324),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_364),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_365),
.B(n_324),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_366),
.B(n_324),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_348),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_348),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_348),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_339),
.B(n_303),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_346),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_348),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_348),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_319),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_455),
.Y(n_460)
);

NAND2x1p5_ASAP7_75t_L g461 ( 
.A(n_425),
.B(n_281),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_395),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_392),
.A2(n_402),
.B(n_398),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_425),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_395),
.B(n_319),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_412),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_403),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_418),
.B(n_300),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_403),
.Y(n_469)
);

NAND2x1p5_ASAP7_75t_L g470 ( 
.A(n_430),
.B(n_281),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_424),
.B(n_300),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_426),
.A2(n_328),
.B(n_281),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_386),
.B(n_416),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_386),
.B(n_325),
.Y(n_475)
);

BUFx12f_ASAP7_75t_SL g476 ( 
.A(n_393),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_440),
.B(n_303),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_R g478 ( 
.A(n_435),
.B(n_429),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_426),
.B(n_328),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_389),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_396),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_53),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_440),
.B(n_447),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_328),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

BUFx5_ASAP7_75t_L g486 ( 
.A(n_407),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_433),
.B(n_287),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_287),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_448),
.B(n_287),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_442),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_438),
.B(n_292),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_443),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_452),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_445),
.B(n_328),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_427),
.B(n_292),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_388),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_292),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_445),
.A2(n_328),
.B(n_302),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_450),
.B(n_328),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_453),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_450),
.B(n_328),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_405),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_428),
.B(n_302),
.Y(n_504)
);

NAND2x1p5_ASAP7_75t_L g505 ( 
.A(n_431),
.B(n_302),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_457),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_458),
.B(n_304),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_388),
.B(n_54),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_304),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_388),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_394),
.B(n_302),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_409),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_449),
.B(n_304),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_304),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_R g518 ( 
.A(n_414),
.B(n_304),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g519 ( 
.A(n_421),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_393),
.B(n_304),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_456),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_387),
.B(n_308),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_393),
.B(n_308),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_399),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_410),
.B(n_300),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_413),
.B(n_308),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_400),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_413),
.B(n_308),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_439),
.B(n_55),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_401),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_56),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_404),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_434),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_399),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_406),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_387),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_387),
.Y(n_537)
);

BUFx2_ASAP7_75t_SL g538 ( 
.A(n_387),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_437),
.B(n_57),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_419),
.B(n_308),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_460),
.B(n_391),
.Y(n_541)
);

BUFx12f_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_488),
.B(n_415),
.Y(n_543)
);

NAND2x1p5_ASAP7_75t_L g544 ( 
.A(n_462),
.B(n_432),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_515),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_488),
.B(n_308),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_489),
.B(n_444),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_466),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_466),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_462),
.B(n_444),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_467),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_498),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_467),
.Y(n_554)
);

AND2x6_ASAP7_75t_L g555 ( 
.A(n_509),
.B(n_429),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_464),
.B(n_436),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_464),
.B(n_436),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_460),
.B(n_397),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

NOR2x1_ASAP7_75t_SL g560 ( 
.A(n_538),
.B(n_276),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_474),
.B(n_38),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_474),
.B(n_39),
.Y(n_562)
);

INVx5_ASAP7_75t_L g563 ( 
.A(n_495),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_515),
.B(n_39),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_493),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_469),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_489),
.B(n_293),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_493),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_510),
.B(n_293),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_506),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_506),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_509),
.B(n_58),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_496),
.B(n_60),
.Y(n_573)
);

NAND2x1p5_ASAP7_75t_L g574 ( 
.A(n_510),
.B(n_293),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_496),
.B(n_63),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_507),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_490),
.B(n_40),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_507),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_498),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_535),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_529),
.B(n_296),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_475),
.B(n_296),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_475),
.B(n_296),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_511),
.Y(n_584)
);

BUFx5_ASAP7_75t_L g585 ( 
.A(n_495),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_535),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_524),
.B(n_40),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_526),
.B(n_296),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_498),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_526),
.B(n_296),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_491),
.B(n_65),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_491),
.B(n_68),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_SL g593 ( 
.A(n_479),
.B(n_300),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_492),
.B(n_70),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_514),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_514),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_497),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_477),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_472),
.Y(n_599)
);

INVx6_ASAP7_75t_L g600 ( 
.A(n_529),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_477),
.B(n_296),
.Y(n_601)
);

NAND2x2_ASAP7_75t_L g602 ( 
.A(n_476),
.B(n_478),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_497),
.B(n_517),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_520),
.B(n_73),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_498),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_517),
.B(n_302),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_552),
.Y(n_607)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_553),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_587),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_542),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_547),
.A2(n_479),
.B1(n_539),
.B2(n_531),
.Y(n_612)
);

BUFx4_ASAP7_75t_SL g613 ( 
.A(n_584),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_461),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_565),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_545),
.Y(n_616)
);

INVxp67_ASAP7_75t_SL g617 ( 
.A(n_603),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_554),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_556),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_563),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_545),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_556),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_557),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_579),
.Y(n_625)
);

BUFx2_ASAP7_75t_SL g626 ( 
.A(n_551),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_579),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_598),
.B(n_483),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_568),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_557),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_550),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_547),
.B(n_540),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

BUFx2_ASAP7_75t_SL g634 ( 
.A(n_551),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_579),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_563),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_541),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_589),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_570),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_589),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_572),
.Y(n_641)
);

CKINVDCx14_ASAP7_75t_R g642 ( 
.A(n_555),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_589),
.Y(n_643)
);

BUFx5_ASAP7_75t_L g644 ( 
.A(n_591),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_543),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_598),
.B(n_483),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_543),
.B(n_540),
.Y(n_647)
);

INVx1_ASAP7_75t_SL g648 ( 
.A(n_564),
.Y(n_648)
);

BUFx6f_ASAP7_75t_SL g649 ( 
.A(n_555),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

NAND2x1p5_ASAP7_75t_L g651 ( 
.A(n_563),
.B(n_529),
.Y(n_651)
);

NAND2x1p5_ASAP7_75t_L g652 ( 
.A(n_563),
.B(n_466),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_605),
.Y(n_653)
);

INVx8_ASAP7_75t_L g654 ( 
.A(n_555),
.Y(n_654)
);

BUFx12f_ASAP7_75t_L g655 ( 
.A(n_544),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_605),
.Y(n_657)
);

NAND2x1p5_ASAP7_75t_L g658 ( 
.A(n_605),
.B(n_466),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_600),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_604),
.B(n_472),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_600),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_604),
.B(n_573),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_576),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_559),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_575),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_597),
.B(n_516),
.Y(n_666)
);

NAND2x1p5_ASAP7_75t_L g667 ( 
.A(n_591),
.B(n_466),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_616),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_612),
.A2(n_600),
.B1(n_597),
.B2(n_603),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_662),
.A2(n_528),
.B1(n_578),
.B2(n_544),
.Y(n_670)
);

INVx1_ASAP7_75t_SL g671 ( 
.A(n_613),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_616),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_607),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_611),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_615),
.Y(n_675)
);

INVx1_ASAP7_75t_SL g676 ( 
.A(n_622),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_622),
.Y(n_677)
);

INVx6_ASAP7_75t_L g678 ( 
.A(n_661),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_662),
.Y(n_679)
);

CKINVDCx11_ASAP7_75t_R g680 ( 
.A(n_610),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_655),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_607),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_629),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_647),
.A2(n_531),
.B1(n_539),
.B2(n_555),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_645),
.A2(n_558),
.B1(n_539),
.B2(n_531),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_645),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_619),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_SL g688 ( 
.A1(n_637),
.A2(n_533),
.B1(n_534),
.B2(n_577),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_639),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_637),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g691 ( 
.A1(n_647),
.A2(n_592),
.B1(n_602),
.B2(n_561),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_632),
.A2(n_592),
.B1(n_562),
.B2(n_575),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_650),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_611),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_663),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_626),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_632),
.A2(n_471),
.B1(n_463),
.B2(n_594),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_619),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_662),
.A2(n_495),
.B1(n_468),
.B2(n_520),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_660),
.A2(n_595),
.B1(n_596),
.B2(n_580),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_664),
.Y(n_701)
);

BUFx2_ASAP7_75t_SL g702 ( 
.A(n_610),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_664),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_660),
.A2(n_586),
.B1(n_461),
.B2(n_470),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_611),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_628),
.Y(n_706)
);

CKINVDCx11_ASAP7_75t_R g707 ( 
.A(n_623),
.Y(n_707)
);

INVx6_ASAP7_75t_L g708 ( 
.A(n_661),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_617),
.B(n_516),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_666),
.B(n_487),
.Y(n_710)
);

BUFx10_ASAP7_75t_L g711 ( 
.A(n_649),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_634),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_646),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_666),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_655),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_648),
.B(n_487),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_SL g717 ( 
.A1(n_624),
.A2(n_519),
.B1(n_504),
.B2(n_505),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_620),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_660),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_641),
.A2(n_495),
.B1(n_523),
.B2(n_599),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_656),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_630),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_681),
.B(n_631),
.Y(n_723)
);

OAI21xp33_ASAP7_75t_L g724 ( 
.A1(n_697),
.A2(n_609),
.B(n_656),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_710),
.B(n_523),
.Y(n_725)
);

INVxp67_ASAP7_75t_SL g726 ( 
.A(n_709),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_674),
.Y(n_727)
);

BUFx12f_ASAP7_75t_L g728 ( 
.A(n_680),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_675),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_692),
.A2(n_665),
.B1(n_641),
.B2(n_614),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_L g731 ( 
.A1(n_685),
.A2(n_706),
.B1(n_713),
.B2(n_684),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_683),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_691),
.A2(n_644),
.B1(n_642),
.B2(n_649),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_710),
.A2(n_593),
.B1(n_473),
.B2(n_665),
.Y(n_734)
);

OAI22xp33_ASAP7_75t_L g735 ( 
.A1(n_696),
.A2(n_593),
.B1(n_614),
.B2(n_633),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_714),
.A2(n_649),
.B1(n_642),
.B2(n_644),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_676),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_669),
.A2(n_644),
.B1(n_501),
.B2(n_480),
.Y(n_738)
);

BUFx4f_ASAP7_75t_SL g739 ( 
.A(n_671),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_717),
.A2(n_644),
.B1(n_501),
.B2(n_480),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_688),
.A2(n_614),
.B1(n_667),
.B2(n_631),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_696),
.A2(n_614),
.B1(n_667),
.B2(n_633),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_718),
.A2(n_644),
.B1(n_566),
.B2(n_654),
.Y(n_743)
);

INVx5_ASAP7_75t_SL g744 ( 
.A(n_674),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_712),
.A2(n_651),
.B1(n_661),
.B2(n_659),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_689),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_718),
.A2(n_722),
.B1(n_707),
.B2(n_695),
.Y(n_747)
);

BUFx12f_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_722),
.B(n_481),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_707),
.A2(n_644),
.B1(n_654),
.B2(n_499),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_677),
.Y(n_751)
);

OAI22xp5_ASAP7_75t_L g752 ( 
.A1(n_712),
.A2(n_651),
.B1(n_661),
.B2(n_659),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_699),
.A2(n_661),
.B1(n_659),
.B2(n_581),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_686),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_673),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_693),
.A2(n_716),
.B1(n_686),
.B2(n_719),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_670),
.A2(n_703),
.B1(n_690),
.B2(n_644),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_673),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_682),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_672),
.B(n_495),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_690),
.A2(n_581),
.B1(n_504),
.B2(n_505),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_702),
.Y(n_762)
);

AOI211xp5_ASAP7_75t_L g763 ( 
.A1(n_721),
.A2(n_525),
.B(n_482),
.C(n_494),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_700),
.A2(n_654),
.B1(n_470),
.B2(n_601),
.Y(n_764)
);

INVx5_ASAP7_75t_SL g765 ( 
.A(n_674),
.Y(n_765)
);

OAI21xp33_ASAP7_75t_L g766 ( 
.A1(n_720),
.A2(n_459),
.B(n_512),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_668),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_682),
.Y(n_768)
);

BUFx8_ASAP7_75t_SL g769 ( 
.A(n_668),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_687),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_672),
.B(n_618),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_687),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_SL g773 ( 
.A1(n_681),
.A2(n_654),
.B1(n_470),
.B2(n_500),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_715),
.A2(n_502),
.B1(n_636),
.B2(n_621),
.Y(n_774)
);

OAI21xp33_ASAP7_75t_L g775 ( 
.A1(n_715),
.A2(n_601),
.B(n_484),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_698),
.A2(n_546),
.B1(n_582),
.B2(n_583),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_698),
.B(n_618),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_701),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_678),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_701),
.A2(n_546),
.B1(n_582),
.B2(n_583),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_SL g781 ( 
.A1(n_704),
.A2(n_513),
.B(n_461),
.Y(n_781)
);

AOI222xp33_ASAP7_75t_L g782 ( 
.A1(n_679),
.A2(n_495),
.B1(n_569),
.B2(n_567),
.C1(n_532),
.C2(n_530),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_SL g783 ( 
.A1(n_674),
.A2(n_513),
.B(n_476),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_726),
.B(n_711),
.Y(n_784)
);

AO22x1_ASAP7_75t_L g785 ( 
.A1(n_741),
.A2(n_711),
.B1(n_705),
.B2(n_694),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_755),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_724),
.A2(n_711),
.B1(n_679),
.B2(n_532),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_731),
.A2(n_679),
.B1(n_708),
.B2(n_678),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_SL g789 ( 
.A1(n_730),
.A2(n_708),
.B1(n_678),
.B2(n_513),
.Y(n_789)
);

OAI222xp33_ASAP7_75t_L g790 ( 
.A1(n_740),
.A2(n_504),
.B1(n_505),
.B2(n_574),
.C1(n_569),
.C2(n_588),
.Y(n_790)
);

OAI222xp33_ASAP7_75t_L g791 ( 
.A1(n_740),
.A2(n_574),
.B1(n_590),
.B2(n_588),
.C1(n_638),
.C2(n_640),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_731),
.A2(n_530),
.B1(n_465),
.B2(n_498),
.Y(n_792)
);

AOI222xp33_ASAP7_75t_L g793 ( 
.A1(n_725),
.A2(n_590),
.B1(n_567),
.B2(n_302),
.C1(n_606),
.C2(n_508),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_756),
.A2(n_708),
.B1(n_678),
.B2(n_606),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_SL g795 ( 
.A1(n_754),
.A2(n_708),
.B1(n_636),
.B2(n_621),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_747),
.A2(n_636),
.B1(n_621),
.B2(n_640),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_781),
.A2(n_763),
.B(n_750),
.Y(n_797)
);

AND2x2_ASAP7_75t_SL g798 ( 
.A(n_750),
.B(n_608),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_L g799 ( 
.A1(n_733),
.A2(n_527),
.B1(n_618),
.B2(n_643),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_756),
.B(n_749),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_SL g801 ( 
.A1(n_757),
.A2(n_635),
.B(n_643),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_737),
.B(n_694),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_751),
.B(n_694),
.Y(n_803)
);

OA21x2_ASAP7_75t_L g804 ( 
.A1(n_775),
.A2(n_522),
.B(n_638),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_747),
.A2(n_527),
.B1(n_635),
.B2(n_643),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_729),
.B(n_694),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_757),
.A2(n_735),
.B1(n_766),
.B2(n_736),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_736),
.A2(n_743),
.B1(n_734),
.B2(n_762),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_761),
.A2(n_738),
.B1(n_734),
.B2(n_748),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_738),
.A2(n_527),
.B1(n_635),
.B2(n_503),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_770),
.Y(n_811)
);

AOI221xp5_ASAP7_75t_L g812 ( 
.A1(n_732),
.A2(n_485),
.B1(n_503),
.B2(n_527),
.C(n_521),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_728),
.A2(n_527),
.B1(n_485),
.B2(n_503),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_773),
.A2(n_485),
.B1(n_585),
.B2(n_548),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_755),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_782),
.A2(n_585),
.B1(n_548),
.B2(n_549),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_758),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_743),
.A2(n_585),
.B1(n_549),
.B2(n_705),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_723),
.A2(n_621),
.B1(n_636),
.B2(n_608),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_783),
.B(n_608),
.C(n_705),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_746),
.B(n_705),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_767),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_742),
.A2(n_585),
.B1(n_521),
.B2(n_653),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_758),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_764),
.A2(n_621),
.B1(n_636),
.B2(n_652),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_764),
.A2(n_652),
.B1(n_658),
.B2(n_653),
.Y(n_826)
);

AOI22xp33_ASAP7_75t_L g827 ( 
.A1(n_779),
.A2(n_585),
.B1(n_521),
.B2(n_653),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_779),
.A2(n_521),
.B1(n_657),
.B2(n_653),
.Y(n_828)
);

OAI211xp5_ASAP7_75t_SL g829 ( 
.A1(n_774),
.A2(n_537),
.B(n_518),
.C(n_536),
.Y(n_829)
);

OAI21xp5_ASAP7_75t_SL g830 ( 
.A1(n_745),
.A2(n_752),
.B(n_753),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_776),
.A2(n_611),
.B1(n_657),
.B2(n_627),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_768),
.B(n_625),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_777),
.B(n_625),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_760),
.A2(n_521),
.B1(n_657),
.B2(n_627),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_771),
.A2(n_657),
.B1(n_627),
.B2(n_625),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_811),
.B(n_768),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_811),
.B(n_778),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_784),
.B(n_759),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_808),
.B(n_772),
.C(n_769),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_809),
.A2(n_739),
.B1(n_776),
.B2(n_780),
.Y(n_840)
);

OAI22x1_ASAP7_75t_L g841 ( 
.A1(n_788),
.A2(n_765),
.B1(n_744),
.B2(n_658),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_822),
.B(n_780),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_786),
.B(n_815),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_800),
.B(n_727),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_807),
.A2(n_765),
.B1(n_744),
.B2(n_727),
.Y(n_845)
);

OAI221xp5_ASAP7_75t_L g846 ( 
.A1(n_797),
.A2(n_727),
.B1(n_627),
.B2(n_625),
.C(n_77),
.Y(n_846)
);

OAI221xp5_ASAP7_75t_L g847 ( 
.A1(n_787),
.A2(n_727),
.B1(n_75),
.B2(n_76),
.C(n_78),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_788),
.A2(n_765),
.B1(n_744),
.B2(n_486),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_786),
.B(n_74),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_792),
.B(n_285),
.C(n_276),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_SL g851 ( 
.A1(n_830),
.A2(n_80),
.B(n_82),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_L g852 ( 
.A(n_793),
.B(n_285),
.C(n_276),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_805),
.B(n_285),
.C(n_276),
.Y(n_853)
);

OA21x2_ASAP7_75t_L g854 ( 
.A1(n_831),
.A2(n_536),
.B(n_560),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_819),
.B(n_820),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_806),
.B(n_83),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_821),
.B(n_87),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_L g858 ( 
.A1(n_796),
.A2(n_285),
.B1(n_276),
.B2(n_538),
.C(n_91),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_802),
.B(n_88),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_803),
.B(n_89),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_815),
.B(n_90),
.Y(n_861)
);

OAI221xp5_ASAP7_75t_SL g862 ( 
.A1(n_801),
.A2(n_794),
.B1(n_799),
.B2(n_816),
.C(n_831),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_817),
.B(n_92),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_L g864 ( 
.A(n_794),
.B(n_285),
.C(n_276),
.Y(n_864)
);

OAI221xp5_ASAP7_75t_L g865 ( 
.A1(n_789),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.C(n_98),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_817),
.B(n_101),
.Y(n_866)
);

AOI221xp5_ASAP7_75t_SL g867 ( 
.A1(n_825),
.A2(n_102),
.B1(n_103),
.B2(n_107),
.C(n_109),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_824),
.B(n_111),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_824),
.B(n_112),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_833),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_SL g871 ( 
.A1(n_795),
.A2(n_114),
.B(n_115),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_832),
.B(n_116),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_L g873 ( 
.A1(n_820),
.A2(n_813),
.B1(n_798),
.B2(n_823),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_832),
.B(n_117),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_804),
.B(n_118),
.Y(n_875)
);

NOR3xp33_ASAP7_75t_L g876 ( 
.A(n_851),
.B(n_846),
.C(n_865),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_L g877 ( 
.A(n_847),
.B(n_785),
.C(n_829),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_870),
.B(n_785),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_839),
.A2(n_798),
.B1(n_814),
.B2(n_818),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_844),
.B(n_804),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_838),
.B(n_791),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_842),
.B(n_804),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_862),
.A2(n_835),
.B1(n_834),
.B2(n_828),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_837),
.B(n_826),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_867),
.B(n_855),
.C(n_858),
.Y(n_885)
);

NAND4xp75_ASAP7_75t_L g886 ( 
.A(n_875),
.B(n_812),
.C(n_790),
.D(n_124),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_843),
.B(n_810),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_SL g888 ( 
.A(n_840),
.B(n_827),
.C(n_123),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_871),
.B(n_537),
.C(n_127),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_SL g890 ( 
.A(n_845),
.B(n_873),
.C(n_872),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_837),
.B(n_120),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_L g892 ( 
.A(n_856),
.B(n_285),
.C(n_129),
.Y(n_892)
);

NAND4xp75_ASAP7_75t_L g893 ( 
.A(n_875),
.B(n_128),
.C(n_130),
.D(n_131),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_843),
.B(n_132),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_852),
.A2(n_136),
.B(n_138),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_836),
.B(n_139),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_L g897 ( 
.A(n_857),
.B(n_860),
.C(n_859),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_836),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_864),
.B(n_537),
.C(n_142),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_898),
.B(n_841),
.Y(n_900)
);

NOR3xp33_ASAP7_75t_SL g901 ( 
.A(n_885),
.B(n_864),
.C(n_853),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_880),
.B(n_841),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_882),
.Y(n_903)
);

NAND4xp75_ASAP7_75t_L g904 ( 
.A(n_890),
.B(n_874),
.C(n_869),
.D(n_849),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_878),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_881),
.B(n_869),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_884),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_887),
.B(n_854),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_897),
.B(n_894),
.Y(n_909)
);

XNOR2x2_ASAP7_75t_L g910 ( 
.A(n_886),
.B(n_853),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_891),
.B(n_854),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_896),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_877),
.B(n_854),
.Y(n_913)
);

XOR2xp5_ASAP7_75t_L g914 ( 
.A(n_888),
.B(n_874),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_877),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_879),
.B(n_854),
.Y(n_916)
);

NOR3xp33_ASAP7_75t_L g917 ( 
.A(n_876),
.B(n_868),
.C(n_863),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_905),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_905),
.Y(n_919)
);

XOR2x2_ASAP7_75t_L g920 ( 
.A(n_904),
.B(n_889),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_900),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_907),
.B(n_899),
.Y(n_922)
);

AO22x2_ASAP7_75t_L g923 ( 
.A1(n_913),
.A2(n_893),
.B1(n_883),
.B2(n_888),
.Y(n_923)
);

XNOR2x1_ASAP7_75t_L g924 ( 
.A(n_915),
.B(n_895),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_909),
.B(n_906),
.Y(n_925)
);

INVxp67_ASAP7_75t_L g926 ( 
.A(n_913),
.Y(n_926)
);

OA22x2_ASAP7_75t_L g927 ( 
.A1(n_914),
.A2(n_866),
.B1(n_849),
.B2(n_861),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_919),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_921),
.Y(n_929)
);

INVxp33_ASAP7_75t_L g930 ( 
.A(n_925),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_918),
.Y(n_931)
);

AOI22x1_ASAP7_75t_L g932 ( 
.A1(n_923),
.A2(n_914),
.B1(n_916),
.B2(n_910),
.Y(n_932)
);

OAI22x1_ASAP7_75t_L g933 ( 
.A1(n_926),
.A2(n_907),
.B1(n_900),
.B2(n_902),
.Y(n_933)
);

OA22x2_ASAP7_75t_L g934 ( 
.A1(n_926),
.A2(n_902),
.B1(n_916),
.B2(n_912),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_922),
.B(n_903),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_923),
.A2(n_917),
.B1(n_904),
.B2(n_901),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_931),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_928),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_929),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_935),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_932),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_934),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_938),
.B(n_930),
.Y(n_943)
);

AOI221xp5_ASAP7_75t_L g944 ( 
.A1(n_941),
.A2(n_936),
.B1(n_933),
.B2(n_932),
.C(n_922),
.Y(n_944)
);

OA22x2_ASAP7_75t_L g945 ( 
.A1(n_941),
.A2(n_920),
.B1(n_924),
.B2(n_908),
.Y(n_945)
);

INVxp67_ASAP7_75t_L g946 ( 
.A(n_942),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_946),
.Y(n_947)
);

AOI221xp5_ASAP7_75t_L g948 ( 
.A1(n_944),
.A2(n_940),
.B1(n_937),
.B2(n_939),
.C(n_908),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_943),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_945),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_948),
.A2(n_927),
.B1(n_911),
.B2(n_892),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_950),
.A2(n_947),
.B1(n_949),
.B2(n_927),
.Y(n_952)
);

AO22x1_ASAP7_75t_L g953 ( 
.A1(n_950),
.A2(n_910),
.B1(n_866),
.B2(n_911),
.Y(n_953)
);

AOI31xp33_ASAP7_75t_L g954 ( 
.A1(n_950),
.A2(n_850),
.A3(n_848),
.B(n_145),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_948),
.A2(n_850),
.B1(n_486),
.B2(n_146),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_950),
.B(n_140),
.Y(n_956)
);

NOR2x2_ASAP7_75t_L g957 ( 
.A(n_953),
.B(n_143),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_956),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_952),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_954),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_951),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_955),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_958),
.Y(n_963)
);

AND3x1_ASAP7_75t_L g964 ( 
.A(n_959),
.B(n_147),
.C(n_152),
.Y(n_964)
);

AND4x1_ASAP7_75t_L g965 ( 
.A(n_960),
.B(n_153),
.C(n_154),
.D(n_158),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_957),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_961),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_967),
.B(n_957),
.C(n_962),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_966),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_966),
.Y(n_970)
);

BUFx8_ASAP7_75t_L g971 ( 
.A(n_963),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_964),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_972),
.A2(n_965),
.B1(n_486),
.B2(n_161),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_969),
.Y(n_974)
);

AOI22xp5_ASAP7_75t_L g975 ( 
.A1(n_970),
.A2(n_486),
.B1(n_160),
.B2(n_164),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_971),
.Y(n_976)
);

AO22x2_ASAP7_75t_L g977 ( 
.A1(n_968),
.A2(n_159),
.B1(n_165),
.B2(n_166),
.Y(n_977)
);

INVxp67_ASAP7_75t_SL g978 ( 
.A(n_976),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_974),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_977),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_978),
.A2(n_973),
.B1(n_975),
.B2(n_486),
.Y(n_981)
);

OAI22xp33_ASAP7_75t_L g982 ( 
.A1(n_980),
.A2(n_167),
.B1(n_169),
.B2(n_170),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_981),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_982),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_984),
.A2(n_979),
.B1(n_486),
.B2(n_175),
.Y(n_985)
);

AOI22xp33_ASAP7_75t_L g986 ( 
.A1(n_983),
.A2(n_486),
.B1(n_174),
.B2(n_176),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_984),
.A2(n_486),
.B1(n_177),
.B2(n_178),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_985),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_987),
.Y(n_989)
);

AOI221xp5_ASAP7_75t_L g990 ( 
.A1(n_989),
.A2(n_986),
.B1(n_180),
.B2(n_182),
.C(n_183),
.Y(n_990)
);

AOI211xp5_ASAP7_75t_L g991 ( 
.A1(n_990),
.A2(n_988),
.B(n_184),
.C(n_185),
.Y(n_991)
);


endmodule