module fake_jpeg_2452_n_168 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_23),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_66),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_49),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_61),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_46),
.B1(n_55),
.B2(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_75),
.B1(n_76),
.B2(n_45),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_46),
.B1(n_45),
.B2(n_52),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_63),
.A2(n_60),
.B1(n_57),
.B2(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_71),
.A2(n_50),
.A3(n_47),
.B1(n_58),
.B2(n_60),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_88),
.B(n_68),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_84),
.B1(n_88),
.B2(n_83),
.Y(n_109)
);

NAND2xp33_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_61),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_86),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_20),
.C(n_40),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_48),
.B(n_54),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_0),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_78),
.B1(n_79),
.B2(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_7),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_43),
.C(n_42),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_85),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_41),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_118),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_100),
.A2(n_92),
.B(n_5),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_127),
.B(n_128),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_104),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_122),
.C(n_123),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_39),
.B(n_38),
.C(n_37),
.Y(n_121)
);

NAND4xp25_ASAP7_75t_SL g137 ( 
.A(n_121),
.B(n_125),
.C(n_21),
.D(n_31),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_6),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_126),
.B1(n_12),
.B2(n_13),
.Y(n_141)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_102),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_99),
.B1(n_101),
.B2(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_7),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_27),
.B(n_26),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_36),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_12),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_136),
.B1(n_141),
.B2(n_124),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_35),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_139),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_135),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_130),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_113),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_145),
.C(n_25),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_34),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_142),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_134),
.A2(n_116),
.B(n_115),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_140),
.C(n_143),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_156),
.C(n_157),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_138),
.C(n_144),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_153),
.B(n_138),
.C(n_144),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_137),
.B1(n_125),
.B2(n_129),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_125),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_149),
.B(n_150),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_161),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_24),
.C(n_14),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_162),
.C(n_14),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_13),
.C(n_15),
.Y(n_166)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_166),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_17),
.Y(n_168)
);


endmodule