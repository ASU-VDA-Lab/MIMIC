module fake_jpeg_1432_n_122 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_16),
.B(n_27),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_60),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_40),
.B1(n_38),
.B2(n_42),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_62),
.B1(n_40),
.B2(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_34),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_36),
.B1(n_43),
.B2(n_41),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_59),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_40),
.C(n_46),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_14),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_67),
.B(n_58),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_50),
.B1(n_46),
.B2(n_51),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_74),
.B1(n_58),
.B2(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_73),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_49),
.B1(n_39),
.B2(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_78),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_74),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_2),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_86),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_71),
.B1(n_18),
.B2(n_19),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_90),
.B(n_7),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_3),
.B(n_4),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_95),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_4),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.C(n_8),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_6),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_100),
.B(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_9),
.Y(n_113)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_88),
.C(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_109),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_108),
.C(n_110),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_8),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_22),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_9),
.B(n_10),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_113),
.B(n_104),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_116),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g116 ( 
.A(n_112),
.B(n_105),
.Y(n_116)
);

OAI31xp33_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_111),
.A3(n_114),
.B(n_107),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_12),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_20),
.B(n_26),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_28),
.C(n_29),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_30),
.Y(n_122)
);


endmodule