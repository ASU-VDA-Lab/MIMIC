module real_aes_1754_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_0), .B(n_130), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_1), .A2(n_124), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_2), .B(n_801), .Y(n_800) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_3), .B(n_141), .Y(n_216) );
INVx1_ASAP7_75t_L g129 ( .A(n_4), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_5), .B(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_6), .B(n_193), .Y(n_490) );
INVx1_ASAP7_75t_L g533 ( .A(n_7), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g801 ( .A(n_8), .Y(n_801) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_9), .Y(n_547) );
NAND2xp33_ASAP7_75t_L g192 ( .A(n_10), .B(n_139), .Y(n_192) );
INVx2_ASAP7_75t_L g121 ( .A(n_11), .Y(n_121) );
AOI221x1_ASAP7_75t_L g123 ( .A1(n_12), .A2(n_25), .B1(n_124), .B2(n_130), .C(n_137), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_13), .Y(n_418) );
AND3x1_ASAP7_75t_L g798 ( .A(n_13), .B(n_41), .C(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_14), .B(n_130), .Y(n_188) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_15), .A2(n_186), .B(n_187), .Y(n_185) );
INVx1_ASAP7_75t_L g499 ( .A(n_16), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_17), .B(n_119), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_18), .B(n_141), .Y(n_200) );
AO21x1_ASAP7_75t_L g211 ( .A1(n_19), .A2(n_130), .B(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_20), .Y(n_784) );
INVx1_ASAP7_75t_L g422 ( .A(n_21), .Y(n_422) );
NOR2xp33_ASAP7_75t_SL g796 ( .A(n_21), .B(n_423), .Y(n_796) );
INVx1_ASAP7_75t_L g497 ( .A(n_22), .Y(n_497) );
INVx1_ASAP7_75t_SL g483 ( .A(n_23), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_24), .B(n_131), .Y(n_461) );
NAND2x1_ASAP7_75t_L g149 ( .A(n_26), .B(n_141), .Y(n_149) );
AOI33xp33_ASAP7_75t_L g514 ( .A1(n_27), .A2(n_56), .A3(n_449), .B1(n_458), .B2(n_515), .B3(n_516), .Y(n_514) );
NAND2x1_ASAP7_75t_L g179 ( .A(n_28), .B(n_139), .Y(n_179) );
INVx1_ASAP7_75t_L g541 ( .A(n_29), .Y(n_541) );
OR2x2_ASAP7_75t_L g122 ( .A(n_30), .B(n_88), .Y(n_122) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_30), .A2(n_88), .B(n_121), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_31), .B(n_474), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_32), .B(n_139), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g771 ( .A1(n_33), .A2(n_34), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_33), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_34), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_35), .B(n_141), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_36), .A2(n_37), .B1(n_108), .B2(n_109), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_36), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_37), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_38), .B(n_139), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_39), .A2(n_124), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g125 ( .A(n_40), .B(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g136 ( .A(n_40), .B(n_129), .Y(n_136) );
INVx1_ASAP7_75t_L g457 ( .A(n_40), .Y(n_457) );
OR2x6_ASAP7_75t_L g420 ( .A(n_41), .B(n_421), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_42), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_43), .B(n_130), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_44), .B(n_474), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_45), .A2(n_154), .B1(n_193), .B2(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_46), .B(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_47), .B(n_131), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_48), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_49), .B(n_139), .Y(n_161) );
INVxp33_ASAP7_75t_L g803 ( .A(n_50), .Y(n_803) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_51), .B(n_186), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_52), .B(n_131), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_53), .A2(n_124), .B(n_178), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_54), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_55), .B(n_139), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_57), .B(n_131), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_58), .Y(n_425) );
INVx1_ASAP7_75t_L g128 ( .A(n_59), .Y(n_128) );
INVx1_ASAP7_75t_L g133 ( .A(n_59), .Y(n_133) );
AND2x2_ASAP7_75t_L g526 ( .A(n_60), .B(n_119), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g531 ( .A1(n_61), .A2(n_77), .B1(n_455), .B2(n_474), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_62), .B(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_63), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_64), .B(n_154), .Y(n_549) );
AOI21xp5_ASAP7_75t_SL g469 ( .A1(n_65), .A2(n_455), .B(n_470), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_66), .A2(n_124), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g493 ( .A(n_67), .Y(n_493) );
AO21x1_ASAP7_75t_L g213 ( .A1(n_68), .A2(n_124), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_69), .B(n_130), .Y(n_170) );
INVx1_ASAP7_75t_L g524 ( .A(n_70), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_71), .B(n_130), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_72), .A2(n_455), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g164 ( .A(n_73), .B(n_120), .Y(n_164) );
INVx1_ASAP7_75t_L g126 ( .A(n_74), .Y(n_126) );
INVx1_ASAP7_75t_L g135 ( .A(n_74), .Y(n_135) );
AND2x2_ASAP7_75t_L g183 ( .A(n_75), .B(n_153), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_76), .B(n_474), .Y(n_517) );
AND2x2_ASAP7_75t_L g485 ( .A(n_78), .B(n_153), .Y(n_485) );
INVx1_ASAP7_75t_L g494 ( .A(n_79), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_80), .A2(n_455), .B(n_482), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_81), .A2(n_455), .B(n_460), .C(n_465), .Y(n_454) );
INVx1_ASAP7_75t_L g423 ( .A(n_82), .Y(n_423) );
AND2x2_ASAP7_75t_L g168 ( .A(n_83), .B(n_153), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_84), .B(n_130), .Y(n_202) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_85), .B(n_153), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_86), .A2(n_455), .B1(n_512), .B2(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g212 ( .A(n_87), .B(n_193), .Y(n_212) );
AND2x2_ASAP7_75t_L g156 ( .A(n_89), .B(n_153), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_90), .B(n_139), .Y(n_201) );
INVx1_ASAP7_75t_L g471 ( .A(n_91), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_92), .B(n_141), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_93), .B(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_94), .A2(n_124), .B(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g518 ( .A(n_95), .B(n_153), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_96), .B(n_141), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_97), .A2(n_539), .B(n_540), .C(n_542), .Y(n_538) );
BUFx2_ASAP7_75t_L g431 ( .A(n_98), .Y(n_431) );
BUFx2_ASAP7_75t_SL g790 ( .A(n_98), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_99), .A2(n_124), .B(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_100), .B(n_131), .Y(n_472) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_791), .B(n_802), .Y(n_101) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_432), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_429), .Y(n_103) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_416), .B(n_424), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
XOR2x1_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx3_ASAP7_75t_L g768 ( .A(n_110), .Y(n_768) );
OAI22xp5_ASAP7_75t_SL g776 ( .A1(n_110), .A2(n_777), .B1(n_779), .B2(n_780), .Y(n_776) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_328), .Y(n_110) );
AND4x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_240), .C(n_267), .D(n_302), .Y(n_111) );
AOI221xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_165), .B1(n_205), .B2(n_220), .C(n_224), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_144), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_115), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OR2x2_ASAP7_75t_L g281 ( .A(n_116), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g336 ( .A(n_116), .B(n_291), .Y(n_336) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g239 ( .A(n_117), .B(n_157), .Y(n_239) );
AND2x4_ASAP7_75t_L g275 ( .A(n_117), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g289 ( .A(n_117), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g206 ( .A(n_118), .Y(n_206) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_118), .Y(n_378) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_123), .B(n_143), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_119), .A2(n_170), .B(n_171), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g182 ( .A(n_119), .Y(n_182) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_119), .A2(n_123), .B(n_143), .Y(n_252) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_SL g120 ( .A(n_121), .B(n_122), .Y(n_120) );
AND2x4_ASAP7_75t_L g193 ( .A(n_121), .B(n_122), .Y(n_193) );
AND2x6_ASAP7_75t_L g124 ( .A(n_125), .B(n_127), .Y(n_124) );
BUFx3_ASAP7_75t_L g452 ( .A(n_125), .Y(n_452) );
AND2x6_ASAP7_75t_L g139 ( .A(n_126), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g459 ( .A(n_126), .Y(n_459) );
AND2x4_ASAP7_75t_L g455 ( .A(n_127), .B(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x4_ASAP7_75t_L g141 ( .A(n_128), .B(n_134), .Y(n_141) );
INVx2_ASAP7_75t_L g449 ( .A(n_128), .Y(n_449) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_129), .Y(n_450) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
INVx1_ASAP7_75t_L g495 ( .A(n_131), .Y(n_495) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_134), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx5_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_136), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_140), .B(n_142), .Y(n_137) );
INVxp67_ASAP7_75t_L g498 ( .A(n_139), .Y(n_498) );
INVxp67_ASAP7_75t_L g500 ( .A(n_141), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_142), .A2(n_149), .B(n_150), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_142), .A2(n_161), .B(n_162), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_142), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_142), .A2(n_179), .B(n_180), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_142), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_142), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_142), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_142), .A2(n_461), .B(n_462), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_142), .A2(n_464), .B(n_471), .C(n_472), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_142), .A2(n_464), .B(n_483), .C(n_484), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_142), .B(n_193), .Y(n_501) );
INVx1_ASAP7_75t_L g512 ( .A(n_142), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_142), .A2(n_464), .B(n_524), .C(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_SL g532 ( .A1(n_142), .A2(n_464), .B(n_533), .C(n_534), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_SL g233 ( .A1(n_144), .A2(n_206), .B(n_234), .C(n_238), .Y(n_233) );
AND2x2_ASAP7_75t_L g254 ( .A(n_144), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_144), .B(n_206), .Y(n_394) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_157), .Y(n_144) );
INVx2_ASAP7_75t_L g274 ( .A(n_145), .Y(n_274) );
BUFx3_ASAP7_75t_L g290 ( .A(n_145), .Y(n_290) );
INVxp67_ASAP7_75t_L g294 ( .A(n_145), .Y(n_294) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_152), .B(n_156), .Y(n_145) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_146), .A2(n_152), .B(n_156), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_152), .A2(n_158), .B(n_164), .Y(n_157) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_152), .A2(n_158), .B(n_164), .Y(n_219) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_152), .A2(n_520), .B(n_526), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_152), .A2(n_153), .B1(n_538), .B2(n_543), .Y(n_537) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_152), .A2(n_520), .B(n_526), .Y(n_556) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_154), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx4f_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
INVx2_ASAP7_75t_L g273 ( .A(n_157), .Y(n_273) );
AND2x2_ASAP7_75t_L g279 ( .A(n_157), .B(n_252), .Y(n_279) );
AND2x2_ASAP7_75t_L g305 ( .A(n_157), .B(n_274), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_159), .B(n_163), .Y(n_158) );
AOI211xp5_ASAP7_75t_L g302 ( .A1(n_165), .A2(n_303), .B(n_306), .C(n_316), .Y(n_302) );
AND2x2_ASAP7_75t_SL g165 ( .A(n_166), .B(n_184), .Y(n_165) );
OAI321xp33_ASAP7_75t_L g277 ( .A1(n_166), .A2(n_225), .A3(n_278), .B1(n_280), .B2(n_281), .C(n_283), .Y(n_277) );
AND2x2_ASAP7_75t_L g398 ( .A(n_166), .B(n_373), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_166), .Y(n_401) );
AND2x2_ASAP7_75t_L g166 ( .A(n_167), .B(n_175), .Y(n_166) );
INVx5_ASAP7_75t_L g223 ( .A(n_167), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_167), .B(n_237), .Y(n_236) );
NOR2x1_ASAP7_75t_SL g268 ( .A(n_167), .B(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g313 ( .A(n_167), .Y(n_313) );
AND2x2_ASAP7_75t_L g415 ( .A(n_167), .B(n_185), .Y(n_415) );
OR2x6_ASAP7_75t_L g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AND2x2_ASAP7_75t_L g222 ( .A(n_175), .B(n_223), .Y(n_222) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
INVx4_ASAP7_75t_L g237 ( .A(n_175), .Y(n_237) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_182), .B(n_183), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_181), .Y(n_176) );
AO21x2_ASAP7_75t_L g478 ( .A1(n_182), .A2(n_479), .B(n_485), .Y(n_478) );
INVx1_ASAP7_75t_L g280 ( .A(n_184), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_R g383 ( .A1(n_184), .A2(n_222), .B(n_254), .C(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g403 ( .A(n_184), .B(n_228), .Y(n_403) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_194), .Y(n_184) );
INVx1_ASAP7_75t_L g221 ( .A(n_185), .Y(n_221) );
INVx2_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
OR2x2_ASAP7_75t_L g246 ( .A(n_185), .B(n_237), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_185), .B(n_269), .Y(n_315) );
BUFx3_ASAP7_75t_L g322 ( .A(n_185), .Y(n_322) );
INVx2_ASAP7_75t_SL g465 ( .A(n_186), .Y(n_465) );
OA21x2_ASAP7_75t_L g530 ( .A1(n_186), .A2(n_531), .B(n_535), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_193), .Y(n_187) );
INVx1_ASAP7_75t_SL g196 ( .A(n_193), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_193), .B(n_218), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_193), .A2(n_469), .B(n_473), .Y(n_468) );
INVx1_ASAP7_75t_L g285 ( .A(n_194), .Y(n_285) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_194), .Y(n_298) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g231 ( .A(n_195), .Y(n_231) );
INVx1_ASAP7_75t_L g340 ( .A(n_195), .Y(n_340) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_203), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_196), .B(n_204), .Y(n_203) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_196), .A2(n_197), .B(n_203), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
AND2x2_ASAP7_75t_L g241 ( .A(n_205), .B(n_242), .Y(n_241) );
OAI31xp33_ASAP7_75t_L g392 ( .A1(n_205), .A2(n_393), .A3(n_395), .B(n_398), .Y(n_392) );
INVx1_ASAP7_75t_SL g410 ( .A(n_205), .Y(n_410) );
AND2x4_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AOI21xp33_ASAP7_75t_L g224 ( .A1(n_206), .A2(n_225), .B(n_233), .Y(n_224) );
NAND2x1_ASAP7_75t_L g304 ( .A(n_206), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_SL g333 ( .A(n_206), .Y(n_333) );
INVx2_ASAP7_75t_L g282 ( .A(n_207), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_207), .B(n_265), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_207), .B(n_264), .Y(n_374) );
NOR2xp33_ASAP7_75t_SL g382 ( .A(n_207), .B(n_333), .Y(n_382) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
AND2x2_ASAP7_75t_SL g251 ( .A(n_208), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g262 ( .A(n_208), .B(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g291 ( .A(n_208), .B(n_273), .Y(n_291) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
BUFx2_ASAP7_75t_L g255 ( .A(n_209), .Y(n_255) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g276 ( .A(n_210), .Y(n_276) );
OAI21x1_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_213), .B(n_217), .Y(n_210) );
INVx1_ASAP7_75t_L g218 ( .A(n_212), .Y(n_218) );
INVx2_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_219), .Y(n_323) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
INVx1_ASAP7_75t_L g259 ( .A(n_221), .Y(n_259) );
AND2x2_ASAP7_75t_L g338 ( .A(n_221), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g249 ( .A(n_222), .B(n_243), .Y(n_249) );
INVx2_ASAP7_75t_SL g297 ( .A(n_222), .Y(n_297) );
INVx4_ASAP7_75t_L g228 ( .A(n_223), .Y(n_228) );
AND2x2_ASAP7_75t_L g326 ( .A(n_223), .B(n_269), .Y(n_326) );
AND2x2_ASAP7_75t_SL g344 ( .A(n_223), .B(n_339), .Y(n_344) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_223), .B(n_237), .Y(n_361) );
INVx1_ASAP7_75t_L g367 ( .A(n_225), .Y(n_367) );
OR2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_229), .Y(n_225) );
INVx1_ASAP7_75t_L g286 ( .A(n_226), .Y(n_286) );
OR2x2_ASAP7_75t_L g299 ( .A(n_226), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_228), .Y(n_226) );
OR2x2_ASAP7_75t_L g351 ( .A(n_227), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g381 ( .A(n_227), .B(n_269), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_228), .B(n_231), .Y(n_257) );
AND2x2_ASAP7_75t_L g349 ( .A(n_228), .B(n_339), .Y(n_349) );
AND2x4_ASAP7_75t_L g411 ( .A(n_228), .B(n_290), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
INVx2_ASAP7_75t_L g235 ( .A(n_230), .Y(n_235) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2xp67_ASAP7_75t_SL g234 ( .A(n_235), .B(n_236), .Y(n_234) );
OAI322xp33_ASAP7_75t_SL g247 ( .A1(n_235), .A2(n_248), .A3(n_250), .B1(n_253), .B2(n_256), .C1(n_258), .C2(n_260), .Y(n_247) );
INVx1_ASAP7_75t_L g405 ( .A(n_235), .Y(n_405) );
OR2x2_ASAP7_75t_L g258 ( .A(n_236), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g284 ( .A(n_237), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_237), .B(n_285), .Y(n_300) );
INVx2_ASAP7_75t_L g327 ( .A(n_237), .Y(n_327) );
AND2x4_ASAP7_75t_L g339 ( .A(n_237), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_239), .B(n_255), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_245), .B(n_247), .Y(n_240) );
AND2x2_ASAP7_75t_L g308 ( .A(n_242), .B(n_275), .Y(n_308) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_243), .B(n_397), .Y(n_396) );
BUFx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
AND2x4_ASAP7_75t_SL g348 ( .A(n_244), .B(n_263), .Y(n_348) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g256 ( .A(n_246), .B(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_249), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g384 ( .A(n_251), .B(n_348), .Y(n_384) );
NOR4xp25_ASAP7_75t_L g388 ( .A(n_251), .B(n_265), .C(n_305), .D(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g265 ( .A(n_252), .B(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g301 ( .A(n_252), .B(n_276), .Y(n_301) );
AND2x4_ASAP7_75t_L g365 ( .A(n_252), .B(n_276), .Y(n_365) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_255), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
OR2x2_ASAP7_75t_L g354 ( .A(n_262), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g408 ( .A(n_262), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_263), .B(n_275), .Y(n_309) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AOI211xp5_ASAP7_75t_SL g267 ( .A1(n_268), .A2(n_270), .B(n_277), .C(n_292), .Y(n_267) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_275), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_273), .B(n_276), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_274), .B(n_279), .Y(n_278) );
BUFx2_ASAP7_75t_L g356 ( .A(n_274), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_275), .B(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g371 ( .A(n_275), .Y(n_371) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .B(n_287), .Y(n_283) );
AND2x4_ASAP7_75t_L g320 ( .A(n_284), .B(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g414 ( .A(n_284), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_SL g318 ( .A(n_290), .Y(n_318) );
AND2x2_ASAP7_75t_L g377 ( .A(n_291), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g391 ( .A(n_291), .Y(n_391) );
O2A1O1Ixp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_299), .C(n_301), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_293), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g369 ( .A(n_294), .B(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g390 ( .A(n_294), .B(n_391), .Y(n_390) );
INVxp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
OR2x2_ASAP7_75t_L g379 ( .A(n_297), .B(n_321), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_300), .A2(n_307), .B1(n_309), .B2(n_310), .Y(n_306) );
INVx1_ASAP7_75t_SL g397 ( .A(n_301), .Y(n_397) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_312), .B(n_321), .Y(n_363) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVxp67_ASAP7_75t_SL g373 ( .A(n_315), .Y(n_373) );
OAI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B1(n_323), .B2(n_324), .Y(n_316) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI21xp5_ASAP7_75t_SL g330 ( .A1(n_321), .A2(n_331), .B(n_334), .Y(n_330) );
AND2x2_ASAP7_75t_L g359 ( .A(n_321), .B(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND3x2_ASAP7_75t_L g325 ( .A(n_322), .B(n_326), .C(n_327), .Y(n_325) );
AND2x2_ASAP7_75t_L g387 ( .A(n_322), .B(n_344), .Y(n_387) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g372 ( .A(n_327), .B(n_373), .Y(n_372) );
NOR2xp67_ASAP7_75t_L g328 ( .A(n_329), .B(n_385), .Y(n_328) );
NAND4xp25_ASAP7_75t_L g329 ( .A(n_330), .B(n_345), .C(n_366), .D(n_383), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B1(n_341), .B2(n_343), .Y(n_334) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_337), .A2(n_351), .B1(n_371), .B2(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g352 ( .A(n_339), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_341), .A2(n_364), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx3_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_349), .B1(n_350), .B2(n_353), .C(n_357), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_362), .B1(n_363), .B2(n_364), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_360), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_360), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B1(n_372), .B2(n_374), .C(n_375), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_371), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_379), .B1(n_380), .B2(n_382), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_381), .A2(n_401), .B(n_402), .C(n_404), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_392), .C(n_399), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_406), .B1(n_409), .B2(n_411), .C(n_412), .Y(n_399) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g428 ( .A(n_417), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OR2x6_ASAP7_75t_SL g767 ( .A(n_418), .B(n_419), .Y(n_767) );
AND2x6_ASAP7_75t_SL g770 ( .A(n_418), .B(n_420), .Y(n_770) );
OR2x2_ASAP7_75t_L g785 ( .A(n_418), .B(n_420), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVxp33_ASAP7_75t_L g786 ( .A(n_424), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
AOI31xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_774), .A3(n_786), .B(n_787), .Y(n_432) );
NAND2xp5_ASAP7_75t_SL g433 ( .A(n_434), .B(n_771), .Y(n_433) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_767), .B1(n_768), .B2(n_769), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g779 ( .A(n_437), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g437 ( .A(n_438), .B(n_618), .C(n_684), .D(n_747), .Y(n_437) );
NOR2x1_ASAP7_75t_L g438 ( .A(n_439), .B(n_581), .Y(n_438) );
OR3x1_ASAP7_75t_L g439 ( .A(n_440), .B(n_551), .C(n_578), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_486), .B(n_507), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_475), .Y(n_442) );
AND2x2_ASAP7_75t_L g681 ( .A(n_443), .B(n_651), .Y(n_681) );
INVx1_ASAP7_75t_L g754 ( .A(n_443), .Y(n_754) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_466), .Y(n_443) );
INVx2_ASAP7_75t_L g506 ( .A(n_444), .Y(n_506) );
HB1xp67_ASAP7_75t_L g569 ( .A(n_444), .Y(n_569) );
AND2x2_ASAP7_75t_L g573 ( .A(n_444), .B(n_489), .Y(n_573) );
AND2x4_ASAP7_75t_L g589 ( .A(n_444), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g593 ( .A(n_444), .Y(n_593) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_454), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_451), .C(n_453), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g474 ( .A(n_448), .B(n_452), .Y(n_474) );
AND2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
OR2x6_ASAP7_75t_L g464 ( .A(n_449), .B(n_459), .Y(n_464) );
INVxp33_ASAP7_75t_L g515 ( .A(n_449), .Y(n_515) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g548 ( .A(n_455), .Y(n_548) );
NOR2x1p5_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx1_ASAP7_75t_L g516 ( .A(n_458), .Y(n_516) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_464), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_492) );
INVxp67_ASAP7_75t_L g539 ( .A(n_464), .Y(n_539) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_465), .A2(n_510), .B(n_518), .Y(n_509) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_465), .A2(n_510), .B(n_518), .Y(n_557) );
AND2x2_ASAP7_75t_L g487 ( .A(n_466), .B(n_488), .Y(n_487) );
INVx4_ASAP7_75t_L g570 ( .A(n_466), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_466), .B(n_560), .Y(n_574) );
INVx2_ASAP7_75t_L g588 ( .A(n_466), .Y(n_588) );
AND2x4_ASAP7_75t_L g592 ( .A(n_466), .B(n_593), .Y(n_592) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_466), .Y(n_627) );
OR2x2_ASAP7_75t_L g633 ( .A(n_466), .B(n_478), .Y(n_633) );
NOR2x1_ASAP7_75t_SL g662 ( .A(n_466), .B(n_489), .Y(n_662) );
NAND2xp5_ASAP7_75t_SL g764 ( .A(n_466), .B(n_736), .Y(n_764) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
INVx1_ASAP7_75t_L g550 ( .A(n_474), .Y(n_550) );
AND2x2_ASAP7_75t_L g661 ( .A(n_475), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2x1_ASAP7_75t_L g695 ( .A(n_476), .B(n_488), .Y(n_695) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g503 ( .A(n_478), .Y(n_503) );
INVx2_ASAP7_75t_L g561 ( .A(n_478), .Y(n_561) );
AND2x2_ASAP7_75t_L g584 ( .A(n_478), .B(n_489), .Y(n_584) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_478), .Y(n_611) );
INVx1_ASAP7_75t_L g652 ( .A(n_478), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_487), .B(n_502), .Y(n_486) );
AND2x2_ASAP7_75t_L g664 ( .A(n_487), .B(n_559), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_488), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g731 ( .A(n_488), .Y(n_731) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g590 ( .A(n_489), .Y(n_590) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_496), .B(n_501), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_495), .B(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_496) );
OAI211xp5_ASAP7_75t_SL g667 ( .A1(n_502), .A2(n_668), .B(n_672), .C(n_678), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_503), .B(n_504), .Y(n_502) );
AND2x2_ASAP7_75t_SL g583 ( .A(n_504), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_SL g714 ( .A(n_504), .Y(n_714) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g636 ( .A(n_506), .B(n_590), .Y(n_636) );
OR2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_527), .Y(n_507) );
AOI32xp33_ASAP7_75t_L g672 ( .A1(n_508), .A2(n_656), .A3(n_673), .B1(n_674), .B2(n_676), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_519), .Y(n_508) );
INVx2_ASAP7_75t_L g598 ( .A(n_509), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_509), .B(n_530), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_511), .B(n_517), .Y(n_510) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g610 ( .A(n_519), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_519), .B(n_536), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_519), .B(n_647), .Y(n_646) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_519), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
OR2x2_ASAP7_75t_L g629 ( .A(n_527), .B(n_630), .Y(n_629) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g580 ( .A(n_528), .B(n_554), .Y(n_580) );
AND2x2_ASAP7_75t_L g729 ( .A(n_528), .B(n_727), .Y(n_729) );
AND2x4_ASAP7_75t_L g528 ( .A(n_529), .B(n_536), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g566 ( .A(n_530), .Y(n_566) );
AND2x4_ASAP7_75t_L g605 ( .A(n_530), .B(n_606), .Y(n_605) );
INVxp67_ASAP7_75t_L g639 ( .A(n_530), .Y(n_639) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_530), .Y(n_647) );
AND2x2_ASAP7_75t_L g656 ( .A(n_530), .B(n_536), .Y(n_656) );
INVx1_ASAP7_75t_L g740 ( .A(n_530), .Y(n_740) );
INVx2_ASAP7_75t_L g577 ( .A(n_536), .Y(n_577) );
INVx1_ASAP7_75t_L g604 ( .A(n_536), .Y(n_604) );
INVx1_ASAP7_75t_L g671 ( .A(n_536), .Y(n_671) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_544), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OAI32xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_562), .A3(n_567), .B1(n_571), .B2(n_575), .Y(n_551) );
INVx1_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_553), .B(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_554), .B(n_614), .Y(n_613) );
AND2x2_ASAP7_75t_L g655 ( .A(n_554), .B(n_656), .Y(n_655) );
INVxp67_ASAP7_75t_L g680 ( .A(n_554), .Y(n_680) );
AND2x2_ASAP7_75t_L g761 ( .A(n_554), .B(n_603), .Y(n_761) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g576 ( .A(n_556), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g675 ( .A(n_556), .B(n_598), .Y(n_675) );
NOR2xp67_ASAP7_75t_L g697 ( .A(n_556), .B(n_577), .Y(n_697) );
NOR2x1_ASAP7_75t_L g739 ( .A(n_556), .B(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g606 ( .A(n_557), .Y(n_606) );
INVx1_ASAP7_75t_L g630 ( .A(n_557), .Y(n_630) );
AND2x2_ASAP7_75t_L g645 ( .A(n_557), .B(n_577), .Y(n_645) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g673 ( .A(n_559), .B(n_662), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_559), .B(n_592), .Y(n_743) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_560), .Y(n_712) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_561), .Y(n_694) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g595 ( .A(n_564), .B(n_596), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_564), .B(n_680), .Y(n_679) );
NOR2xp67_ASAP7_75t_SL g766 ( .A(n_564), .B(n_704), .Y(n_766) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g623 ( .A(n_566), .B(n_577), .Y(n_623) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_567), .B(n_633), .Y(n_691) );
INVx2_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_SL g657 ( .A(n_568), .B(n_584), .Y(n_657) );
AND2x4_ASAP7_75t_SL g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2x1_ASAP7_75t_L g616 ( .A(n_570), .B(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g722 ( .A(n_570), .B(n_593), .Y(n_722) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_570), .Y(n_751) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_571), .B(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
OR2x2_ASAP7_75t_L g693 ( .A(n_572), .B(n_694), .Y(n_693) );
NOR2x1_ASAP7_75t_L g758 ( .A(n_572), .B(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g682 ( .A(n_573), .B(n_627), .Y(n_682) );
INVxp33_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_576), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g756 ( .A(n_576), .B(n_638), .Y(n_756) );
INVx2_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_599), .Y(n_581) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_585), .B(n_594), .Y(n_582) );
AND2x2_ASAP7_75t_L g717 ( .A(n_584), .B(n_592), .Y(n_717) );
NAND2xp33_ASAP7_75t_R g585 ( .A(n_586), .B(n_591), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g759 ( .A(n_588), .Y(n_759) );
INVx4_ASAP7_75t_L g617 ( .A(n_589), .Y(n_617) );
INVx1_ASAP7_75t_L g736 ( .A(n_590), .Y(n_736) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g730 ( .A(n_592), .B(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_592), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_595), .A2(n_660), .B1(n_764), .B2(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g624 ( .A(n_598), .B(n_610), .Y(n_624) );
AND2x2_ASAP7_75t_L g638 ( .A(n_598), .B(n_639), .Y(n_638) );
A2O1A1Ixp33_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_607), .B(n_612), .C(n_615), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx3_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g686 ( .A(n_602), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g614 ( .A(n_603), .Y(n_614) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g674 ( .A(n_604), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g683 ( .A(n_604), .B(n_605), .Y(n_683) );
INVx1_ASAP7_75t_L g715 ( .A(n_604), .Y(n_715) );
AND2x4_ASAP7_75t_L g696 ( .A(n_605), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g718 ( .A(n_605), .B(n_609), .Y(n_718) );
AND2x2_ASAP7_75t_L g726 ( .A(n_605), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g701 ( .A(n_609), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_609), .B(n_623), .Y(n_703) );
AND2x2_ASAP7_75t_L g706 ( .A(n_609), .B(n_656), .Y(n_706) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_610), .B(n_671), .Y(n_720) );
AND2x2_ASAP7_75t_L g648 ( .A(n_611), .B(n_636), .Y(n_648) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g744 ( .A(n_614), .B(n_624), .Y(n_744) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_616), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g628 ( .A(n_617), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_617), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_658), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_642), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_625), .B1(n_629), .B2(n_631), .C1(n_634), .C2(n_637), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_627), .B(n_636), .Y(n_635) );
OR2x6_ASAP7_75t_L g707 ( .A(n_627), .B(n_677), .Y(n_707) );
NAND5xp2_ASAP7_75t_L g710 ( .A(n_627), .B(n_630), .C(n_646), .D(n_711), .E(n_713), .Y(n_710) );
NAND2x1_ASAP7_75t_L g746 ( .A(n_628), .B(n_632), .Y(n_746) );
INVx2_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NOR2x1_ASAP7_75t_L g676 ( .A(n_633), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_635), .A2(n_726), .B1(n_729), .B2(n_730), .Y(n_725) );
INVx2_ASAP7_75t_L g677 ( .A(n_636), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_636), .B(n_652), .Y(n_689) );
INVx3_ASAP7_75t_L g724 ( .A(n_637), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
AND2x2_ASAP7_75t_L g669 ( .A(n_638), .B(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g702 ( .A(n_638), .Y(n_702) );
INVx2_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g665 ( .A(n_641), .B(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_643), .B(n_654), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_648), .B(n_649), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g653 ( .A(n_645), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_648), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_653), .Y(n_649) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x4_ASAP7_75t_SL g735 ( .A(n_652), .B(n_736), .Y(n_735) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_659), .B(n_667), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B(n_665), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
BUFx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g704 ( .A(n_675), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B1(n_682), .B2(n_683), .Y(n_678) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_708), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .C(n_698), .Y(n_685) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
BUFx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OA21x2_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B(n_696), .Y(n_690) );
NAND2xp33_ASAP7_75t_SL g692 ( .A(n_693), .B(n_695), .Y(n_692) );
AOI21xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_705), .B(n_707), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .B(n_703), .C(n_704), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_702), .A2(n_742), .B1(n_744), .B2(n_745), .Y(n_741) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_732), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g709 ( .A(n_710), .B(n_716), .C(n_723), .D(n_725), .Y(n_709) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g721 ( .A(n_712), .B(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_L g752 ( .A(n_715), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_719), .B2(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_721), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI21xp5_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_737), .B(n_741), .Y(n_732) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_762), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B(n_753), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B1(n_757), .B2(n_760), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
CKINVDCx11_ASAP7_75t_R g778 ( .A(n_767), .Y(n_778) );
CKINVDCx11_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_770), .Y(n_782) );
INVx1_ASAP7_75t_L g775 ( .A(n_771), .Y(n_775) );
AOI21xp33_ASAP7_75t_SL g774 ( .A1(n_775), .A2(n_776), .B(n_783), .Y(n_774) );
INVx1_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx4_ASAP7_75t_SL g780 ( .A(n_781), .Y(n_780) );
INVx3_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_788), .Y(n_787) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx8_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_SL g791 ( .A(n_792), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_793), .Y(n_792) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_794), .Y(n_805) );
OR2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
CKINVDCx16_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
endmodule