module fake_jpeg_14664_n_23 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_23);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_23;

wire n_13;
wire n_21;
wire n_10;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_7),
.B(n_4),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx3_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_11),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_16),
.C(n_12),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_12),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_15),
.B(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_21),
.B(n_0),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_1),
.C(n_9),
.Y(n_23)
);


endmodule