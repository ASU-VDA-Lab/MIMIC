module fake_jpeg_1298_n_209 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_209);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_1),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_17),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_66),
.CON(n_75),
.SN(n_75)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_72),
.B1(n_65),
.B2(n_57),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_67),
.B1(n_61),
.B2(n_53),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_88),
.B1(n_86),
.B2(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_84),
.B(n_87),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_85),
.A2(n_51),
.B1(n_66),
.B2(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_71),
.Y(n_87)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_57),
.B1(n_67),
.B2(n_72),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_100),
.B1(n_51),
.B2(n_73),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_91),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_109),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_72),
.B1(n_65),
.B2(n_69),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_52),
.B1(n_59),
.B2(n_58),
.Y(n_120)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_63),
.C(n_54),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_69),
.C(n_56),
.Y(n_130)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_113),
.Y(n_116)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_103),
.B1(n_100),
.B2(n_110),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_114),
.A2(n_118),
.B1(n_122),
.B2(n_131),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_37),
.B(n_35),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_70),
.B1(n_73),
.B2(n_63),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_120),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_102),
.B1(n_108),
.B2(n_104),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_62),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_124),
.B(n_125),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_66),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_131),
.C(n_130),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_55),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_0),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_49),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_56),
.B(n_2),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_135),
.A2(n_7),
.B(n_9),
.Y(n_168)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_138),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_116),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_150),
.C(n_153),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_138),
.C(n_150),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_133),
.A2(n_3),
.B(n_4),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_120),
.A2(n_48),
.B1(n_47),
.B2(n_46),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_149),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_38),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_121),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_4),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_31),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_30),
.C(n_29),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_161),
.C(n_165),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_154),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_27),
.C(n_22),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_21),
.B(n_6),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_168),
.B1(n_175),
.B2(n_166),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_166),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_10),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_174),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_157),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_183),
.C(n_171),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_135),
.B(n_144),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_184),
.B1(n_186),
.B2(n_169),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_145),
.C(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_148),
.B1(n_12),
.B2(n_13),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_161),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_162),
.C(n_167),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_192),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_172),
.C(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_194),
.A2(n_164),
.B(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_181),
.B1(n_176),
.B2(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g201 ( 
.A1(n_199),
.A2(n_193),
.A3(n_191),
.B1(n_192),
.B2(n_173),
.C1(n_19),
.C2(n_20),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_198),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_202),
.Y(n_204)
);

OAI21x1_ASAP7_75t_SL g205 ( 
.A1(n_204),
.A2(n_200),
.B(n_195),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_197),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_196),
.C(n_14),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_11),
.C(n_14),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_208),
.A2(n_16),
.B(n_17),
.Y(n_209)
);


endmodule