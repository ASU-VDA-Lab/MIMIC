module fake_jpeg_26379_n_338 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_14),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_19),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_28),
.Y(n_69)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_20),
.B1(n_18),
.B2(n_27),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_57),
.B1(n_63),
.B2(n_33),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_66),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_43),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_38),
.A2(n_20),
.B1(n_27),
.B2(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_33),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_20),
.B1(n_26),
.B2(n_29),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_26),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_73),
.B(n_85),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_74),
.B(n_80),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_50),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_76),
.A2(n_93),
.B1(n_99),
.B2(n_100),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_77),
.A2(n_79),
.B1(n_84),
.B2(n_98),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_68),
.A2(n_45),
.B1(n_24),
.B2(n_18),
.Y(n_79)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_42),
.CI(n_44),
.CON(n_80),
.SN(n_80)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_18),
.B1(n_67),
.B2(n_54),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_56),
.B1(n_48),
.B2(n_64),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_32),
.B1(n_34),
.B2(n_41),
.Y(n_110)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_51),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_95),
.Y(n_113)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_25),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_44),
.C(n_39),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_35),
.C(n_41),
.Y(n_111)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_96),
.Y(n_109)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_23),
.B1(n_33),
.B2(n_30),
.Y(n_99)
);

AO22x2_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_44),
.B1(n_41),
.B2(n_39),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_60),
.B1(n_31),
.B2(n_17),
.Y(n_133)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_103),
.B(n_104),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_59),
.B(n_34),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_53),
.B1(n_24),
.B2(n_59),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_107),
.A2(n_133),
.B1(n_117),
.B2(n_108),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_110),
.A2(n_102),
.B1(n_91),
.B2(n_82),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_94),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_119),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_87),
.A2(n_32),
.B1(n_34),
.B2(n_39),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_126),
.B1(n_97),
.B2(n_96),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_72),
.A2(n_32),
.B1(n_25),
.B2(n_30),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_76),
.A2(n_0),
.B(n_1),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_131),
.B(n_82),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_17),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_25),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_25),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_111),
.B1(n_132),
.B2(n_120),
.Y(n_165)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_137),
.Y(n_171)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_80),
.B(n_95),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_138),
.A2(n_139),
.B(n_154),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_80),
.B(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_142),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_164),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_144),
.A2(n_166),
.B1(n_133),
.B2(n_128),
.Y(n_178)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_126),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_149),
.B1(n_158),
.B2(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_75),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_157),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g148 ( 
.A(n_106),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_81),
.B1(n_88),
.B2(n_92),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_150),
.A2(n_128),
.B1(n_112),
.B2(n_91),
.Y(n_186)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_108),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_156),
.A2(n_160),
.B(n_133),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_105),
.B(n_83),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_83),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_163),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_101),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_160),
.B1(n_154),
.B2(n_139),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_129),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_179),
.B(n_0),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_198),
.B1(n_134),
.B2(n_164),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_136),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_147),
.B(n_113),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_178),
.A2(n_186),
.B1(n_187),
.B2(n_194),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_160),
.A2(n_125),
.B(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_183),
.Y(n_210)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_184),
.B(n_199),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_141),
.A2(n_127),
.B1(n_131),
.B2(n_122),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_157),
.B(n_131),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_191),
.B(n_192),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_110),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_143),
.B(n_101),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_196),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_86),
.B1(n_90),
.B2(n_30),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_138),
.A2(n_16),
.B(n_17),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_22),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_86),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_144),
.A2(n_30),
.B1(n_31),
.B2(n_17),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_166),
.A2(n_16),
.B1(n_22),
.B2(n_31),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_52),
.C(n_31),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_31),
.C(n_17),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_201),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_174),
.A2(n_153),
.B1(n_151),
.B2(n_137),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_203),
.A2(n_204),
.B1(n_211),
.B2(n_212),
.Y(n_232)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_201),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_214),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_16),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_216),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_220),
.C(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_170),
.A2(n_31),
.B1(n_17),
.B2(n_16),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_179),
.A2(n_17),
.B1(n_31),
.B2(n_22),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_213),
.A2(n_229),
.B(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_189),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_22),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_15),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_219),
.B(n_225),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_168),
.B(n_15),
.C(n_13),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_223),
.A2(n_192),
.B1(n_199),
.B2(n_185),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_189),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_168),
.B(n_12),
.C(n_11),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_176),
.B(n_12),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_228),
.Y(n_233)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_190),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_2),
.Y(n_230)
);

AO21x2_ASAP7_75t_L g231 ( 
.A1(n_217),
.A2(n_184),
.B(n_186),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_231),
.A2(n_245),
.B1(n_247),
.B2(n_223),
.Y(n_262)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_246),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_239),
.A2(n_241),
.B1(n_253),
.B2(n_255),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_216),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_221),
.A2(n_190),
.B1(n_183),
.B2(n_181),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_187),
.B1(n_197),
.B2(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_172),
.B1(n_180),
.B2(n_173),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_167),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_221),
.A2(n_185),
.B1(n_191),
.B2(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_177),
.C(n_173),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_230),
.C(n_207),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_167),
.B1(n_177),
.B2(n_175),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_256),
.B(n_259),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

AOI221xp5_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_224),
.B1(n_212),
.B2(n_230),
.C(n_220),
.Y(n_259)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_218),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_266),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_233),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_265),
.B(n_258),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_244),
.B(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_255),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_270),
.Y(n_276)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_209),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_278)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_241),
.Y(n_272)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_207),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_2),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_231),
.B1(n_245),
.B2(n_232),
.Y(n_277)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_238),
.C(n_239),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_280),
.C(n_283),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_238),
.C(n_232),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_231),
.C(n_250),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_231),
.B1(n_250),
.B2(n_235),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_288),
.A2(n_289),
.B1(n_264),
.B2(n_260),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_231),
.B1(n_169),
.B2(n_11),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_269),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_2),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_273),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_304),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_276),
.Y(n_297)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_297),
.Y(n_312)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_262),
.B(n_256),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_276),
.B(n_285),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_286),
.A2(n_263),
.B1(n_169),
.B2(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_301),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_279),
.B(n_280),
.C(n_278),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_9),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_303),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_9),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_281),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_3),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_306),
.A2(n_298),
.B(n_292),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_307),
.A2(n_309),
.B(n_313),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_277),
.B1(n_288),
.B2(n_284),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_294),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_310),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_295),
.A2(n_3),
.B(n_4),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_3),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_314),
.B(n_4),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_319),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_301),
.C(n_294),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_320),
.B(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_5),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_321),
.B(n_324),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_296),
.B(n_7),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_308),
.B(n_6),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_315),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_315),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_325),
.C(n_312),
.Y(n_332)
);

AOI21xp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_326),
.B(n_332),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_330),
.B(n_329),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_311),
.B(n_7),
.Y(n_336)
);

AOI211xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_8),
.C(n_316),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g338 ( 
.A(n_337),
.B(n_8),
.Y(n_338)
);


endmodule