module fake_aes_11968_n_657 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_657);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_657;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx16_ASAP7_75t_R g78 ( .A(n_60), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_70), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_32), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_74), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_30), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_29), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_14), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_28), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_44), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
INVx2_ASAP7_75t_L g89 ( .A(n_57), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_19), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_72), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_6), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_50), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_47), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_68), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_3), .Y(n_98) );
BUFx2_ASAP7_75t_L g99 ( .A(n_36), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_3), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_9), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_58), .Y(n_102) );
XOR2xp5_ASAP7_75t_L g103 ( .A(n_66), .B(n_10), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_48), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_41), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_65), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_33), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_2), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_25), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_69), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_27), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_31), .Y(n_116) );
INVxp67_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_53), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_62), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_40), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_52), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
INVx3_ASAP7_75t_L g123 ( .A(n_98), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_89), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_87), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_99), .B(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
BUFx2_ASAP7_75t_L g131 ( .A(n_99), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_104), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_101), .B(n_0), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_84), .B(n_1), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
INVxp33_ASAP7_75t_SL g137 ( .A(n_103), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_92), .A2(n_1), .B1(n_2), .B2(n_4), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_105), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_83), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_100), .B(n_4), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_92), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_110), .B(n_5), .Y(n_146) );
OAI22x1_ASAP7_75t_L g147 ( .A1(n_103), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_78), .B(n_7), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_111), .B(n_8), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_85), .B(n_11), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_86), .B(n_11), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_95), .B(n_12), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_97), .B(n_13), .Y(n_154) );
INVxp67_ASAP7_75t_L g155 ( .A(n_102), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_106), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g157 ( .A1(n_118), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_107), .B(n_15), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_129), .B(n_113), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_136), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_129), .B(n_109), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_131), .B(n_121), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_129), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g166 ( .A(n_137), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_131), .Y(n_170) );
BUFx4f_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
OR2x6_ASAP7_75t_L g172 ( .A(n_140), .B(n_117), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_136), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_123), .Y(n_174) );
AND2x6_ASAP7_75t_L g175 ( .A(n_152), .B(n_114), .Y(n_175) );
INVx5_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_149), .Y(n_177) );
BUFx10_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_148), .Y(n_180) );
HB1xp67_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_123), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_123), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_122), .B(n_116), .Y(n_186) );
OR2x6_ASAP7_75t_L g187 ( .A(n_140), .B(n_108), .Y(n_187) );
NOR2x1p5_ASAP7_75t_L g188 ( .A(n_145), .B(n_121), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_157), .Y(n_189) );
BUFx3_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
AND2x6_ASAP7_75t_L g191 ( .A(n_149), .B(n_120), .Y(n_191) );
BUFx4f_ASAP7_75t_L g192 ( .A(n_149), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_155), .B(n_91), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_149), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_136), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_143), .B(n_91), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_127), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_122), .A2(n_119), .B1(n_115), .B2(n_93), .Y(n_199) );
AND2x6_ASAP7_75t_L g200 ( .A(n_128), .B(n_90), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_128), .B(n_93), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_133), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_143), .B(n_90), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_159), .A2(n_130), .B1(n_156), .B2(n_138), .Y(n_204) );
OR2x6_ASAP7_75t_L g205 ( .A(n_188), .B(n_147), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_193), .B(n_142), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_197), .B(n_130), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_203), .B(n_158), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_163), .B(n_154), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_198), .Y(n_210) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_159), .A2(n_134), .B1(n_151), .B2(n_150), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_192), .B(n_133), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_170), .B(n_135), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_164), .B(n_144), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_202), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_159), .A2(n_156), .B1(n_153), .B2(n_138), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_181), .B(n_147), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_164), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_160), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_159), .A2(n_156), .B1(n_153), .B2(n_138), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_192), .B(n_133), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_164), .B(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_171), .B(n_79), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_159), .A2(n_153), .B1(n_127), .B2(n_126), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_201), .B(n_132), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_192), .B(n_132), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_201), .B(n_126), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_200), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_200), .B(n_127), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_200), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_199), .B(n_112), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_200), .B(n_81), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_165), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_167), .B(n_141), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_172), .B(n_139), .Y(n_236) );
INVxp67_ASAP7_75t_SL g237 ( .A(n_171), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_200), .B(n_81), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_199), .B(n_112), .Y(n_239) );
INVxp33_ASAP7_75t_L g240 ( .A(n_186), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_178), .B(n_79), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
AOI22xp5_ASAP7_75t_L g243 ( .A1(n_162), .A2(n_125), .B1(n_124), .B2(n_139), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_178), .B(n_125), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_162), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_177), .A2(n_124), .B(n_17), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_162), .A2(n_16), .B1(n_20), .B2(n_21), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_162), .B(n_16), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g249 ( .A(n_175), .B(n_22), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_162), .B(n_23), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_178), .B(n_24), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_191), .A2(n_26), .B1(n_37), .B2(n_38), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_195), .B(n_39), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_191), .B(n_42), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_179), .B(n_43), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_191), .B(n_45), .Y(n_257) );
BUFx8_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_220), .Y(n_259) );
NOR2xp67_ASAP7_75t_L g260 ( .A(n_236), .B(n_166), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_213), .B(n_172), .Y(n_261) );
O2A1O1Ixp5_ASAP7_75t_L g262 ( .A1(n_251), .A2(n_186), .B(n_179), .C(n_184), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_206), .B(n_166), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_218), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_206), .B(n_189), .Y(n_266) );
NOR2xp33_ASAP7_75t_R g267 ( .A(n_232), .B(n_189), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_219), .B(n_179), .Y(n_268) );
INVx4_ASAP7_75t_L g269 ( .A(n_218), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_208), .A2(n_184), .B(n_174), .Y(n_270) );
OAI21xp33_ASAP7_75t_SL g271 ( .A1(n_207), .A2(n_184), .B(n_187), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g272 ( .A1(n_234), .A2(n_174), .B(n_185), .C(n_190), .Y(n_272) );
O2A1O1Ixp5_ASAP7_75t_SL g273 ( .A1(n_251), .A2(n_161), .B(n_196), .C(n_176), .Y(n_273) );
OR2x6_ASAP7_75t_SL g274 ( .A(n_205), .B(n_187), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_223), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_229), .B(n_176), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_237), .B(n_191), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_239), .B(n_172), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_SL g279 ( .A1(n_255), .A2(n_185), .B(n_194), .C(n_168), .Y(n_279) );
INVx4_ASAP7_75t_L g280 ( .A(n_229), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_223), .Y(n_281) );
NOR2xp33_ASAP7_75t_R g282 ( .A(n_249), .B(n_191), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_209), .B(n_172), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_230), .A2(n_190), .B(n_183), .Y(n_284) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_242), .A2(n_183), .B(n_176), .C(n_168), .Y(n_285) );
NOR2xp67_ASAP7_75t_SL g286 ( .A(n_229), .B(n_175), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_205), .B(n_187), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_244), .A2(n_176), .B(n_194), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_210), .Y(n_289) );
AOI21xp5_ASAP7_75t_L g290 ( .A1(n_212), .A2(n_182), .B(n_173), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_215), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_205), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_214), .A2(n_175), .B1(n_187), .B2(n_182), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_229), .B(n_196), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g295 ( .A1(n_226), .A2(n_173), .B(n_175), .C(n_196), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_214), .B(n_175), .Y(n_296) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_228), .A2(n_196), .B(n_161), .C(n_51), .Y(n_297) );
NAND2xp33_ASAP7_75t_L g298 ( .A(n_245), .B(n_161), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_211), .A2(n_161), .B1(n_49), .B2(n_54), .Y(n_299) );
NOR2xp33_ASAP7_75t_R g300 ( .A(n_248), .B(n_46), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_235), .B(n_55), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_235), .B(n_56), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g303 ( .A1(n_212), .A2(n_59), .B(n_61), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_222), .A2(n_64), .B(n_67), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g305 ( .A1(n_204), .A2(n_71), .B1(n_73), .B2(n_75), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_266), .A2(n_240), .B1(n_241), .B2(n_224), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_271), .A2(n_227), .B(n_222), .C(n_244), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_259), .B(n_210), .Y(n_308) );
O2A1O1Ixp33_ASAP7_75t_SL g309 ( .A1(n_272), .A2(n_250), .B(n_257), .C(n_247), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_258), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_SL g311 ( .A1(n_301), .A2(n_256), .B(n_246), .C(n_254), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_291), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_279), .A2(n_227), .B(n_256), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_275), .Y(n_314) );
O2A1O1Ixp5_ASAP7_75t_L g315 ( .A1(n_262), .A2(n_254), .B(n_233), .C(n_238), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_283), .B(n_216), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_267), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_273), .A2(n_252), .B(n_253), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_263), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_264), .A2(n_252), .B(n_231), .C(n_221), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_268), .A2(n_243), .B(n_225), .C(n_77), .Y(n_321) );
A2O1A1Ixp33_ASAP7_75t_L g322 ( .A1(n_270), .A2(n_268), .B(n_293), .C(n_301), .Y(n_322) );
NOR2xp67_ASAP7_75t_SL g323 ( .A(n_292), .B(n_280), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_258), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_281), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g326 ( .A1(n_270), .A2(n_302), .B(n_295), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g327 ( .A1(n_302), .A2(n_284), .B(n_289), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_285), .A2(n_304), .B(n_303), .C(n_299), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g329 ( .A(n_287), .B(n_260), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_280), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_261), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_290), .A2(n_297), .B(n_296), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_277), .A2(n_278), .B1(n_269), .B2(n_274), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_282), .B(n_304), .Y(n_334) );
O2A1O1Ixp33_ASAP7_75t_SL g335 ( .A1(n_303), .A2(n_305), .B(n_276), .C(n_290), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_294), .Y(n_336) );
AO31x2_ASAP7_75t_L g337 ( .A1(n_288), .A2(n_265), .A3(n_269), .B(n_300), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g338 ( .A(n_286), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_308), .Y(n_339) );
AO31x2_ASAP7_75t_L g340 ( .A1(n_322), .A2(n_294), .A3(n_298), .B(n_277), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_311), .A2(n_328), .B(n_335), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_311), .A2(n_328), .B(n_335), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_312), .B(n_329), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_330), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_319), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_327), .A2(n_326), .B(n_332), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_309), .A2(n_334), .B(n_322), .Y(n_347) );
AO31x2_ASAP7_75t_L g348 ( .A1(n_313), .A2(n_336), .A3(n_316), .B(n_325), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_331), .B(n_306), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_333), .B(n_317), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_314), .B(n_323), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_336), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_330), .Y(n_353) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_318), .A2(n_315), .B(n_334), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_320), .B(n_307), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
AO31x2_ASAP7_75t_L g358 ( .A1(n_309), .A2(n_337), .A3(n_321), .B(n_338), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_310), .A2(n_283), .B1(n_266), .B2(n_264), .C(n_217), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_337), .A2(n_326), .B(n_322), .Y(n_360) );
AO31x2_ASAP7_75t_L g361 ( .A1(n_337), .A2(n_322), .A3(n_313), .B(n_299), .Y(n_361) );
OAI22xp5_ASAP7_75t_SL g362 ( .A1(n_324), .A2(n_137), .B1(n_145), .B2(n_172), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_317), .B(n_137), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_322), .A2(n_271), .B(n_270), .C(n_307), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_312), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_352), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_344), .Y(n_368) );
INVxp67_ASAP7_75t_SL g369 ( .A(n_357), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_365), .A2(n_356), .B(n_346), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
AO21x2_ASAP7_75t_L g372 ( .A1(n_341), .A2(n_342), .B(n_347), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_363), .B(n_348), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_366), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_365), .A2(n_354), .B(n_346), .Y(n_375) );
AO21x2_ASAP7_75t_L g376 ( .A1(n_349), .A2(n_366), .B(n_350), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_363), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_344), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_348), .B(n_360), .Y(n_379) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_359), .A2(n_360), .B(n_345), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_357), .Y(n_381) );
BUFx3_ASAP7_75t_L g382 ( .A(n_353), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_348), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_348), .B(n_360), .Y(n_384) );
AO21x2_ASAP7_75t_L g385 ( .A1(n_355), .A2(n_351), .B(n_361), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_353), .B1(n_343), .B2(n_357), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_348), .B(n_340), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_361), .A2(n_354), .B(n_358), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_340), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_340), .B(n_361), .Y(n_391) );
INVx2_ASAP7_75t_SL g392 ( .A(n_343), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_340), .B(n_343), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_340), .A2(n_361), .B(n_358), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_358), .B(n_361), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_358), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_358), .B(n_364), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_382), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_392), .B(n_362), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_374), .B(n_377), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_388), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_373), .B(n_367), .Y(n_402) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_382), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_374), .B(n_376), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_373), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_373), .B(n_367), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_397), .B(n_376), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_388), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_376), .B(n_380), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_376), .B(n_380), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_383), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_397), .B(n_377), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_383), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_382), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_392), .A2(n_397), .B1(n_386), .B2(n_368), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_386), .A2(n_393), .B1(n_392), .B2(n_391), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
AND2x4_ASAP7_75t_SL g420 ( .A(n_368), .B(n_378), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_371), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_368), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_371), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_379), .B(n_384), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_381), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_381), .B(n_384), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_385), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_393), .B(n_385), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_391), .B(n_384), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_391), .B(n_379), .Y(n_431) );
INVxp67_ASAP7_75t_SL g432 ( .A(n_369), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_379), .B(n_385), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_378), .Y(n_434) );
INVx5_ASAP7_75t_L g435 ( .A(n_378), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_385), .B(n_370), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_387), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_385), .B(n_370), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_390), .B(n_387), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_430), .B(n_390), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_430), .B(n_394), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_405), .B(n_394), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_424), .B(n_395), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_405), .B(n_426), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_431), .B(n_389), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_431), .B(n_389), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_433), .B(n_389), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_433), .B(n_389), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_402), .B(n_395), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_402), .B(n_389), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_407), .B(n_395), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_407), .B(n_396), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_424), .B(n_396), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_436), .B(n_396), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_436), .B(n_372), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_436), .B(n_372), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_426), .B(n_372), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_413), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_421), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_421), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_438), .B(n_372), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_438), .B(n_375), .Y(n_464) );
INVx5_ASAP7_75t_L g465 ( .A(n_435), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_438), .B(n_375), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_401), .Y(n_467) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_429), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_426), .B(n_437), .Y(n_469) );
AND2x2_ASAP7_75t_SL g470 ( .A(n_406), .B(n_417), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_414), .B(n_408), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_426), .B(n_437), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_423), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_435), .B(n_434), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_400), .B(n_423), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_415), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_440), .B(n_415), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_415), .B(n_414), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_404), .Y(n_479) );
NOR2x1_ASAP7_75t_L g480 ( .A(n_406), .B(n_429), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_429), .B(n_428), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_408), .B(n_428), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_404), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_399), .B(n_420), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_409), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_410), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_398), .B(n_403), .Y(n_487) );
NOR2x1_ASAP7_75t_SL g488 ( .A(n_435), .B(n_434), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_429), .B(n_419), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_419), .B(n_427), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_416), .B(n_422), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_425), .B(n_419), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_441), .B(n_417), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_477), .B(n_432), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_471), .B(n_410), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_470), .A2(n_418), .B1(n_439), .B2(n_427), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_446), .B(n_425), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_477), .B(n_420), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_461), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_442), .B(n_420), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_442), .B(n_411), .Y(n_501) );
NAND3xp33_ASAP7_75t_L g502 ( .A(n_468), .B(n_411), .C(n_412), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_470), .A2(n_435), .B1(n_412), .B2(n_425), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_441), .B(n_435), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_467), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_446), .B(n_425), .Y(n_506) );
INVx1_ASAP7_75t_SL g507 ( .A(n_487), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_447), .B(n_435), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g509 ( .A(n_465), .B(n_474), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
INVx2_ASAP7_75t_SL g511 ( .A(n_465), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_484), .B(n_487), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_467), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_471), .B(n_482), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_482), .B(n_444), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_462), .Y(n_516) );
BUFx2_ASAP7_75t_L g517 ( .A(n_465), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_469), .B(n_472), .Y(n_518) );
INVxp67_ASAP7_75t_L g519 ( .A(n_488), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_462), .Y(n_520) );
NAND2x1_ASAP7_75t_L g521 ( .A(n_480), .B(n_488), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_447), .B(n_478), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_491), .B(n_444), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_469), .B(n_472), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_451), .B(n_453), .Y(n_526) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_470), .B(n_450), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_455), .B(n_478), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_467), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_473), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_449), .B(n_450), .Y(n_531) );
OR2x6_ASAP7_75t_L g532 ( .A(n_480), .B(n_459), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_465), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_449), .B(n_455), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_452), .B(n_475), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_452), .B(n_445), .Y(n_536) );
INVx4_ASAP7_75t_L g537 ( .A(n_465), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_454), .B(n_443), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_454), .B(n_443), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_448), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_445), .B(n_481), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_445), .B(n_481), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_445), .B(n_443), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_443), .B(n_463), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_448), .B(n_460), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_460), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_476), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_507), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_499), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_544), .B(n_459), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_505), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_505), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_510), .Y(n_553) );
INVx2_ASAP7_75t_SL g554 ( .A(n_537), .Y(n_554) );
NAND2xp33_ASAP7_75t_L g555 ( .A(n_511), .B(n_465), .Y(n_555) );
INVxp67_ASAP7_75t_SL g556 ( .A(n_519), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_524), .B(n_483), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_513), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_495), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_514), .B(n_479), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_516), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_520), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_512), .B(n_479), .Y(n_564) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_527), .A2(n_483), .B1(n_459), .B2(n_458), .C(n_457), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_544), .B(n_459), .Y(n_566) );
OAI222xp33_ASAP7_75t_L g567 ( .A1(n_519), .A2(n_457), .B1(n_458), .B2(n_463), .C1(n_476), .C2(n_464), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_536), .B(n_464), .Y(n_568) );
INVxp67_ASAP7_75t_SL g569 ( .A(n_521), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_512), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_531), .B(n_489), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_536), .B(n_466), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_518), .B(n_466), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_525), .B(n_489), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_517), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_540), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_546), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_513), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_522), .B(n_490), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_496), .A2(n_490), .B(n_456), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_547), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_528), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_497), .B(n_456), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_529), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_545), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_527), .A2(n_468), .B1(n_492), .B2(n_486), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_497), .B(n_492), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_524), .B(n_485), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_589), .B(n_493), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_560), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_560), .Y(n_592) );
AOI22xp5_ASAP7_75t_L g593 ( .A1(n_581), .A2(n_496), .B1(n_501), .B2(n_500), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_564), .B(n_535), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_586), .Y(n_595) );
OAI31xp33_ASAP7_75t_L g596 ( .A1(n_569), .A2(n_509), .A3(n_511), .B(n_533), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_554), .Y(n_597) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_548), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_570), .B(n_515), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_586), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_559), .B(n_534), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_583), .B(n_526), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_557), .B(n_542), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_555), .A2(n_537), .B(n_509), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_582), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_554), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_573), .B(n_538), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_582), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_573), .B(n_539), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_549), .Y(n_610) );
NOR3xp33_ASAP7_75t_L g611 ( .A(n_581), .B(n_537), .C(n_502), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_550), .B(n_541), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_551), .Y(n_613) );
OAI211xp5_ASAP7_75t_SL g614 ( .A1(n_565), .A2(n_503), .B(n_508), .C(n_504), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_575), .B(n_543), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_604), .A2(n_556), .B(n_567), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_599), .B(n_575), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g618 ( .A1(n_599), .A2(n_572), .B1(n_568), .B2(n_563), .C(n_561), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_606), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_601), .B(n_571), .Y(n_620) );
INVx1_ASAP7_75t_SL g621 ( .A(n_606), .Y(n_621) );
OAI21xp5_ASAP7_75t_SL g622 ( .A1(n_596), .A2(n_587), .B(n_498), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_532), .B(n_494), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_595), .B(n_553), .Y(n_624) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_611), .A2(n_566), .B(n_550), .C(n_572), .Y(n_625) );
AOI221x1_ASAP7_75t_SL g626 ( .A1(n_602), .A2(n_553), .B1(n_578), .B2(n_577), .C(n_576), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_611), .A2(n_568), .B1(n_576), .B2(n_561), .C(n_578), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_598), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_593), .B(n_574), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_591), .B(n_574), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_594), .A2(n_614), .B1(n_592), .B2(n_590), .C(n_600), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_617), .B(n_603), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_631), .B(n_615), .C(n_603), .D(n_597), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_628), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_621), .Y(n_635) );
AO22x2_ASAP7_75t_L g636 ( .A1(n_616), .A2(n_605), .B1(n_610), .B2(n_608), .Y(n_636) );
AOI221x1_ASAP7_75t_L g637 ( .A1(n_625), .A2(n_629), .B1(n_623), .B2(n_619), .C(n_624), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_622), .A2(n_615), .B(n_607), .C(n_609), .Y(n_638) );
OAI321xp33_ASAP7_75t_L g639 ( .A1(n_627), .A2(n_532), .A3(n_566), .B1(n_563), .B2(n_562), .C(n_577), .Y(n_639) );
OAI211xp5_ASAP7_75t_L g640 ( .A1(n_618), .A2(n_549), .B(n_562), .C(n_612), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_635), .B(n_626), .Y(n_641) );
NAND4xp25_ASAP7_75t_SL g642 ( .A(n_637), .B(n_630), .C(n_620), .D(n_624), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_634), .Y(n_643) );
AND4x1_ASAP7_75t_L g644 ( .A(n_638), .B(n_588), .C(n_584), .D(n_506), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_636), .A2(n_571), .B1(n_580), .B2(n_532), .Y(n_645) );
NOR3xp33_ASAP7_75t_SL g646 ( .A(n_642), .B(n_639), .C(n_633), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_643), .B(n_636), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_641), .A2(n_640), .B(n_632), .C(n_580), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_646), .B(n_644), .Y(n_649) );
XOR2xp5_ASAP7_75t_L g650 ( .A(n_647), .B(n_645), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_650), .A2(n_648), .B1(n_613), .B2(n_579), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_649), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_652), .Y(n_653) );
AOI222xp33_ASAP7_75t_SL g654 ( .A1(n_653), .A2(n_651), .B1(n_585), .B2(n_579), .C1(n_558), .C2(n_552), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_654), .A2(n_468), .B1(n_585), .B2(n_558), .Y(n_655) );
OAI32xp33_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_552), .A3(n_551), .B1(n_588), .B2(n_584), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g657 ( .A1(n_656), .A2(n_468), .B(n_506), .C(n_529), .Y(n_657) );
endmodule