module fake_ibex_2057_n_936 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_936);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_936;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_457;
wire n_357;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_158;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_580;
wire n_543;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_157;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_456;
wire n_368;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_264;
wire n_198;
wire n_164;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_159;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g157 ( 
.A(n_27),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_136),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_99),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_42),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_47),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_76),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_52),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_77),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_144),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_37),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_7),
.B(n_93),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_57),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_70),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_48),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_84),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_26),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_30),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_91),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_105),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_56),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_33),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_41),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_90),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_17),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_71),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_53),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_11),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_72),
.Y(n_202)
);

BUFx2_ASAP7_75t_SL g203 ( 
.A(n_40),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_153),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_59),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_152),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_35),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_92),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_6),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_68),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_39),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_101),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_36),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_6),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_15),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_145),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_104),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_51),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_74),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_43),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_140),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_60),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_50),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_1),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_73),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_32),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_139),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_18),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_102),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_82),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_33),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_11),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_67),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_58),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_79),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_155),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_69),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_123),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_66),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_64),
.B(n_88),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_75),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_113),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_55),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_8),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_8),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_15),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_107),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_61),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g261 ( 
.A(n_95),
.B(n_116),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_89),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_97),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_19),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_80),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_25),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_98),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_132),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_186),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_162),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_187),
.Y(n_273)
);

AND2x4_ASAP7_75t_L g274 ( 
.A(n_186),
.B(n_0),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_215),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_171),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_187),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_249),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_178),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_249),
.Y(n_282)
);

BUFx8_ASAP7_75t_L g283 ( 
.A(n_190),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_249),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_219),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_252),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_252),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_222),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_171),
.Y(n_291)
);

OAI22x1_ASAP7_75t_SL g292 ( 
.A1(n_175),
.A2(n_174),
.B1(n_267),
.B2(n_198),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_173),
.A2(n_217),
.B1(n_177),
.B2(n_241),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_187),
.B(n_214),
.Y(n_294)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_159),
.B(n_44),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_169),
.B(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_195),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_174),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_187),
.Y(n_300)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_267),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_195),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_2),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_214),
.A2(n_81),
.B(n_156),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_157),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_227),
.A2(n_78),
.B(n_154),
.Y(n_306)
);

AND2x4_ASAP7_75t_L g307 ( 
.A(n_197),
.B(n_3),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_185),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_197),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_187),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_194),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_202),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_187),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_202),
.B(n_5),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_187),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_199),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_227),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_207),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_252),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_237),
.B(n_10),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_251),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_194),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_238),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_209),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_198),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_244),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_239),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_239),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_211),
.Y(n_332)
);

AND2x4_ASAP7_75t_L g333 ( 
.A(n_259),
.B(n_12),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_213),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_257),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_220),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_266),
.B(n_165),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_322),
.Y(n_341)
);

AND2x4_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_167),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_273),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_333),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_339),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_281),
.B(n_168),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_339),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_333),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_333),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_L g354 ( 
.A(n_323),
.B(n_268),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_276),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_301),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_339),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_312),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_279),
.B(n_268),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_308),
.B(n_269),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_278),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_300),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_272),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_300),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_286),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_335),
.B(n_269),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_313),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_316),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_286),
.B(n_223),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_L g376 ( 
.A(n_296),
.B(n_256),
.C(n_234),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_312),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_335),
.B(n_293),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_307),
.B(n_172),
.Y(n_383)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_323),
.Y(n_384)
);

CKINVDCx6p67_ASAP7_75t_R g385 ( 
.A(n_295),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_307),
.B(n_158),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g388 ( 
.A1(n_303),
.A2(n_258),
.B1(n_232),
.B2(n_203),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_315),
.B(n_160),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_315),
.B(n_161),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_315),
.B(n_163),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_331),
.Y(n_393)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_271),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_323),
.B(n_295),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_274),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_277),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

OAI22xp33_ASAP7_75t_L g399 ( 
.A1(n_311),
.A2(n_175),
.B1(n_246),
.B2(n_229),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_277),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_334),
.Y(n_401)
);

OAI22xp33_ASAP7_75t_L g402 ( 
.A1(n_299),
.A2(n_229),
.B1(n_246),
.B2(n_253),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_291),
.B(n_166),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_314),
.B(n_181),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_326),
.B(n_179),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_277),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_280),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_280),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_280),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_332),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_280),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_272),
.B(n_180),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_282),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_337),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_271),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_305),
.B(n_182),
.Y(n_417)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_340),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_283),
.B(n_188),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_274),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_L g421 ( 
.A(n_338),
.B(n_176),
.C(n_183),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_324),
.Y(n_422)
);

BUFx10_ASAP7_75t_L g423 ( 
.A(n_324),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_327),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_291),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_271),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_309),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_337),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_275),
.Y(n_429)
);

INVx3_ASAP7_75t_L g430 ( 
.A(n_275),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_284),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_284),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_309),
.B(n_189),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_284),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_309),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_426),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_319),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_327),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_344),
.A2(n_336),
.B(n_319),
.C(n_294),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_321),
.C(n_319),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_417),
.B(n_336),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_342),
.B(n_336),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_342),
.A2(n_283),
.B1(n_328),
.B2(n_317),
.Y(n_444)
);

AND2x6_ASAP7_75t_SL g445 ( 
.A(n_375),
.B(n_292),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_297),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_298),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_362),
.B(n_302),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_369),
.Y(n_449)
);

A2O1A1Ixp33_ASAP7_75t_L g450 ( 
.A1(n_344),
.A2(n_294),
.B(n_304),
.C(n_306),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_350),
.B(n_193),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_405),
.B(n_200),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_352),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_204),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_416),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g456 ( 
.A(n_352),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_369),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_411),
.B(n_205),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_386),
.B(n_184),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_346),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_367),
.B(n_325),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_352),
.A2(n_325),
.B1(n_210),
.B2(n_216),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_365),
.B(n_325),
.Y(n_465)
);

A2O1A1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_353),
.A2(n_304),
.B(n_306),
.C(n_192),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_346),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_429),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_383),
.B(n_212),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_221),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_383),
.B(n_233),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_365),
.B(n_164),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_383),
.B(n_353),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_353),
.B(n_243),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_396),
.B(n_248),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_355),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_420),
.B(n_254),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_420),
.B(n_255),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_378),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_355),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_382),
.B(n_261),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_389),
.B(n_260),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_394),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g487 ( 
.A(n_402),
.B(n_231),
.C(n_201),
.Y(n_487)
);

NOR2x1p5_ASAP7_75t_L g488 ( 
.A(n_385),
.B(n_262),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

AND2x2_ASAP7_75t_SL g490 ( 
.A(n_354),
.B(n_206),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_390),
.B(n_263),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g492 ( 
.A(n_421),
.B(n_250),
.C(n_218),
.Y(n_492)
);

AO22x2_ASAP7_75t_L g493 ( 
.A1(n_391),
.A2(n_230),
.B1(n_224),
.B2(n_225),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_361),
.B(n_13),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_404),
.B(n_170),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_360),
.B(n_235),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_360),
.B(n_226),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_380),
.B(n_228),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_371),
.B(n_236),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_343),
.B(n_242),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_379),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_380),
.B(n_245),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_394),
.Y(n_503)
);

OAI221xp5_ASAP7_75t_L g504 ( 
.A1(n_388),
.A2(n_247),
.B1(n_289),
.B2(n_284),
.C(n_287),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_354),
.B(n_289),
.C(n_320),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_424),
.A2(n_289),
.B1(n_320),
.B2(n_288),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_379),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_381),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_381),
.Y(n_510)
);

BUFx4f_ASAP7_75t_L g511 ( 
.A(n_387),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_365),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_387),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_423),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_403),
.B(n_289),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_413),
.B(n_14),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_393),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.Y(n_518)
);

NOR3xp33_ASAP7_75t_L g519 ( 
.A(n_433),
.B(n_16),
.C(n_20),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_427),
.B(n_270),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_427),
.B(n_270),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_487),
.B(n_422),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_466),
.A2(n_366),
.B(n_358),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_474),
.A2(n_425),
.B(n_384),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_509),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_448),
.B(n_393),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_449),
.B(n_423),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_437),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_457),
.B(n_423),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_514),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g531 ( 
.A1(n_450),
.A2(n_456),
.B(n_453),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_511),
.B(n_457),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_366),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_444),
.B(n_422),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_368),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_448),
.B(n_443),
.Y(n_537)
);

BUFx4f_ASAP7_75t_L g538 ( 
.A(n_512),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_435),
.B(n_398),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_454),
.B(n_427),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_L g541 ( 
.A1(n_440),
.A2(n_372),
.B(n_368),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_511),
.A2(n_401),
.B1(n_409),
.B2(n_398),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_516),
.A2(n_373),
.B(n_372),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_452),
.B(n_374),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_471),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_515),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_439),
.B(n_487),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_477),
.A2(n_363),
.B(n_359),
.Y(n_549)
);

O2A1O1Ixp33_ASAP7_75t_L g550 ( 
.A1(n_441),
.A2(n_415),
.B(n_409),
.C(n_428),
.Y(n_550)
);

CKINVDCx10_ASAP7_75t_R g551 ( 
.A(n_483),
.Y(n_551)
);

NAND2x1p5_ASAP7_75t_L g552 ( 
.A(n_488),
.B(n_415),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_481),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_480),
.A2(n_370),
.B(n_364),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_463),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_459),
.A2(n_468),
.B(n_476),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_501),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_499),
.B(n_21),
.Y(n_558)
);

A2O1A1Ixp33_ASAP7_75t_L g559 ( 
.A1(n_446),
.A2(n_345),
.B(n_351),
.C(n_349),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_507),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_449),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_341),
.B(n_347),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_517),
.B(n_22),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_473),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_510),
.B(n_348),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_519),
.A2(n_357),
.B(n_432),
.C(n_431),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_513),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_518),
.Y(n_568)
);

O2A1O1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_519),
.A2(n_434),
.B(n_432),
.C(n_431),
.Y(n_569)
);

O2A1O1Ixp33_ASAP7_75t_SL g570 ( 
.A1(n_500),
.A2(n_495),
.B(n_506),
.C(n_498),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_446),
.B(n_23),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_447),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_499),
.B(n_23),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_461),
.B(n_24),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_447),
.B(n_24),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_475),
.B(n_270),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_460),
.B(n_25),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_438),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_490),
.A2(n_493),
.B1(n_461),
.B2(n_518),
.Y(n_581)
);

AND2x6_ASAP7_75t_SL g582 ( 
.A(n_483),
.B(n_26),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_469),
.A2(n_472),
.B(n_470),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_497),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_483),
.B(n_27),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_455),
.Y(n_587)
);

OAI321xp33_ASAP7_75t_L g588 ( 
.A1(n_504),
.A2(n_285),
.A3(n_287),
.B1(n_288),
.B2(n_320),
.C(n_407),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_493),
.B(n_28),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_464),
.B(n_29),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_485),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_494),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_464),
.B(n_29),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_496),
.A2(n_478),
.B1(n_482),
.B2(n_467),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_484),
.B(n_30),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_465),
.B(n_285),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_451),
.B(n_31),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g601 ( 
.A1(n_521),
.A2(n_502),
.B(n_489),
.C(n_503),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_491),
.B(n_31),
.Y(n_602)
);

NOR4xp25_ASAP7_75t_L g603 ( 
.A(n_581),
.B(n_479),
.C(n_505),
.D(n_521),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_561),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_528),
.B(n_508),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_593),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_551),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g608 ( 
.A(n_568),
.B(n_46),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_555),
.Y(n_609)
);

BUFx12f_ASAP7_75t_L g610 ( 
.A(n_582),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_546),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_584),
.A2(n_288),
.B1(n_320),
.B2(n_400),
.Y(n_612)
);

BUFx12f_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_537),
.B(n_32),
.Y(n_614)
);

AND3x4_ASAP7_75t_L g615 ( 
.A(n_576),
.B(n_34),
.C(n_35),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_564),
.Y(n_616)
);

AOI22xp5_ASAP7_75t_L g617 ( 
.A1(n_548),
.A2(n_408),
.B1(n_406),
.B2(n_397),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_525),
.Y(n_618)
);

A2O1A1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_544),
.A2(n_414),
.B(n_412),
.C(n_410),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_530),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_545),
.B(n_38),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_534),
.B(n_38),
.Y(n_622)
);

BUFx4_ASAP7_75t_SL g623 ( 
.A(n_594),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_585),
.B(n_39),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_533),
.B(n_54),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_576),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_542),
.A2(n_414),
.B1(n_410),
.B2(n_62),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_538),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_533),
.A2(n_410),
.B(n_63),
.Y(n_629)
);

O2A1O1Ixp5_ASAP7_75t_L g630 ( 
.A1(n_574),
.A2(n_558),
.B(n_598),
.C(n_575),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_526),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_547),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_553),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_572),
.B(n_532),
.Y(n_635)
);

NAND2x1p5_ASAP7_75t_L g636 ( 
.A(n_547),
.B(n_94),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_529),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_522),
.B(n_96),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

NOR2x1_ASAP7_75t_SL g640 ( 
.A(n_567),
.B(n_100),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_108),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_589),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_552),
.B(n_111),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_552),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_570),
.A2(n_549),
.B(n_554),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_579),
.B(n_112),
.Y(n_646)
);

OAI22x1_ASAP7_75t_L g647 ( 
.A1(n_591),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_535),
.A2(n_120),
.B1(n_122),
.B2(n_127),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_536),
.B(n_129),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_573),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_580),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_541),
.A2(n_133),
.B(n_134),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_L g653 ( 
.A1(n_550),
.A2(n_143),
.B(n_146),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_599),
.B(n_147),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_543),
.A2(n_524),
.B(n_565),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_539),
.Y(n_656)
);

AOI21xp33_ASAP7_75t_L g657 ( 
.A1(n_566),
.A2(n_569),
.B(n_596),
.Y(n_657)
);

AO31x2_ASAP7_75t_L g658 ( 
.A1(n_559),
.A2(n_601),
.A3(n_595),
.B(n_592),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_563),
.B(n_602),
.Y(n_659)
);

O2A1O1Ixp5_ASAP7_75t_L g660 ( 
.A1(n_540),
.A2(n_578),
.B(n_597),
.C(n_590),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_587),
.A2(n_600),
.B(n_588),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_528),
.B(n_545),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_581),
.B(n_519),
.C(n_566),
.Y(n_663)
);

AO31x2_ASAP7_75t_L g664 ( 
.A1(n_584),
.A2(n_466),
.A3(n_450),
.B(n_531),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g665 ( 
.A1(n_531),
.A2(n_466),
.B(n_450),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_538),
.Y(n_667)
);

OAI21x1_ASAP7_75t_L g668 ( 
.A1(n_523),
.A2(n_531),
.B(n_562),
.Y(n_668)
);

OAI21x1_ASAP7_75t_L g669 ( 
.A1(n_523),
.A2(n_531),
.B(n_562),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_561),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_537),
.B(n_418),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_571),
.A2(n_395),
.B(n_574),
.C(n_558),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_534),
.B(n_457),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_546),
.Y(n_674)
);

OAI22x1_ASAP7_75t_L g675 ( 
.A1(n_584),
.A2(n_324),
.B1(n_327),
.B2(n_424),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_531),
.A2(n_556),
.B(n_583),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_531),
.A2(n_556),
.B(n_583),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_546),
.Y(n_678)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_607),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_634),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_626),
.B(n_628),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_663),
.A2(n_615),
.B1(n_622),
.B2(n_627),
.Y(n_682)
);

AO31x2_ASAP7_75t_L g683 ( 
.A1(n_619),
.A2(n_642),
.A3(n_655),
.B(n_627),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_633),
.Y(n_684)
);

AO32x2_ASAP7_75t_L g685 ( 
.A1(n_631),
.A2(n_603),
.A3(n_664),
.B1(n_663),
.B2(n_658),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_605),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_616),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_639),
.B(n_666),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_650),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_674),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_678),
.Y(n_691)
);

AO21x2_ASAP7_75t_L g692 ( 
.A1(n_657),
.A2(n_629),
.B(n_608),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_609),
.B(n_675),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_673),
.B(n_611),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_609),
.B(n_644),
.Y(n_695)
);

INVx4_ASAP7_75t_L g696 ( 
.A(n_604),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_637),
.B(n_670),
.Y(n_697)
);

CKINVDCx6p67_ASAP7_75t_R g698 ( 
.A(n_613),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_624),
.Y(n_699)
);

AO31x2_ASAP7_75t_L g700 ( 
.A1(n_647),
.A2(n_625),
.A3(n_631),
.B(n_640),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_635),
.B(n_667),
.Y(n_701)
);

AO21x2_ASAP7_75t_L g702 ( 
.A1(n_608),
.A2(n_603),
.B(n_652),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_659),
.A2(n_630),
.B(n_614),
.C(n_660),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_611),
.B(n_621),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_635),
.B(n_632),
.Y(n_705)
);

INVx5_ASAP7_75t_L g706 ( 
.A(n_649),
.Y(n_706)
);

AO21x2_ASAP7_75t_L g707 ( 
.A1(n_652),
.A2(n_661),
.B(n_612),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_651),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_636),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_606),
.B(n_638),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_636),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_648),
.B(n_643),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_618),
.Y(n_713)
);

INVx6_ASAP7_75t_L g714 ( 
.A(n_610),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_606),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_623),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_641),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_620),
.Y(n_718)
);

OAI21x1_ASAP7_75t_L g719 ( 
.A1(n_617),
.A2(n_654),
.B(n_646),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_649),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_658),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_658),
.A2(n_656),
.B(n_544),
.C(n_662),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_656),
.B(n_662),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_656),
.B(n_662),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_609),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_662),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_662),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_662),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_671),
.B(n_457),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_662),
.Y(n_730)
);

CKINVDCx6p67_ASAP7_75t_R g731 ( 
.A(n_613),
.Y(n_731)
);

NOR3xp33_ASAP7_75t_L g732 ( 
.A(n_673),
.B(n_424),
.C(n_534),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_628),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_673),
.A2(n_522),
.B1(n_534),
.B2(n_385),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_662),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_662),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_626),
.A2(n_527),
.B1(n_522),
.B2(n_327),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_645),
.A2(n_677),
.A3(n_676),
.B(n_584),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_671),
.B(n_418),
.Y(n_739)
);

OAI211xp5_ASAP7_75t_L g740 ( 
.A1(n_673),
.A2(n_444),
.B(n_581),
.C(n_311),
.Y(n_740)
);

O2A1O1Ixp33_ASAP7_75t_L g741 ( 
.A1(n_671),
.A2(n_659),
.B(n_548),
.C(n_622),
.Y(n_741)
);

NAND3xp33_ASAP7_75t_L g742 ( 
.A(n_663),
.B(n_653),
.C(n_672),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_673),
.A2(n_522),
.B1(n_584),
.B2(n_534),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_609),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_656),
.A2(n_584),
.B1(n_581),
.B2(n_568),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_671),
.B(n_457),
.Y(n_746)
);

OA21x2_ASAP7_75t_L g747 ( 
.A1(n_665),
.A2(n_669),
.B(n_668),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_723),
.B(n_724),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_739),
.Y(n_749)
);

OR2x6_ASAP7_75t_L g750 ( 
.A(n_712),
.B(n_745),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_695),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_725),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_689),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_726),
.B(n_727),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_680),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_728),
.B(n_730),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_709),
.B(n_711),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_706),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_738),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_735),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_736),
.Y(n_761)
);

NOR2x1_ASAP7_75t_SL g762 ( 
.A(n_706),
.B(n_745),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_688),
.Y(n_763)
);

AOI22xp33_ASAP7_75t_L g764 ( 
.A1(n_732),
.A2(n_682),
.B1(n_743),
.B2(n_734),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_741),
.A2(n_722),
.B(n_703),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_682),
.B(n_712),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_747),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_691),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_740),
.A2(n_742),
.B(n_719),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_733),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_729),
.B(n_746),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_743),
.A2(n_737),
.B1(n_699),
.B2(n_717),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_708),
.Y(n_773)
);

INVx4_ASAP7_75t_L g774 ( 
.A(n_706),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_720),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_740),
.B(n_694),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_684),
.B(n_690),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_744),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_733),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_721),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_687),
.B(n_686),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_715),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_705),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_701),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_696),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_696),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_698),
.Y(n_787)
);

BUFx2_ASAP7_75t_SL g788 ( 
.A(n_701),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_693),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_718),
.Y(n_790)
);

INVxp67_ASAP7_75t_L g791 ( 
.A(n_697),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_710),
.A2(n_686),
.B1(n_681),
.B2(n_707),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_685),
.B(n_704),
.Y(n_793)
);

BUFx2_ASAP7_75t_SL g794 ( 
.A(n_716),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_685),
.B(n_704),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_685),
.B(n_713),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_683),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_683),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_700),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_702),
.B(n_692),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_755),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_753),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_768),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_780),
.Y(n_804)
);

BUFx3_ASAP7_75t_L g805 ( 
.A(n_779),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_793),
.B(n_692),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_793),
.B(n_714),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_779),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_764),
.A2(n_714),
.B1(n_731),
.B2(n_679),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_795),
.B(n_750),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_776),
.B(n_778),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_750),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_789),
.B(n_772),
.C(n_765),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_748),
.Y(n_814)
);

BUFx3_ASAP7_75t_L g815 ( 
.A(n_779),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_770),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_775),
.B(n_750),
.Y(n_817)
);

NAND2x1p5_ASAP7_75t_L g818 ( 
.A(n_774),
.B(n_758),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_796),
.B(n_754),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_762),
.B(n_799),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_773),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_796),
.B(n_769),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_770),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_786),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_760),
.B(n_761),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_767),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_785),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_777),
.B(n_763),
.Y(n_828)
);

AND2x4_ASAP7_75t_SL g829 ( 
.A(n_774),
.B(n_785),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_752),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_797),
.B(n_798),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_751),
.B(n_790),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_756),
.B(n_783),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_790),
.B(n_781),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_782),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_819),
.B(n_822),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_819),
.B(n_797),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_829),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_822),
.B(n_800),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_801),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_802),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_826),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_814),
.B(n_771),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_810),
.B(n_800),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_810),
.B(n_759),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_817),
.B(n_762),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_828),
.B(n_749),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_811),
.B(n_766),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_803),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_805),
.B(n_792),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_821),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_835),
.Y(n_852)
);

NAND4xp25_ASAP7_75t_L g853 ( 
.A(n_813),
.B(n_791),
.C(n_787),
.D(n_784),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_824),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_825),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_809),
.B(n_794),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_805),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_804),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_842),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_854),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_836),
.B(n_806),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_846),
.B(n_820),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_836),
.B(n_830),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_853),
.A2(n_812),
.B1(n_807),
.B2(n_817),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_843),
.B(n_794),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_857),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_858),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_855),
.B(n_807),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_839),
.B(n_812),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_839),
.B(n_831),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_837),
.B(n_832),
.Y(n_871)
);

OR3x2_ASAP7_75t_L g872 ( 
.A(n_848),
.B(n_832),
.C(n_834),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_844),
.B(n_831),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_870),
.B(n_837),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_R g875 ( 
.A(n_862),
.B(n_808),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_870),
.B(n_840),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_866),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_860),
.B(n_863),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_859),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_861),
.B(n_841),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_861),
.B(n_844),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_867),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_873),
.B(n_845),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_866),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_862),
.B(n_846),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_873),
.B(n_871),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_874),
.B(n_868),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_883),
.B(n_881),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_876),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_884),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_884),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_885),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_877),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_SL g894 ( 
.A1(n_875),
.A2(n_838),
.B(n_865),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_880),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_883),
.B(n_869),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_885),
.A2(n_815),
.B(n_862),
.C(n_878),
.Y(n_897)
);

AOI222xp33_ASAP7_75t_L g898 ( 
.A1(n_881),
.A2(n_847),
.B1(n_869),
.B2(n_856),
.C1(n_833),
.C2(n_852),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_894),
.A2(n_885),
.B(n_815),
.C(n_862),
.Y(n_899)
);

OA21x2_ASAP7_75t_L g900 ( 
.A1(n_894),
.A2(n_879),
.B(n_882),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_889),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_895),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_898),
.B(n_886),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_892),
.Y(n_904)
);

OAI21xp33_ASAP7_75t_SL g905 ( 
.A1(n_903),
.A2(n_890),
.B(n_888),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_901),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_899),
.B(n_897),
.Y(n_907)
);

AOI21xp33_ASAP7_75t_L g908 ( 
.A1(n_905),
.A2(n_900),
.B(n_902),
.Y(n_908)
);

OR2x2_ASAP7_75t_L g909 ( 
.A(n_906),
.B(n_904),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_909),
.Y(n_910)
);

NAND4xp25_ASAP7_75t_L g911 ( 
.A(n_908),
.B(n_907),
.C(n_899),
.D(n_864),
.Y(n_911)
);

NOR2x1_ASAP7_75t_L g912 ( 
.A(n_911),
.B(n_900),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_910),
.B(n_891),
.C(n_904),
.Y(n_913)
);

XNOR2xp5_ASAP7_75t_L g914 ( 
.A(n_912),
.B(n_900),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_913),
.B(n_893),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_915),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_915),
.Y(n_917)
);

NOR2x1_ASAP7_75t_L g918 ( 
.A(n_914),
.B(n_892),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_916),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_918),
.B(n_877),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_917),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_917),
.A2(n_808),
.B1(n_857),
.B2(n_887),
.Y(n_922)
);

NOR2x1p5_ASAP7_75t_L g923 ( 
.A(n_916),
.B(n_896),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_919),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_921),
.B(n_849),
.Y(n_925)
);

AOI22x1_ASAP7_75t_L g926 ( 
.A1(n_923),
.A2(n_758),
.B1(n_818),
.B2(n_788),
.Y(n_926)
);

XNOR2x1_ASAP7_75t_L g927 ( 
.A(n_922),
.B(n_757),
.Y(n_927)
);

OA22x2_ASAP7_75t_L g928 ( 
.A1(n_920),
.A2(n_829),
.B1(n_850),
.B2(n_823),
.Y(n_928)
);

AOI22xp5_ASAP7_75t_L g929 ( 
.A1(n_919),
.A2(n_872),
.B1(n_757),
.B2(n_788),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_924),
.A2(n_827),
.B1(n_816),
.B2(n_823),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_927),
.B(n_851),
.Y(n_931)
);

AOI21xp33_ASAP7_75t_SL g932 ( 
.A1(n_928),
.A2(n_818),
.B(n_757),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_930),
.B(n_925),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_933),
.B(n_926),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_934),
.B(n_932),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_935),
.A2(n_931),
.B1(n_929),
.B2(n_872),
.Y(n_936)
);


endmodule