module fake_jpeg_16583_n_122 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_SL g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_0),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_16),
.B1(n_21),
.B2(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_14),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_14),
.Y(n_47)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_40),
.A2(n_44),
.B1(n_50),
.B2(n_18),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_29),
.B(n_18),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_17),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_16),
.B1(n_19),
.B2(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_35),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_53),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_33),
.C(n_32),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_24),
.C(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_33),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_36),
.B1(n_34),
.B2(n_23),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_59),
.B1(n_65),
.B2(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_19),
.B1(n_25),
.B2(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_17),
.B1(n_20),
.B2(n_28),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_69),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_76),
.Y(n_82)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_38),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_78),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_87),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_64),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_72),
.C(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_51),
.Y(n_87)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_56),
.B1(n_39),
.B2(n_38),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_74),
.B1(n_54),
.B2(n_70),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_42),
.B(n_63),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_89),
.A2(n_75),
.B(n_43),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_71),
.A2(n_64),
.B1(n_65),
.B2(n_60),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_90),
.A2(n_61),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_82),
.C(n_83),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_42),
.B(n_61),
.Y(n_94)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_66),
.B1(n_24),
.B2(n_27),
.C(n_12),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_85),
.C(n_46),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_79),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_104),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_88),
.B1(n_82),
.B2(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_105),
.B1(n_94),
.B2(n_91),
.Y(n_106)
);

FAx1_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_90),
.CI(n_88),
.CON(n_104),
.SN(n_104)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_110),
.C(n_111),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_92),
.C(n_98),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_107),
.A2(n_108),
.B1(n_2),
.B2(n_3),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_102),
.B1(n_101),
.B2(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_84),
.C(n_27),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_115),
.C(n_113),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_109),
.A2(n_9),
.B1(n_11),
.B2(n_6),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_116),
.B(n_117),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_107),
.C(n_4),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_120),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g122 ( 
.A(n_121),
.Y(n_122)
);


endmodule