module real_jpeg_12754_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_3),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_3),
.A2(n_54),
.B1(n_57),
.B2(n_63),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_3),
.A2(n_30),
.B1(n_36),
.B2(n_63),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_59),
.B1(n_60),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_4),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_4),
.A2(n_54),
.B1(n_57),
.B2(n_119),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_119),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_4),
.A2(n_30),
.B1(n_36),
.B2(n_119),
.Y(n_257)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_54),
.B1(n_57),
.B2(n_182),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_6),
.A2(n_41),
.B1(n_42),
.B2(n_182),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_6),
.A2(n_30),
.B1(n_36),
.B2(n_182),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_7),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_7),
.A2(n_54),
.B1(n_57),
.B2(n_65),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_65),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_7),
.A2(n_30),
.B1(n_36),
.B2(n_65),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_8),
.A2(n_54),
.B1(n_57),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_8),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_73),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_8),
.A2(n_41),
.B1(n_42),
.B2(n_73),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_8),
.A2(n_30),
.B1(n_36),
.B2(n_73),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_30),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_9),
.A2(n_35),
.B1(n_54),
.B2(n_57),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_9),
.A2(n_35),
.B1(n_59),
.B2(n_60),
.Y(n_325)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_11),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_13),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_13),
.A2(n_54),
.B1(n_57),
.B2(n_155),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_155),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_13),
.A2(n_30),
.B1(n_36),
.B2(n_155),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_14),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g194 ( 
.A1(n_14),
.A2(n_59),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_185),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_14),
.B(n_57),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_174),
.Y(n_247)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_42),
.B(n_45),
.C(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_14),
.B(n_81),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_14),
.B(n_33),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_14),
.B(n_50),
.Y(n_274)
);

AOI21xp33_ASAP7_75t_L g283 ( 
.A1(n_14),
.A2(n_57),
.B(n_233),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_15),
.A2(n_49),
.B1(n_54),
.B2(n_57),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_15),
.A2(n_30),
.B1(n_36),
.B2(n_49),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_15),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_16),
.A2(n_40),
.B1(n_54),
.B2(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_16),
.A2(n_40),
.B1(n_59),
.B2(n_60),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_16),
.A2(n_30),
.B1(n_36),
.B2(n_40),
.Y(n_146)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_321),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_308),
.B(n_320),
.Y(n_19)
);

AO21x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_133),
.B(n_305),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_120),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_96),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_23),
.B(n_96),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_66),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_82),
.C(n_94),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_51),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_25),
.A2(n_26),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_27),
.A2(n_28),
.B1(n_51),
.B2(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_27),
.A2(n_28),
.B1(n_37),
.B2(n_38),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_34),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_33),
.B1(n_34),
.B2(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_29),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_29),
.A2(n_33),
.B1(n_146),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_29),
.A2(n_33),
.B1(n_170),
.B2(n_212),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_29),
.A2(n_33),
.B1(n_212),
.B2(n_236),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_29),
.A2(n_33),
.B1(n_236),
.B2(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_29),
.A2(n_33),
.B1(n_174),
.B2(n_269),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_29),
.A2(n_33),
.B1(n_262),
.B2(n_269),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_30),
.B(n_271),
.Y(n_270)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_32),
.A2(n_110),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_32),
.A2(n_144),
.B1(n_261),
.B2(n_263),
.Y(n_260)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_36),
.A2(n_46),
.B(n_174),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_39),
.A2(n_43),
.B1(n_50),
.B2(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_41),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_41),
.A2(n_42),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_41),
.A2(n_57),
.A3(n_78),
.B1(n_232),
.B2(n_234),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_42),
.B(n_77),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_43),
.A2(n_50),
.B(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_43),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_43),
.A2(n_50),
.B1(n_149),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_43),
.A2(n_50),
.B1(n_200),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_43),
.A2(n_50),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_43),
.A2(n_50),
.B1(n_248),
.B2(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_47),
.A2(n_114),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_47),
.A2(n_150),
.B1(n_227),
.B2(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_51),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_64),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_52),
.A2(n_53),
.B1(n_85),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_52),
.A2(n_53),
.B1(n_118),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_52),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_52),
.A2(n_53),
.B1(n_181),
.B2(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_53),
.Y(n_185)
);

OA22x2_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_57),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g171 ( 
.A1(n_54),
.A2(n_56),
.A3(n_59),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_55),
.B(n_57),
.Y(n_172)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_60),
.B(n_174),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_82),
.B1(n_94),
.B2(n_95),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_68),
.B(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_72),
.A2(n_75),
.B1(n_76),
.B2(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_80),
.B1(n_81),
.B2(n_91),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_74),
.A2(n_81),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_74),
.A2(n_81),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_74),
.A2(n_81),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_76),
.B1(n_92),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_75),
.A2(n_76),
.B1(n_116),
.B2(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_75),
.A2(n_76),
.B1(n_177),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_75),
.A2(n_76),
.B1(n_208),
.B2(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_76),
.Y(n_81)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_83),
.A2(n_84),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_88),
.C(n_90),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_84),
.B(n_123),
.C(n_126),
.Y(n_309)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_93),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_88),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_93),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_88),
.B(n_129),
.C(n_131),
.Y(n_319)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_102),
.C(n_104),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_97),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_157)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.C(n_117),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_106),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_117),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_120),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_121),
.B(n_122),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_130),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_132),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_158),
.B(n_304),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_156),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_135),
.B(n_156),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_140),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_151),
.C(n_153),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_142),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_143),
.B(n_147),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_153),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_188),
.B(n_303),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_186),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_160),
.B(n_186),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_165),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_166),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_175),
.C(n_179),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_168),
.A2(n_169),
.B1(n_171),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_171),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_173),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_179),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_183),
.A2(n_185),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_183),
.A2(n_185),
.B1(n_316),
.B2(n_325),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_219),
.B(n_297),
.C(n_302),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_213),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_190),
.B(n_213),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_203),
.C(n_205),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_191),
.A2(n_192),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_193),
.B(n_197),
.C(n_202),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_203),
.B(n_205),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_206),
.B(n_224),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_211),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_215),
.B(n_216),
.C(n_217),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_296),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_240),
.B(n_295),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_237),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_222),
.B(n_237),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_223),
.B(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_225),
.A2(n_228),
.B1(n_229),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_225),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_230),
.A2(n_231),
.B1(n_235),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_238),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_289),
.B(n_294),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_278),
.B(n_288),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_258),
.B(n_277),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_251),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_244),
.B(n_251),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_256),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_254),
.C(n_256),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_266),
.B(n_276),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_260),
.B(n_264),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_272),
.B(n_275),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_273),
.B(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_286),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_284),
.C(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_299),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_319),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_328),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_326),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);


endmodule