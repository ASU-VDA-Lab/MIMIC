module fake_jpeg_22995_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_152;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_19),
.B(n_2),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_38),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_30),
.B1(n_34),
.B2(n_21),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_55),
.Y(n_88)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_63),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_66),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_65),
.B(n_74),
.Y(n_118)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_69),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_75),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_41),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_71),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_30),
.B1(n_21),
.B2(n_27),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_45),
.A2(n_30),
.B1(n_21),
.B2(n_27),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_44),
.A2(n_34),
.B1(n_22),
.B2(n_18),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_34),
.B1(n_22),
.B2(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_35),
.B1(n_22),
.B2(n_18),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_35),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_85),
.B(n_104),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_87),
.Y(n_124)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_92),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_78),
.B(n_72),
.C(n_35),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_7),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_33),
.B1(n_37),
.B2(n_36),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_59),
.B(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_97),
.B(n_24),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_66),
.B(n_23),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_67),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_3),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_23),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_113),
.Y(n_134)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_7),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_54),
.A2(n_26),
.B1(n_37),
.B2(n_36),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_111),
.A2(n_115),
.B1(n_24),
.B2(n_23),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_59),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_58),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_56),
.A2(n_31),
.B(n_29),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_28),
.B(n_25),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_56),
.B1(n_28),
.B2(n_25),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_120),
.A2(n_150),
.B1(n_112),
.B2(n_93),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_121),
.A2(n_129),
.B(n_142),
.Y(n_173)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_123),
.Y(n_158)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_130),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_131),
.B1(n_132),
.B2(n_136),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_128),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_103),
.A2(n_76),
.B(n_23),
.C(n_5),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_96),
.A2(n_23),
.B1(n_17),
.B2(n_7),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_114),
.B1(n_98),
.B2(n_116),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_85),
.B(n_3),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_145),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_4),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_148),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_9),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_118),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_88),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_17),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_104),
.B(n_115),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_115),
.B1(n_95),
.B2(n_89),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_9),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_151),
.A2(n_99),
.B1(n_107),
.B2(n_100),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_153),
.A2(n_156),
.B1(n_167),
.B2(n_170),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_100),
.B1(n_108),
.B2(n_95),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_159),
.B(n_165),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g163 ( 
.A1(n_129),
.A2(n_101),
.B(n_109),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_163),
.A2(n_14),
.B(n_15),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_130),
.A2(n_102),
.B1(n_101),
.B2(n_83),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_86),
.B(n_94),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_169),
.A2(n_180),
.B(n_127),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_142),
.A2(n_119),
.B1(n_145),
.B2(n_137),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_119),
.A2(n_83),
.B1(n_106),
.B2(n_93),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_175),
.B1(n_183),
.B2(n_143),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_86),
.C(n_94),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_140),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_174),
.B(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_133),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_9),
.B(n_11),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_181),
.A2(n_135),
.B(n_147),
.Y(n_198)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_121),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_184),
.A2(n_191),
.B1(n_195),
.B2(n_206),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_139),
.Y(n_187)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_187),
.A2(n_194),
.B(n_176),
.Y(n_221)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_188),
.B(n_190),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_138),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_192),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_160),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_140),
.B1(n_126),
.B2(n_143),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_162),
.B(n_166),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_196),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_167),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_177),
.B1(n_173),
.B2(n_174),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_160),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_199),
.B(n_209),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_123),
.B(n_135),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_184),
.Y(n_223)
);

OA21x2_ASAP7_75t_SL g201 ( 
.A1(n_168),
.A2(n_11),
.B(n_12),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_201),
.B(n_181),
.Y(n_213)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_164),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_208)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_208),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_213),
.A2(n_233),
.B(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_159),
.Y(n_214)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

AOI22x1_ASAP7_75t_L g215 ( 
.A1(n_201),
.A2(n_163),
.B1(n_154),
.B2(n_177),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_221),
.B(n_185),
.C(n_194),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_155),
.C(n_170),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_222),
.C(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_217),
.B(n_227),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_186),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_219),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_187),
.C(n_202),
.Y(n_222)
);

INVx13_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_226),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_210),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_229),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_231),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_163),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_211),
.B(n_205),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_189),
.B(n_161),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_193),
.B1(n_203),
.B2(n_207),
.Y(n_235)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_202),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_244),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_240),
.C(n_242),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_194),
.B1(n_211),
.B2(n_206),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_187),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_216),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_212),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_247),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_198),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_209),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_224),
.C(n_228),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_227),
.B(n_215),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_260),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_214),
.C(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_237),
.C(n_235),
.Y(n_274)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_257),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_249),
.B(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_226),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_264),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_215),
.B(n_231),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_266),
.B1(n_218),
.B2(n_246),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

NAND4xp25_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_231),
.C(n_213),
.D(n_205),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_268),
.B(n_243),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_236),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_271),
.C(n_274),
.Y(n_283)
);

INVx11_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_243),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_277),
.B(n_265),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_280),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_262),
.B(n_247),
.Y(n_280)
);

NOR4xp25_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_262),
.C(n_266),
.D(n_261),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_281),
.A2(n_288),
.B(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_258),
.C(n_255),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_257),
.C(n_254),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_258),
.C(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_287),
.C(n_152),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_267),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_289),
.A2(n_284),
.B(n_283),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_285),
.A2(n_279),
.B1(n_254),
.B2(n_270),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_282),
.B(n_272),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_284),
.B(n_287),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_285),
.A2(n_218),
.B1(n_267),
.B2(n_244),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_294),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_16),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_297),
.A2(n_292),
.A3(n_268),
.B1(n_219),
.B2(n_152),
.C1(n_179),
.C2(n_180),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_295),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_182),
.C1(n_208),
.C2(n_298),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_301),
.B(n_16),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_302),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_305),
.Y(n_306)
);


endmodule