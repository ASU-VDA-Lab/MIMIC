module fake_jpeg_15566_n_137 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx2_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_5),
.Y(n_17)
);

HB1xp67_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_29),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_21),
.B1(n_15),
.B2(n_16),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_33),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_22),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

AOI32xp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_16),
.A3(n_28),
.B1(n_17),
.B2(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_13),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_24),
.B1(n_29),
.B2(n_12),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_29),
.B1(n_24),
.B2(n_20),
.Y(n_53)
);

OAI32xp33_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_14),
.A3(n_17),
.B1(n_27),
.B2(n_19),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_59),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_24),
.B1(n_30),
.B2(n_31),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_39),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_19),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_13),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_68),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_76),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_11),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_30),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_11),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_30),
.Y(n_93)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_58),
.B1(n_57),
.B2(n_51),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_79),
.B1(n_3),
.B2(n_4),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_27),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_86),
.C(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_70),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_90),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_27),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_94),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_75),
.B(n_68),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_96),
.B(n_98),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_76),
.C(n_65),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_101),
.C(n_102),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_75),
.B(n_65),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_64),
.C(n_66),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_63),
.C(n_69),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_103),
.B(n_84),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_105),
.A2(n_87),
.B1(n_82),
.B2(n_91),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_85),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_112),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_97),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g124 ( 
.A(n_116),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_89),
.B(n_97),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_98),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_114),
.A2(n_82),
.B1(n_94),
.B2(n_103),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_119),
.A2(n_95),
.B1(n_80),
.B2(n_79),
.Y(n_123)
);

AOI31xp67_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_111),
.A3(n_95),
.B(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_122),
.B(n_123),
.C(n_119),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_8),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_8),
.B(n_9),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_120),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_129),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_9),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_131),
.B(n_2),
.Y(n_135)
);

NOR2xp67_ASAP7_75t_SL g132 ( 
.A(n_127),
.B(n_11),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_132),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_134),
.Y(n_137)
);


endmodule