module fake_netlist_1_11188_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_13;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g10 ( .A(n_4), .B(n_9), .Y(n_10) );
BUFx6f_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_7), .A2(n_3), .B1(n_0), .B2(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
OR2x6_ASAP7_75t_L g16 ( .A(n_15), .B(n_0), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_12), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_11), .Y(n_19) );
OR2x6_ASAP7_75t_L g20 ( .A(n_16), .B(n_10), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_16), .Y(n_23) );
AOI211x1_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_10), .B(n_19), .C(n_16), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_23), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_18), .Y(n_29) );
AOI21xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_22), .B(n_17), .Y(n_30) );
CKINVDCx16_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
CKINVDCx20_ASAP7_75t_R g32 ( .A(n_28), .Y(n_32) );
XNOR2x1_ASAP7_75t_L g33 ( .A(n_30), .B(n_13), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
AOI21xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_24), .B(n_11), .Y(n_35) );
AOI22xp5_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_31), .B1(n_33), .B2(n_11), .Y(n_36) );
OA331x2_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_34), .A3(n_2), .B1(n_3), .B2(n_5), .B3(n_1), .C1(n_8), .Y(n_37) );
endmodule