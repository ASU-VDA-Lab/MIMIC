module fake_jpeg_30104_n_489 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_489);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_489;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_434;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_419;
wire n_133;
wire n_378;
wire n_132;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_361;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_11),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_7),
.B(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_5),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_48),
.B(n_50),
.Y(n_129)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_51),
.B(n_54),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_24),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_55),
.B(n_59),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_63),
.Y(n_120)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_64),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_65),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g117 ( 
.A(n_68),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_14),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_79),
.Y(n_139)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_85),
.Y(n_146)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_21),
.B(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_90),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_86),
.B(n_87),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_16),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_95),
.Y(n_115)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_46),
.B1(n_26),
.B2(n_43),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_41),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_41),
.B1(n_45),
.B2(n_30),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_100),
.A2(n_111),
.B1(n_125),
.B2(n_134),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_31),
.B1(n_38),
.B2(n_44),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_104),
.A2(n_106),
.B1(n_113),
.B2(n_135),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_76),
.A2(n_40),
.B1(n_23),
.B2(n_42),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_57),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_112),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_81),
.B1(n_57),
.B2(n_69),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_68),
.A2(n_31),
.B(n_44),
.C(n_43),
.Y(n_114)
);

NOR2x1_ASAP7_75t_L g182 ( 
.A(n_114),
.B(n_17),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_68),
.A2(n_46),
.B1(n_26),
.B2(n_39),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_118),
.A2(n_124),
.B1(n_143),
.B2(n_145),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_63),
.A2(n_46),
.B1(n_26),
.B2(n_39),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_62),
.A2(n_30),
.B1(n_32),
.B2(n_27),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_91),
.A2(n_27),
.B(n_32),
.C(n_42),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_53),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_90),
.B(n_23),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_0),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_82),
.A2(n_34),
.B1(n_19),
.B2(n_26),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_93),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_70),
.A2(n_34),
.B1(n_26),
.B2(n_46),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_65),
.A2(n_85),
.B1(n_80),
.B2(n_77),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_136),
.A2(n_142),
.B1(n_88),
.B2(n_72),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_46),
.B1(n_17),
.B2(n_13),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_58),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_92),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_126),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_151),
.B(n_155),
.Y(n_230)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_121),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_153),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_156),
.B(n_161),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_183),
.B1(n_195),
.B2(n_159),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_159),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_97),
.B(n_9),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_160),
.B(n_171),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_121),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_162),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_168),
.Y(n_223)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_129),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_170),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_49),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_97),
.B(n_8),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_172),
.Y(n_226)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

INVx13_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_106),
.A2(n_61),
.B1(n_83),
.B2(n_64),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_179),
.B1(n_190),
.B2(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_184),
.Y(n_212)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_178),
.Y(n_203)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_114),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_115),
.C(n_113),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_188),
.C(n_98),
.Y(n_224)
);

OR2x4_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_193),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_116),
.A2(n_89),
.B1(n_60),
.B2(n_56),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_116),
.B(n_111),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_60),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_186),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_56),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_146),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_191),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_17),
.C(n_10),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_119),
.B(n_10),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_189),
.B(n_196),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_137),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

BUFx8_ASAP7_75t_L g192 ( 
.A(n_109),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_192),
.Y(n_200)
);

NAND2x1_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_149),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_120),
.B(n_0),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_120),
.B(n_0),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_99),
.B(n_1),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_198),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_99),
.B(n_1),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_103),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_204),
.B(n_227),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_211),
.Y(n_254)
);

CKINVDCx12_ASAP7_75t_R g207 ( 
.A(n_153),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_179),
.A2(n_136),
.B(n_109),
.C(n_150),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_208),
.A2(n_195),
.B(n_183),
.Y(n_251)
);

NOR2x1p5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_150),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_155),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_144),
.B1(n_138),
.B2(n_139),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_216),
.A2(n_176),
.B1(n_172),
.B2(n_166),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_180),
.A2(n_102),
.B1(n_109),
.B2(n_149),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_220),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_188),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_181),
.B(n_122),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g229 ( 
.A(n_182),
.B(n_122),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_229),
.B(n_185),
.Y(n_256)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_157),
.A2(n_139),
.B1(n_138),
.B2(n_137),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_237),
.B1(n_175),
.B2(n_154),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_151),
.A2(n_107),
.B1(n_108),
.B2(n_123),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_167),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_153),
.Y(n_248)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_169),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_240),
.B(n_246),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_215),
.A2(n_180),
.B1(n_159),
.B2(n_193),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_184),
.C(n_170),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_265),
.C(n_235),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_244),
.A2(n_251),
.B(n_256),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_245),
.B(n_257),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_247),
.Y(n_285)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_248),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_249),
.A2(n_250),
.B1(n_266),
.B2(n_208),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_211),
.A2(n_154),
.B1(n_177),
.B2(n_193),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_171),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_259),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_202),
.B(n_187),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_260),
.A2(n_268),
.B1(n_271),
.B2(n_208),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_194),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_262),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_168),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_221),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_263),
.Y(n_306)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_215),
.A2(n_186),
.B(n_197),
.C(n_198),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_264),
.A2(n_273),
.B(n_228),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_230),
.B1(n_212),
.B2(n_233),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_206),
.A2(n_158),
.B1(n_190),
.B2(n_123),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_269),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_163),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_272),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_206),
.A2(n_158),
.B1(n_190),
.B2(n_123),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_205),
.B(n_189),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_225),
.A2(n_196),
.B(n_190),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_173),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_274),
.B(n_200),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_231),
.B(n_173),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_200),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_205),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_276),
.B(n_292),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_250),
.A2(n_206),
.B1(n_235),
.B2(n_204),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_279),
.A2(n_291),
.B1(n_296),
.B2(n_310),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_293),
.C(n_243),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_268),
.A2(n_229),
.B1(n_227),
.B2(n_237),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_262),
.B(n_214),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_287),
.B(n_261),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_208),
.B1(n_232),
.B2(n_222),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_289),
.A2(n_290),
.B1(n_254),
.B2(n_249),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_218),
.Y(n_293)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_295),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_254),
.A2(n_216),
.B1(n_208),
.B2(n_214),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_268),
.A2(n_218),
.B1(n_228),
.B2(n_190),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_301),
.B(n_303),
.Y(n_330)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_248),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_244),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_244),
.A2(n_199),
.B(n_213),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_241),
.B(n_274),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_254),
.A2(n_222),
.B1(n_174),
.B2(n_213),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_311),
.B(n_326),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_313),
.A2(n_296),
.B1(n_310),
.B2(n_279),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_265),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_319),
.C(n_293),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_SL g318 ( 
.A(n_283),
.B(n_256),
.C(n_292),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_318),
.A2(n_325),
.B(n_264),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_272),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_278),
.Y(n_357)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_300),
.Y(n_321)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_321),
.Y(n_352)
);

OR2x2_ASAP7_75t_L g363 ( 
.A(n_323),
.B(n_274),
.Y(n_363)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_300),
.Y(n_324)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_271),
.B1(n_255),
.B2(n_244),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_255),
.B(n_274),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_327),
.A2(n_331),
.B(n_343),
.Y(n_366)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_302),
.Y(n_328)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_283),
.A2(n_258),
.B(n_266),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_332),
.Y(n_349)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_333),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_288),
.A2(n_306),
.B1(n_253),
.B2(n_289),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_334),
.A2(n_310),
.B1(n_291),
.B2(n_298),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_282),
.B(n_259),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_335),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_278),
.B(n_272),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_340),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_288),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_338),
.Y(n_346)
);

NOR4xp25_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_281),
.C(n_294),
.D(n_246),
.Y(n_351)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_282),
.B(n_264),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_341),
.B(n_273),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_287),
.B(n_275),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_342),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_303),
.B(n_271),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_345),
.C(n_354),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_293),
.C(n_276),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_347),
.A2(n_350),
.B1(n_343),
.B2(n_337),
.Y(n_376)
);

OA21x2_ASAP7_75t_SL g384 ( 
.A1(n_351),
.A2(n_362),
.B(n_341),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_319),
.B(n_276),
.C(n_286),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_355),
.B(n_374),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_357),
.B(n_370),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_313),
.A2(n_290),
.B1(n_281),
.B2(n_294),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_361),
.A2(n_329),
.B1(n_251),
.B2(n_333),
.Y(n_386)
);

NOR3xp33_ASAP7_75t_SL g362 ( 
.A(n_318),
.B(n_246),
.C(n_252),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_372),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_339),
.A2(n_306),
.B1(n_260),
.B2(n_301),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_364),
.A2(n_369),
.B1(n_363),
.B2(n_360),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_240),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_365),
.B(n_368),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_317),
.B(n_240),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_342),
.A2(n_260),
.B1(n_299),
.B2(n_285),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_252),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_327),
.B(n_273),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_373),
.C(n_329),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_314),
.B(n_331),
.C(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_376),
.A2(n_386),
.B1(n_396),
.B2(n_346),
.Y(n_410)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_352),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_381),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_366),
.A2(n_314),
.B(n_325),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_379),
.A2(n_382),
.B(n_397),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_348),
.A2(n_330),
.B1(n_311),
.B2(n_326),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_392),
.B1(n_358),
.B2(n_367),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_353),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_366),
.A2(n_337),
.B(n_343),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g403 ( 
.A(n_384),
.B(n_362),
.CI(n_365),
.CON(n_403),
.SN(n_403)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_353),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_385),
.A2(n_399),
.B1(n_400),
.B2(n_349),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_387),
.B(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_344),
.B(n_336),
.C(n_309),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_394),
.C(n_354),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_297),
.B(n_328),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_390),
.B(n_322),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_355),
.B(n_251),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_340),
.C(n_324),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_350),
.A2(n_321),
.B1(n_315),
.B2(n_312),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_373),
.A2(n_315),
.B(n_312),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_371),
.A2(n_299),
.B(n_285),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_356),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_411),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_394),
.B(n_370),
.C(n_357),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_414),
.C(n_417),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_404),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_387),
.B(n_360),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_408),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_395),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_418),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_376),
.B1(n_396),
.B2(n_398),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_368),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_359),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_413),
.B(n_415),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_361),
.C(n_367),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_349),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_416),
.A2(n_421),
.B1(n_390),
.B2(n_253),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_284),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_284),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_419),
.A2(n_375),
.B(n_385),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_253),
.B1(n_247),
.B2(n_267),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_403),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_424),
.Y(n_443)
);

AOI211xp5_ASAP7_75t_SL g423 ( 
.A1(n_405),
.A2(n_393),
.B(n_378),
.C(n_386),
.Y(n_423)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_423),
.Y(n_449)
);

BUFx4f_ASAP7_75t_SL g424 ( 
.A(n_408),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_403),
.B(n_242),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_425),
.B(n_429),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_426),
.A2(n_263),
.B1(n_245),
.B2(n_209),
.Y(n_451)
);

OAI221xp5_ASAP7_75t_L g427 ( 
.A1(n_416),
.A2(n_397),
.B1(n_378),
.B2(n_379),
.C(n_405),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_427),
.B(n_428),
.Y(n_445)
);

OAI221xp5_ASAP7_75t_L g428 ( 
.A1(n_412),
.A2(n_400),
.B1(n_399),
.B2(n_377),
.C(n_381),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_433),
.B(n_410),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_414),
.B(n_391),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_437),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_401),
.B(n_389),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_439),
.B(n_451),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_431),
.A2(n_417),
.B1(n_421),
.B2(n_418),
.Y(n_440)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_440),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_426),
.A2(n_407),
.B(n_420),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_201),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_432),
.A2(n_407),
.B(n_411),
.Y(n_444)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_444),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_402),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_446),
.B(n_452),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_429),
.B(n_420),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_438),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_430),
.A2(n_238),
.B(n_257),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_450),
.A2(n_424),
.B(n_192),
.Y(n_456)
);

OAI221xp5_ASAP7_75t_L g452 ( 
.A1(n_423),
.A2(n_210),
.B1(n_201),
.B2(n_209),
.C(n_219),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_436),
.A2(n_210),
.B1(n_219),
.B2(n_203),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_453),
.B(n_451),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_203),
.C(n_178),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_164),
.C(n_152),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_455),
.A2(n_140),
.B1(n_148),
.B2(n_96),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_456),
.B(n_460),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_464),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_441),
.B(n_434),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_446),
.B(n_424),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_462),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_443),
.B(n_162),
.Y(n_462)
);

AOI322xp5_ASAP7_75t_L g468 ( 
.A1(n_466),
.A2(n_445),
.A3(n_449),
.B1(n_448),
.B2(n_442),
.C1(n_447),
.C2(n_122),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_107),
.C(n_165),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_128),
.C(n_132),
.Y(n_474)
);

AOI322xp5_ASAP7_75t_L g480 ( 
.A1(n_468),
.A2(n_466),
.A3(n_467),
.B1(n_459),
.B2(n_7),
.C1(n_4),
.C2(n_6),
.Y(n_480)
);

AOI322xp5_ASAP7_75t_L g470 ( 
.A1(n_465),
.A2(n_440),
.A3(n_454),
.B1(n_148),
.B2(n_109),
.C1(n_140),
.C2(n_108),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_470),
.A2(n_473),
.B1(n_477),
.B2(n_3),
.Y(n_479)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

AOI322xp5_ASAP7_75t_L g473 ( 
.A1(n_457),
.A2(n_148),
.A3(n_96),
.B1(n_132),
.B2(n_130),
.C1(n_192),
.C2(n_98),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_474),
.B(n_464),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_192),
.C(n_2),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_476),
.A2(n_6),
.B(n_7),
.Y(n_482)
);

AOI322xp5_ASAP7_75t_L g477 ( 
.A1(n_463),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_478),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_479),
.B(n_480),
.C(n_482),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_459),
.C(n_6),
.Y(n_483)
);

AOI321xp33_ASAP7_75t_L g486 ( 
.A1(n_483),
.A2(n_469),
.A3(n_474),
.B1(n_475),
.B2(n_476),
.C(n_480),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_486),
.B(n_475),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_487),
.B(n_488),
.C(n_485),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_481),
.Y(n_488)
);


endmodule