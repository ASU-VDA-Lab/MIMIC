module real_aes_7293_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_749;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_1), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_1), .Y(n_460) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_2), .A2(n_151), .B(n_156), .C(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_3), .A2(n_146), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g508 ( .A(n_4), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_5), .B(n_184), .Y(n_250) );
AOI21xp33_ASAP7_75t_L g515 ( .A1(n_6), .A2(n_146), .B(n_516), .Y(n_515) );
AND2x6_ASAP7_75t_L g151 ( .A(n_7), .B(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_8), .A2(n_281), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g163 ( .A(n_9), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_10), .B(n_116), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_10), .B(n_43), .Y(n_127) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_11), .A2(n_33), .B1(n_463), .B2(n_464), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_11), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_12), .B(n_161), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_13), .B(n_208), .Y(n_487) );
INVx1_ASAP7_75t_L g520 ( .A(n_14), .Y(n_520) );
INVx1_ASAP7_75t_L g144 ( .A(n_15), .Y(n_144) );
INVx1_ASAP7_75t_L g499 ( .A(n_16), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g177 ( .A1(n_17), .A2(n_164), .B(n_178), .C(n_182), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_18), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_19), .B(n_478), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_20), .B(n_146), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_21), .B(n_290), .Y(n_289) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_22), .A2(n_208), .B(n_209), .C(n_211), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_23), .B(n_184), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_24), .B(n_161), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_25), .A2(n_180), .B(n_182), .C(n_498), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_26), .B(n_161), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g232 ( .A(n_27), .Y(n_232) );
INVx1_ASAP7_75t_L g220 ( .A(n_28), .Y(n_220) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_29), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_30), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_31), .B(n_161), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_32), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g463 ( .A(n_33), .Y(n_463) );
INVx1_ASAP7_75t_L g286 ( .A(n_34), .Y(n_286) );
INVx1_ASAP7_75t_L g528 ( .A(n_35), .Y(n_528) );
INVx2_ASAP7_75t_L g149 ( .A(n_36), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_37), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_38), .A2(n_208), .B(n_246), .C(n_248), .Y(n_245) );
INVxp67_ASAP7_75t_L g287 ( .A(n_39), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_40), .A2(n_156), .B(n_219), .C(n_225), .Y(n_218) );
CKINVDCx14_ASAP7_75t_R g244 ( .A(n_41), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_42), .A2(n_151), .B(n_156), .C(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g116 ( .A(n_43), .Y(n_116) );
INVx1_ASAP7_75t_L g527 ( .A(n_44), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g159 ( .A1(n_45), .A2(n_160), .B(n_162), .C(n_165), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_46), .B(n_161), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_47), .A2(n_105), .B1(n_117), .B2(n_754), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_48), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g283 ( .A(n_49), .Y(n_283) );
INVx1_ASAP7_75t_L g206 ( .A(n_50), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_51), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_52), .B(n_146), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_53), .A2(n_156), .B1(n_211), .B2(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_54), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_55), .Y(n_505) );
CKINVDCx14_ASAP7_75t_R g154 ( .A(n_56), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_57), .A2(n_160), .B(n_248), .C(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_58), .Y(n_565) );
INVx1_ASAP7_75t_L g517 ( .A(n_59), .Y(n_517) );
INVx1_ASAP7_75t_L g152 ( .A(n_60), .Y(n_152) );
INVx1_ASAP7_75t_L g143 ( .A(n_61), .Y(n_143) );
INVx1_ASAP7_75t_SL g247 ( .A(n_62), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_63), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_64), .B(n_184), .Y(n_213) );
INVx1_ASAP7_75t_L g235 ( .A(n_65), .Y(n_235) );
A2O1A1Ixp33_ASAP7_75t_SL g536 ( .A1(n_66), .A2(n_248), .B(n_478), .C(n_537), .Y(n_536) );
INVxp67_ASAP7_75t_L g538 ( .A(n_67), .Y(n_538) );
INVx1_ASAP7_75t_L g113 ( .A(n_68), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_69), .A2(n_146), .B(n_153), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_70), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_71), .A2(n_146), .B(n_175), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_72), .Y(n_531) );
INVx1_ASAP7_75t_L g559 ( .A(n_73), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_74), .A2(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g176 ( .A(n_75), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g217 ( .A(n_76), .Y(n_217) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_77), .A2(n_78), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_77), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_78), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_79), .A2(n_151), .B(n_156), .C(n_561), .Y(n_560) );
AOI22xp5_ASAP7_75t_SL g454 ( .A1(n_80), .A2(n_125), .B1(n_455), .B2(n_749), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_81), .A2(n_146), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g179 ( .A(n_82), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_83), .B(n_221), .Y(n_476) );
INVx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
INVx1_ASAP7_75t_L g195 ( .A(n_85), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_86), .B(n_478), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_87), .A2(n_151), .B(n_156), .C(n_507), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_88), .B(n_110), .C(n_111), .Y(n_109) );
OR2x2_ASAP7_75t_L g124 ( .A(n_88), .B(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g747 ( .A(n_88), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_89), .A2(n_156), .B(n_234), .C(n_237), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_90), .A2(n_92), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_90), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_91), .B(n_140), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_92), .Y(n_130) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_93), .A2(n_151), .B(n_156), .C(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_94), .Y(n_491) );
INVx1_ASAP7_75t_L g535 ( .A(n_95), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g496 ( .A(n_96), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_97), .B(n_221), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_98), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_99), .B(n_169), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_100), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g210 ( .A(n_101), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_102), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g457 ( .A(n_102), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_103), .A2(n_146), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g754 ( .A(n_107), .Y(n_754) );
AND2x2_ASAP7_75t_SL g107 ( .A(n_108), .B(n_114), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
AND2x2_ASAP7_75t_L g126 ( .A(n_110), .B(n_127), .Y(n_126) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_122), .B(n_453), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g753 ( .A(n_120), .Y(n_753) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_128), .B(n_450), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_124), .Y(n_452) );
NOR2x2_ASAP7_75t_L g751 ( .A(n_125), .B(n_747), .Y(n_751) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B1(n_133), .B2(n_449), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_129), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_130), .B(n_189), .Y(n_511) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
XOR2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_446), .Y(n_133) );
INVx2_ASAP7_75t_L g748 ( .A(n_134), .Y(n_748) );
OR2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_376), .Y(n_134) );
NAND5xp2_ASAP7_75t_L g135 ( .A(n_136), .B(n_291), .C(n_323), .D(n_340), .E(n_363), .Y(n_135) );
AOI221xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_214), .B1(n_251), .B2(n_255), .C(n_259), .Y(n_136) );
INVx1_ASAP7_75t_L g403 ( .A(n_137), .Y(n_403) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_186), .Y(n_137) );
AND3x2_ASAP7_75t_L g378 ( .A(n_138), .B(n_188), .C(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_171), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_139), .B(n_257), .Y(n_256) );
BUFx3_ASAP7_75t_L g266 ( .A(n_139), .Y(n_266) );
AND2x2_ASAP7_75t_L g270 ( .A(n_139), .B(n_202), .Y(n_270) );
INVx2_ASAP7_75t_L g300 ( .A(n_139), .Y(n_300) );
OR2x2_ASAP7_75t_L g311 ( .A(n_139), .B(n_203), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_139), .B(n_187), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_139), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g390 ( .A(n_139), .B(n_203), .Y(n_390) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_145), .B(n_168), .Y(n_139) );
INVx1_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g216 ( .A1(n_140), .A2(n_192), .B(n_217), .C(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g240 ( .A(n_140), .Y(n_240) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_140), .A2(n_494), .B(n_500), .Y(n_493) );
AND2x2_ASAP7_75t_SL g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x2_ASAP7_75t_L g170 ( .A(n_141), .B(n_142), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx2_ASAP7_75t_L g281 ( .A(n_146), .Y(n_281) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_147), .B(n_151), .Y(n_192) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g224 ( .A(n_148), .Y(n_224) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
INVx1_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
INVx1_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
INVx3_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
INVx1_ASAP7_75t_L g478 ( .A(n_150), .Y(n_478) );
INVx4_ASAP7_75t_SL g167 ( .A(n_151), .Y(n_167) );
BUFx3_ASAP7_75t_L g225 ( .A(n_151), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g153 ( .A1(n_154), .A2(n_155), .B(n_159), .C(n_167), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_SL g175 ( .A1(n_155), .A2(n_167), .B(n_176), .C(n_177), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_SL g205 ( .A1(n_155), .A2(n_167), .B(n_206), .C(n_207), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_155), .A2(n_167), .B(n_244), .C(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_SL g282 ( .A1(n_155), .A2(n_167), .B(n_283), .C(n_284), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_155), .A2(n_167), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_155), .A2(n_167), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_155), .A2(n_167), .B(n_535), .C(n_536), .Y(n_534) );
INVx5_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx3_ASAP7_75t_L g166 ( .A(n_157), .Y(n_166) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_157), .Y(n_249) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g208 ( .A(n_161), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
INVx5_ASAP7_75t_L g221 ( .A(n_164), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_164), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_164), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
INVx1_ASAP7_75t_L g237 ( .A(n_167), .Y(n_237) );
OAI22xp33_ASAP7_75t_L g524 ( .A1(n_167), .A2(n_192), .B1(n_525), .B2(n_529), .Y(n_524) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_169), .Y(n_173) );
INVx4_ASAP7_75t_L g185 ( .A(n_169), .Y(n_185) );
OA21x2_ASAP7_75t_L g532 ( .A1(n_169), .A2(n_533), .B(n_539), .Y(n_532) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g278 ( .A(n_170), .Y(n_278) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_171), .Y(n_269) );
AND2x2_ASAP7_75t_L g331 ( .A(n_171), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_171), .B(n_187), .Y(n_350) );
INVx1_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
OR2x2_ASAP7_75t_L g258 ( .A(n_172), .B(n_187), .Y(n_258) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_172), .Y(n_265) );
AND2x2_ASAP7_75t_L g317 ( .A(n_172), .B(n_203), .Y(n_317) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_172), .B(n_186), .C(n_300), .Y(n_342) );
AND2x2_ASAP7_75t_L g407 ( .A(n_172), .B(n_188), .Y(n_407) );
AND2x2_ASAP7_75t_L g441 ( .A(n_172), .B(n_187), .Y(n_441) );
OA21x2_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_183), .Y(n_172) );
OA21x2_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_204), .B(n_213), .Y(n_203) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_173), .A2(n_242), .B(n_250), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_180), .B(n_210), .Y(n_209) );
OAI22xp33_ASAP7_75t_L g285 ( .A1(n_180), .A2(n_221), .B1(n_286), .B2(n_287), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_180), .B(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g197 ( .A(n_181), .Y(n_197) );
OAI22xp5_ASAP7_75t_SL g526 ( .A1(n_181), .A2(n_197), .B1(n_527), .B2(n_528), .Y(n_526) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_184), .A2(n_515), .B(n_521), .Y(n_514) );
INVx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_185), .B(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_185), .B(n_227), .Y(n_226) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_185), .A2(n_231), .B(n_238), .Y(n_230) );
NOR2xp33_ASAP7_75t_SL g479 ( .A(n_185), .B(n_480), .Y(n_479) );
INVxp67_ASAP7_75t_L g267 ( .A(n_186), .Y(n_267) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_202), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_187), .B(n_300), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_187), .B(n_331), .Y(n_339) );
AND2x2_ASAP7_75t_L g389 ( .A(n_187), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g417 ( .A(n_187), .Y(n_417) );
INVx4_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x2_ASAP7_75t_L g324 ( .A(n_188), .B(n_317), .Y(n_324) );
BUFx3_ASAP7_75t_L g356 ( .A(n_188), .Y(n_356) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_200), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_189), .B(n_491), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_189), .B(n_565), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_192), .A2(n_232), .B(n_233), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_192), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_192), .A2(n_559), .B(n_560), .Y(n_558) );
O2A1O1Ixp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_198), .C(n_199), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g234 ( .A1(n_196), .A2(n_199), .B(n_235), .C(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_199), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_199), .A2(n_562), .B(n_563), .Y(n_561) );
INVx2_ASAP7_75t_L g332 ( .A(n_202), .Y(n_332) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_203), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_208), .B(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g510 ( .A(n_211), .Y(n_510) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_214), .A2(n_392), .B1(n_394), .B2(n_395), .Y(n_391) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_228), .Y(n_214) );
AND2x2_ASAP7_75t_L g251 ( .A(n_215), .B(n_252), .Y(n_251) );
INVx3_ASAP7_75t_SL g262 ( .A(n_215), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_215), .B(n_295), .Y(n_327) );
OR2x2_ASAP7_75t_L g346 ( .A(n_215), .B(n_229), .Y(n_346) );
AND2x2_ASAP7_75t_L g351 ( .A(n_215), .B(n_303), .Y(n_351) );
AND2x2_ASAP7_75t_L g354 ( .A(n_215), .B(n_296), .Y(n_354) );
AND2x2_ASAP7_75t_L g366 ( .A(n_215), .B(n_241), .Y(n_366) );
AND2x2_ASAP7_75t_L g382 ( .A(n_215), .B(n_230), .Y(n_382) );
AND2x4_ASAP7_75t_L g385 ( .A(n_215), .B(n_253), .Y(n_385) );
OR2x2_ASAP7_75t_L g402 ( .A(n_215), .B(n_338), .Y(n_402) );
OR2x2_ASAP7_75t_L g433 ( .A(n_215), .B(n_275), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_215), .B(n_361), .Y(n_435) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_226), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_222), .C(n_223), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_221), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_224), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g309 ( .A(n_228), .B(n_273), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_228), .B(n_296), .Y(n_428) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_241), .Y(n_228) );
AND2x2_ASAP7_75t_L g261 ( .A(n_229), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g295 ( .A(n_229), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g303 ( .A(n_229), .B(n_275), .Y(n_303) );
AND2x2_ASAP7_75t_L g321 ( .A(n_229), .B(n_253), .Y(n_321) );
OR2x2_ASAP7_75t_L g338 ( .A(n_229), .B(n_296), .Y(n_338) );
INVx2_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
BUFx2_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
AND2x2_ASAP7_75t_L g361 ( .A(n_230), .B(n_241), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g290 ( .A(n_240), .Y(n_290) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_240), .A2(n_483), .B(n_490), .Y(n_482) );
INVx2_ASAP7_75t_L g253 ( .A(n_241), .Y(n_253) );
INVx1_ASAP7_75t_L g373 ( .A(n_241), .Y(n_373) );
AND2x2_ASAP7_75t_L g423 ( .A(n_241), .B(n_262), .Y(n_423) );
INVx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_249), .Y(n_488) );
AND2x2_ASAP7_75t_L g272 ( .A(n_252), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g307 ( .A(n_252), .B(n_262), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_252), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
AND2x2_ASAP7_75t_L g294 ( .A(n_253), .B(n_262), .Y(n_294) );
OR2x2_ASAP7_75t_L g410 ( .A(n_254), .B(n_384), .Y(n_410) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_257), .B(n_390), .Y(n_396) );
INVx2_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
OAI32xp33_ASAP7_75t_L g352 ( .A1(n_258), .A2(n_353), .A3(n_355), .B1(n_357), .B2(n_358), .Y(n_352) );
OR2x2_ASAP7_75t_L g369 ( .A(n_258), .B(n_311), .Y(n_369) );
OAI21xp33_ASAP7_75t_SL g394 ( .A1(n_258), .A2(n_268), .B(n_299), .Y(n_394) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_263), .B1(n_268), .B2(n_271), .Y(n_259) );
INVxp33_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_261), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_262), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g320 ( .A(n_262), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g420 ( .A(n_262), .B(n_361), .Y(n_420) );
OR2x2_ASAP7_75t_L g444 ( .A(n_262), .B(n_338), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g427 ( .A1(n_263), .A2(n_326), .B(n_428), .Y(n_427) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g304 ( .A(n_265), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_265), .B(n_270), .Y(n_322) );
AND2x2_ASAP7_75t_L g344 ( .A(n_266), .B(n_317), .Y(n_344) );
INVx1_ASAP7_75t_L g357 ( .A(n_266), .Y(n_357) );
OR2x2_ASAP7_75t_L g362 ( .A(n_266), .B(n_296), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_269), .B(n_311), .Y(n_310) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_270), .A2(n_293), .B1(n_298), .B2(n_302), .Y(n_292) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_273), .A2(n_335), .B1(n_342), .B2(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_L g419 ( .A(n_273), .B(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_275), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g438 ( .A(n_275), .B(n_321), .Y(n_438) );
AO21x2_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_279), .B(n_288), .Y(n_275) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_276), .A2(n_558), .B(n_564), .Y(n_557) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI21xp5_ASAP7_75t_SL g472 ( .A1(n_277), .A2(n_473), .B(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_278), .A2(n_504), .B(n_511), .Y(n_503) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_278), .A2(n_524), .B(n_530), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_278), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_280), .A2(n_289), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_304), .B1(n_305), .B2(n_310), .C(n_312), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_294), .B(n_296), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_294), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g313 ( .A(n_295), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_295), .A2(n_401), .B(n_402), .C(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_L g405 ( .A(n_295), .B(n_385), .Y(n_405) );
O2A1O1Ixp33_ASAP7_75t_SL g443 ( .A1(n_295), .A2(n_384), .B(n_444), .C(n_445), .Y(n_443) );
BUFx3_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_299), .B(n_356), .Y(n_399) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_299), .A2(n_419), .B(n_421), .C(n_427), .Y(n_418) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVxp67_ASAP7_75t_L g379 ( .A(n_301), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_303), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g323 ( .A1(n_307), .A2(n_324), .B(n_325), .C(n_333), .Y(n_323) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g408 ( .A(n_311), .Y(n_408) );
OR2x2_ASAP7_75t_L g425 ( .A(n_311), .B(n_355), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_319), .B2(n_322), .Y(n_312) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_314), .A2(n_326), .B1(n_327), .B2(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_318), .Y(n_315) );
OR2x2_ASAP7_75t_L g412 ( .A(n_316), .B(n_356), .Y(n_412) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g367 ( .A(n_317), .B(n_357), .Y(n_367) );
INVx1_ASAP7_75t_L g375 ( .A(n_318), .Y(n_375) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_321), .B(n_335), .Y(n_383) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_331), .B(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g440 ( .A(n_332), .Y(n_440) );
AOI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_336), .B(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_335), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_335), .B(n_366), .Y(n_365) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_335), .B(n_361), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_335), .B(n_382), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g397 ( .A1(n_335), .A2(n_345), .B(n_385), .C(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
AOI221xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_345), .B1(n_347), .B2(n_351), .C(n_352), .Y(n_340) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_349), .B(n_357), .Y(n_431) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_351), .A2(n_366), .B(n_368), .C(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_354), .B(n_361), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_355), .B(n_408), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
INVxp33_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
AOI21xp33_ASAP7_75t_SL g371 ( .A1(n_360), .A2(n_372), .B(n_374), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_360), .B(n_433), .Y(n_432) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_361), .B(n_415), .Y(n_414) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B1(n_368), .B2(n_370), .C(n_371), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_367), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g401 ( .A(n_373), .Y(n_401) );
NAND5xp2_ASAP7_75t_L g376 ( .A(n_377), .B(n_404), .C(n_418), .D(n_429), .E(n_442), .Y(n_376) );
AOI211xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_387), .C(n_400), .Y(n_377) );
INVx2_ASAP7_75t_SL g424 ( .A(n_378), .Y(n_424) );
NAND4xp25_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .C(n_384), .D(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_386), .A2(n_388), .B(n_391), .C(n_397), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_389), .A2(n_430), .B1(n_432), .B2(n_434), .C(n_436), .Y(n_429) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI221xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_406), .B1(n_409), .B2(n_411), .C(n_413), .Y(n_404) );
AND2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_412), .A2(n_435), .B1(n_437), .B2(n_439), .Y(n_436) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g453 ( .A(n_450), .B(n_454), .C(n_752), .Y(n_453) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
XOR2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_465), .Y(n_455) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_745), .B1(n_746), .B2(n_748), .Y(n_465) );
AND2x2_ASAP7_75t_SL g466 ( .A(n_467), .B(n_714), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_607), .C(n_680), .Y(n_467) );
OAI211xp5_ASAP7_75t_SL g468 ( .A1(n_469), .A2(n_501), .B(n_540), .C(n_591), .Y(n_468) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .Y(n_470) );
AND2x2_ASAP7_75t_L g556 ( .A(n_471), .B(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g574 ( .A(n_471), .Y(n_574) );
INVx2_ASAP7_75t_L g589 ( .A(n_471), .Y(n_589) );
INVx1_ASAP7_75t_L g619 ( .A(n_471), .Y(n_619) );
AND2x2_ASAP7_75t_L g669 ( .A(n_471), .B(n_590), .Y(n_669) );
AOI32xp33_ASAP7_75t_L g696 ( .A1(n_471), .A2(n_624), .A3(n_697), .B1(n_699), .B2(n_700), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_471), .B(n_546), .Y(n_702) );
AND2x2_ASAP7_75t_L g729 ( .A(n_471), .B(n_572), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_471), .B(n_738), .Y(n_737) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_479), .Y(n_471) );
AND2x2_ASAP7_75t_L g618 ( .A(n_481), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g640 ( .A(n_481), .Y(n_640) );
AND2x2_ASAP7_75t_L g725 ( .A(n_481), .B(n_556), .Y(n_725) );
AND2x2_ASAP7_75t_L g728 ( .A(n_481), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_492), .Y(n_481) );
INVx2_ASAP7_75t_L g548 ( .A(n_482), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_482), .B(n_572), .Y(n_578) );
AND2x2_ASAP7_75t_L g588 ( .A(n_482), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g624 ( .A(n_482), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_489), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_488), .Y(n_485) );
AND2x2_ASAP7_75t_L g566 ( .A(n_492), .B(n_548), .Y(n_566) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
AND2x2_ASAP7_75t_L g590 ( .A(n_493), .B(n_572), .Y(n_590) );
AND2x2_ASAP7_75t_L g659 ( .A(n_493), .B(n_557), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
OR2x2_ASAP7_75t_L g554 ( .A(n_502), .B(n_523), .Y(n_554) );
INVx1_ASAP7_75t_L g632 ( .A(n_502), .Y(n_632) );
AND2x2_ASAP7_75t_L g646 ( .A(n_502), .B(n_647), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_502), .B(n_522), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_502), .B(n_644), .Y(n_698) );
AND2x2_ASAP7_75t_L g706 ( .A(n_502), .B(n_707), .Y(n_706) );
INVx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx3_ASAP7_75t_L g544 ( .A(n_503), .Y(n_544) );
AND2x2_ASAP7_75t_L g613 ( .A(n_503), .B(n_523), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_512), .B(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g740 ( .A(n_512), .Y(n_740) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_522), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_513), .B(n_584), .Y(n_606) );
OR2x2_ASAP7_75t_L g635 ( .A(n_513), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g667 ( .A(n_513), .B(n_647), .Y(n_667) );
INVx1_ASAP7_75t_SL g687 ( .A(n_513), .Y(n_687) );
AND2x2_ASAP7_75t_L g691 ( .A(n_513), .B(n_553), .Y(n_691) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_SL g545 ( .A(n_514), .B(n_522), .Y(n_545) );
AND2x2_ASAP7_75t_L g552 ( .A(n_514), .B(n_532), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_514), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g594 ( .A(n_514), .B(n_576), .Y(n_594) );
INVx1_ASAP7_75t_SL g601 ( .A(n_514), .Y(n_601) );
BUFx2_ASAP7_75t_L g612 ( .A(n_514), .Y(n_612) );
AND2x2_ASAP7_75t_L g628 ( .A(n_514), .B(n_544), .Y(n_628) );
AND2x2_ASAP7_75t_L g643 ( .A(n_514), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g707 ( .A(n_514), .B(n_523), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_522), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g631 ( .A(n_522), .B(n_632), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_522), .A2(n_649), .B1(n_652), .B2(n_655), .C(n_660), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_522), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_532), .Y(n_522) );
INVx3_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
BUFx2_ASAP7_75t_L g586 ( .A(n_532), .Y(n_586) );
AND2x2_ASAP7_75t_L g600 ( .A(n_532), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g617 ( .A(n_532), .Y(n_617) );
OR2x2_ASAP7_75t_L g636 ( .A(n_532), .B(n_576), .Y(n_636) );
INVx3_ASAP7_75t_L g644 ( .A(n_532), .Y(n_644) );
AND2x2_ASAP7_75t_L g647 ( .A(n_532), .B(n_576), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B1(n_550), .B2(n_555), .C(n_567), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_545), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_543), .B(n_616), .Y(n_741) );
OR2x2_ASAP7_75t_L g744 ( .A(n_543), .B(n_575), .Y(n_744) );
INVx1_ASAP7_75t_SL g543 ( .A(n_544), .Y(n_543) );
OAI221xp5_ASAP7_75t_SL g567 ( .A1(n_544), .A2(n_568), .B1(n_575), .B2(n_577), .C(n_580), .Y(n_567) );
AND2x2_ASAP7_75t_L g584 ( .A(n_544), .B(n_576), .Y(n_584) );
AND2x2_ASAP7_75t_L g592 ( .A(n_544), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_544), .B(n_600), .Y(n_599) );
NAND2x1_ASAP7_75t_L g642 ( .A(n_544), .B(n_643), .Y(n_642) );
OR2x2_ASAP7_75t_L g694 ( .A(n_544), .B(n_636), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_546), .A2(n_654), .B1(n_683), .B2(n_685), .Y(n_682) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI322xp5_ASAP7_75t_L g591 ( .A1(n_547), .A2(n_556), .A3(n_592), .B1(n_595), .B2(n_598), .C1(n_602), .C2(n_605), .Y(n_591) );
OR2x2_ASAP7_75t_L g603 ( .A(n_547), .B(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_548), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g582 ( .A(n_548), .B(n_557), .Y(n_582) );
INVx1_ASAP7_75t_L g597 ( .A(n_548), .Y(n_597) );
AND2x2_ASAP7_75t_L g663 ( .A(n_548), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g573 ( .A(n_549), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g664 ( .A(n_549), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_549), .B(n_572), .Y(n_738) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_553), .B(n_687), .Y(n_686) );
INVx3_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g638 ( .A(n_554), .B(n_585), .Y(n_638) );
OR2x2_ASAP7_75t_L g735 ( .A(n_554), .B(n_586), .Y(n_735) );
INVx1_ASAP7_75t_L g716 ( .A(n_555), .Y(n_716) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_566), .Y(n_555) );
INVx4_ASAP7_75t_L g604 ( .A(n_556), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_556), .B(n_623), .Y(n_629) );
INVx2_ASAP7_75t_L g572 ( .A(n_557), .Y(n_572) );
INVx1_ASAP7_75t_L g654 ( .A(n_566), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_566), .B(n_626), .Y(n_695) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_568), .A2(n_642), .B(n_645), .Y(n_641) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_573), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g626 ( .A(n_572), .Y(n_626) );
INVx1_ASAP7_75t_L g653 ( .A(n_572), .Y(n_653) );
INVx1_ASAP7_75t_L g579 ( .A(n_573), .Y(n_579) );
AND2x2_ASAP7_75t_L g581 ( .A(n_573), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g677 ( .A(n_574), .B(n_663), .Y(n_677) );
AND2x2_ASAP7_75t_L g699 ( .A(n_574), .B(n_659), .Y(n_699) );
BUFx2_ASAP7_75t_L g651 ( .A(n_576), .Y(n_651) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AOI32xp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .A3(n_584), .B1(n_585), .B2(n_587), .Y(n_580) );
INVx1_ASAP7_75t_L g661 ( .A(n_581), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_581), .A2(n_709), .B1(n_710), .B2(n_712), .Y(n_708) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_584), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_584), .B(n_643), .Y(n_684) );
AND2x2_ASAP7_75t_L g731 ( .A(n_584), .B(n_616), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_585), .B(n_632), .Y(n_679) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g732 ( .A(n_587), .Y(n_732) );
AND2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx1_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_590), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g704 ( .A(n_590), .B(n_624), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_590), .B(n_619), .Y(n_711) );
INVx1_ASAP7_75t_SL g693 ( .A(n_592), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_593), .B(n_644), .Y(n_671) );
NOR4xp25_ASAP7_75t_L g717 ( .A(n_593), .B(n_616), .C(n_718), .D(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_594), .B(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVxp67_ASAP7_75t_L g674 ( .A(n_597), .Y(n_674) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g724 ( .A1(n_600), .A2(n_691), .B(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_L g616 ( .A(n_601), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g665 ( .A(n_604), .Y(n_665) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND4xp25_ASAP7_75t_SL g607 ( .A(n_608), .B(n_633), .C(n_648), .D(n_668), .Y(n_607) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_614), .B(n_618), .C(n_620), .Y(n_608) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g700 ( .A(n_613), .B(n_643), .Y(n_700) );
AND2x2_ASAP7_75t_L g709 ( .A(n_613), .B(n_687), .Y(n_709) );
INVx3_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_616), .B(n_651), .Y(n_713) );
AND2x2_ASAP7_75t_L g625 ( .A(n_619), .B(n_626), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_627), .B1(n_629), .B2(n_630), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
AND2x2_ASAP7_75t_L g723 ( .A(n_623), .B(n_669), .Y(n_723) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_625), .B(n_674), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_626), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
O2A1O1Ixp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_637), .B(n_639), .C(n_641), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_634), .A2(n_669), .B1(n_670), .B2(n_672), .C(n_675), .Y(n_668) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g726 ( .A1(n_642), .A2(n_727), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_643), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_651), .B(n_720), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g681 ( .A(n_653), .Y(n_681) );
INVx1_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_656), .A2(n_676), .B1(n_678), .B2(n_679), .Y(n_675) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_666), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_665), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_676), .A2(n_702), .B1(n_740), .B2(n_741), .C(n_742), .Y(n_739) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g721 ( .A(n_678), .Y(n_721) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_688), .C(n_708), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_692), .C(n_701), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B(n_695), .C(n_696), .Y(n_692) );
INVx1_ASAP7_75t_L g720 ( .A(n_698), .Y(n_720) );
OAI21xp5_ASAP7_75t_SL g742 ( .A1(n_699), .A2(n_725), .B(n_743), .Y(n_742) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_703), .B(n_705), .Y(n_701) );
INVx1_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g734 ( .A1(n_711), .A2(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_726), .C(n_739), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_716), .A2(n_717), .B(n_722), .C(n_724), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
CKINVDCx14_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
endmodule