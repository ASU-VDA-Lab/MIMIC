module fake_jpeg_12746_n_85 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx8_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_45),
.Y(n_49)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_0),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_29),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_3),
.B(n_4),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_59),
.B1(n_23),
.B2(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_62),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_63),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_6),
.B(n_7),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_3),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_32),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_5),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_5),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_27),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_32),
.C(n_27),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_68),
.B(n_70),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_6),
.C(n_17),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_72),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_21),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_75),
.B(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_67),
.B(n_66),
.Y(n_79)
);

XNOR2x1_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_79),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_74),
.B1(n_70),
.B2(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_26),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_25),
.Y(n_85)
);


endmodule