module real_jpeg_25591_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_221;
wire n_292;
wire n_215;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_273;
wire n_253;
wire n_89;

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_0),
.B(n_43),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_0),
.B(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_0),
.B(n_31),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_0),
.B(n_17),
.Y(n_231)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_45),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_36),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_2),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_5),
.B(n_43),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_5),
.B(n_25),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_5),
.B(n_36),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_5),
.B(n_31),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_5),
.B(n_62),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_5),
.B(n_45),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_6),
.B(n_51),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_6),
.B(n_25),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_6),
.B(n_31),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_6),
.B(n_62),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_6),
.B(n_36),
.Y(n_233)
);

INVx8_ASAP7_75t_SL g53 ( 
.A(n_7),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_8),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_8),
.B(n_51),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_8),
.B(n_25),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_8),
.B(n_31),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_8),
.B(n_45),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_8),
.B(n_36),
.Y(n_196)
);

NAND2x1_ASAP7_75t_SL g211 ( 
.A(n_8),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_8),
.B(n_43),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_9),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_9),
.B(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_9),
.B(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_9),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_9),
.B(n_31),
.Y(n_239)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_11),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_43),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_11),
.B(n_31),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_11),
.B(n_135),
.Y(n_134)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_12),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_13),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_13),
.B(n_43),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_13),
.B(n_25),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_13),
.B(n_45),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_13),
.B(n_36),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_13),
.B(n_51),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_16),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_16),
.B(n_51),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_16),
.B(n_45),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_16),
.B(n_43),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_16),
.B(n_31),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_16),
.B(n_36),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_16),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_16),
.B(n_25),
.Y(n_246)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_17),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_155),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_33),
.B2(n_38),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_32),
.B(n_147),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_38),
.B1(n_60),
.B2(n_64),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_33),
.B(n_57),
.C(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_34),
.B(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_35),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_47),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_41),
.B(n_42),
.CI(n_44),
.CON(n_71),
.SN(n_71)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx24_ASAP7_75t_SL g304 ( 
.A(n_47),
.Y(n_304)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_49),
.CI(n_50),
.CON(n_47),
.SN(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_52),
.B(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_65),
.C(n_71),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_56),
.B(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_64),
.B1(n_66),
.B2(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g212 ( 
.A(n_63),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_66),
.C(n_67),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_65),
.B(n_71),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_66),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_67),
.A2(n_68),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g301 ( 
.A(n_71),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_86),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_84),
.C(n_85),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_75),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.C(n_81),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_78),
.CI(n_81),
.CON(n_95),
.SN(n_95)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_85),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_88),
.Y(n_90)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_106),
.C(n_110),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_106),
.CI(n_110),
.CON(n_125),
.SN(n_125)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.C(n_102),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_95),
.B(n_292),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_95),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_96),
.B(n_102),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.C(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_97),
.A2(n_98),
.B1(n_100),
.B2(n_101),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_99),
.B(n_279),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_107),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_122),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_119),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_119),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_114),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_122),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_129),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_124),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_299)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_125),
.Y(n_300)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_129),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_142),
.C(n_144),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_130),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.C(n_138),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_131),
.B(n_285),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_133),
.A2(n_134),
.B(n_137),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_133),
.B(n_138),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.C(n_141),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_139),
.B(n_140),
.CI(n_141),
.CON(n_258),
.SN(n_258)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_142),
.B(n_144),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_151),
.C(n_153),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_145),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_150),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_146),
.B(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_149),
.B(n_150),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_297),
.C(n_298),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_287),
.C(n_288),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_272),
.C(n_273),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_251),
.C(n_252),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_226),
.C(n_227),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_189),
.C(n_200),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_175),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_170),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_170),
.C(n_175),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_165),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_171),
.B(n_173),
.C(n_174),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_183),
.C(n_184),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_177),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_188),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_199),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_193),
.A2(n_194),
.B1(n_199),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_222),
.C(n_223),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.C(n_215),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_222)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_240),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_241),
.C(n_250),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_236),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_235),
.C(n_236),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_234),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_231),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_234),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g306 ( 
.A(n_236),
.Y(n_306)
);

FAx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.CI(n_239),
.CON(n_236),
.SN(n_236)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_238),
.C(n_239),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_250),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_248),
.B2(n_249),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_244),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_247),
.C(n_249),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_248),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_264),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_256),
.C(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_260),
.C(n_263),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g302 ( 
.A(n_258),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_267),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_268),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_282),
.B2(n_286),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_283),
.C(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_278),
.C(n_280),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_295),
.B2(n_296),
.Y(n_288)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_293),
.C(n_295),
.Y(n_297)
);


endmodule