module fake_jpeg_28107_n_285 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_285);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_49),
.Y(n_66)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

AOI32xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_31),
.A3(n_33),
.B1(n_27),
.B2(n_28),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_62),
.Y(n_86)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_24),
.B1(n_25),
.B2(n_20),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_27),
.B1(n_31),
.B2(n_33),
.Y(n_76)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_60),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_27),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_29),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_33),
.B1(n_31),
.B2(n_35),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_46),
.B1(n_38),
.B2(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_80),
.B1(n_46),
.B2(n_37),
.Y(n_92)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_79),
.B1(n_66),
.B2(n_24),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_64),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_66),
.A2(n_24),
.B1(n_35),
.B2(n_25),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_31),
.B1(n_33),
.B2(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_50),
.Y(n_98)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_87),
.A2(n_88),
.B1(n_37),
.B2(n_47),
.Y(n_94)
);

OAI22x1_ASAP7_75t_L g88 ( 
.A1(n_52),
.A2(n_30),
.B1(n_46),
.B2(n_37),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_75),
.A2(n_65),
.B1(n_54),
.B2(n_52),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_97),
.B1(n_105),
.B2(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_65),
.B1(n_59),
.B2(n_63),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_62),
.B(n_68),
.C(n_34),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_87),
.B(n_18),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_78),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_34),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_91),
.Y(n_123)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_75),
.A2(n_51),
.B1(n_35),
.B2(n_34),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_41),
.B1(n_53),
.B2(n_67),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_98),
.B(n_84),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_17),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_17),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_50),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_103),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_20),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_73),
.A2(n_35),
.B1(n_66),
.B2(n_55),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_20),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_107),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_21),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_77),
.B1(n_83),
.B2(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_129),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_88),
.C(n_80),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_70),
.C(n_36),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_112),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_88),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_93),
.B1(n_82),
.B2(n_15),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_87),
.B1(n_84),
.B2(n_72),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_118),
.A2(n_121),
.B1(n_15),
.B2(n_24),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_97),
.B1(n_90),
.B2(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_123),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_87),
.B1(n_72),
.B2(n_77),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_18),
.B(n_14),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_92),
.B1(n_107),
.B2(n_96),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_110),
.B1(n_127),
.B2(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_127),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_128),
.A2(n_105),
.B(n_90),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_106),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g130 ( 
.A(n_104),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_130),
.A2(n_64),
.B1(n_57),
.B2(n_70),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_135),
.B1(n_139),
.B2(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_133),
.A2(n_137),
.B1(n_153),
.B2(n_154),
.Y(n_158)
);

AO21x2_ASAP7_75t_SL g134 ( 
.A1(n_118),
.A2(n_91),
.B(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_100),
.B1(n_15),
.B2(n_25),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_143),
.B1(n_146),
.B2(n_147),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_141),
.B(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_70),
.B1(n_22),
.B2(n_39),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_110),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_112),
.A2(n_70),
.B(n_11),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_149),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_22),
.B1(n_39),
.B2(n_64),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_22),
.B1(n_14),
.B2(n_18),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_19),
.B(n_14),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_128),
.A2(n_21),
.B1(n_16),
.B2(n_19),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_150),
.A2(n_116),
.B1(n_129),
.B2(n_111),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_16),
.B1(n_30),
.B2(n_23),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_12),
.B1(n_32),
.B2(n_36),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_123),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_171),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_160),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_114),
.C(n_120),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_174),
.C(n_175),
.Y(n_182)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_165),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_163),
.A2(n_133),
.B1(n_154),
.B2(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_113),
.Y(n_164)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_166),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_178),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_153),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_172),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_109),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_173),
.B(n_137),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_116),
.C(n_117),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_130),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_152),
.B(n_130),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_145),
.C(n_141),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_146),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_177),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_130),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_134),
.B1(n_140),
.B2(n_138),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_186),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_157),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_135),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_171),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_134),
.C(n_149),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_163),
.B(n_147),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_197),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_143),
.B1(n_150),
.B2(n_12),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_157),
.B1(n_170),
.B2(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_160),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_202),
.A2(n_217),
.B1(n_188),
.B2(n_199),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_204),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_182),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_212),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_161),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_219),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_174),
.C(n_159),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_198),
.C(n_200),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_156),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_197),
.B(n_193),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_158),
.B1(n_167),
.B2(n_36),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_227),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_230),
.C(n_214),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_229),
.B1(n_209),
.B2(n_207),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_203),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_210),
.A2(n_188),
.B1(n_196),
.B2(n_198),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_190),
.C(n_196),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_181),
.B(n_8),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_231),
.A2(n_7),
.B(n_11),
.Y(n_242)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_235),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_211),
.A2(n_181),
.B1(n_36),
.B2(n_32),
.Y(n_233)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_233),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_201),
.B(n_26),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_205),
.C(n_219),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_246),
.C(n_235),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_1),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_215),
.B1(n_1),
.B2(n_2),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_6),
.B1(n_10),
.B2(n_9),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_26),
.C(n_2),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_228),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_250),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_220),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_224),
.B(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_251),
.B(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_257),
.C(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_225),
.C(n_2),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_247),
.B(n_243),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_266),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_246),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_268),
.Y(n_272)
);

NOR2xp67_ASAP7_75t_SL g264 ( 
.A(n_255),
.B(n_242),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_5),
.B(n_7),
.Y(n_274)
);

INVxp33_ASAP7_75t_L g265 ( 
.A(n_257),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_258),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_274),
.C(n_261),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_3),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_272),
.B(n_273),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_5),
.B(n_6),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_269),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_276),
.A2(n_275),
.B(n_5),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_261),
.B(n_270),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_278),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_280),
.A2(n_279),
.B(n_5),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_10),
.C(n_9),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_2),
.C(n_9),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_9),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_10),
.Y(n_285)
);


endmodule