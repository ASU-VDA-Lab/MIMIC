module fake_aes_7897_n_715 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_715);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_715;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_42), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_38), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_54), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_58), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_17), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_52), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_69), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_35), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_20), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_28), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_43), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_22), .Y(n_92) );
HB1xp67_ASAP7_75t_L g93 ( .A(n_11), .Y(n_93) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_75), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_21), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_15), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_53), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_60), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_31), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_55), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_29), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_41), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_62), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_34), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_76), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_49), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_1), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_45), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_44), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_6), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_72), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_56), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_67), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_57), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_39), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_8), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_1), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_3), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_51), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_30), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_40), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_9), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_2), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_59), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_93), .B(n_0), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_104), .B(n_0), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_111), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_104), .B(n_2), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_104), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_84), .B(n_3), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_111), .B(n_4), .Y(n_135) );
CKINVDCx11_ASAP7_75t_R g136 ( .A(n_79), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_119), .B(n_4), .Y(n_137) );
BUFx2_ASAP7_75t_L g138 ( .A(n_118), .Y(n_138) );
OA21x2_ASAP7_75t_L g139 ( .A1(n_81), .A2(n_32), .B(n_73), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_120), .B(n_5), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_80), .B(n_5), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_82), .Y(n_142) );
CKINVDCx11_ASAP7_75t_R g143 ( .A(n_79), .Y(n_143) );
NOR2xp33_ASAP7_75t_SL g144 ( .A(n_127), .B(n_33), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_118), .B(n_7), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_92), .B(n_7), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_85), .B(n_8), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_92), .B(n_10), .Y(n_152) );
INVxp67_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_94), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_88), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_117), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_97), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_117), .Y(n_160) );
INVx3_ASAP7_75t_L g161 ( .A(n_123), .Y(n_161) );
AND2x2_ASAP7_75t_L g162 ( .A(n_83), .B(n_10), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_100), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_102), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_103), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_83), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_94), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_90), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_114), .B(n_12), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_153), .B(n_126), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_142), .B(n_126), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_138), .B(n_113), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_142), .B(n_122), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
OAI22xp33_ASAP7_75t_L g180 ( .A1(n_138), .A2(n_90), .B1(n_107), .B2(n_113), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_151), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
OR2x2_ASAP7_75t_L g184 ( .A(n_133), .B(n_115), .Y(n_184) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_162), .B(n_94), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_135), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_134), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_154), .B(n_115), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_171), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_171), .B(n_110), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_154), .B(n_121), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_128), .B(n_114), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_171), .B(n_95), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_156), .B(n_112), .Y(n_196) );
OA22x2_ASAP7_75t_L g197 ( .A1(n_135), .A2(n_96), .B1(n_89), .B2(n_106), .Y(n_197) );
AND2x6_ASAP7_75t_L g198 ( .A(n_171), .B(n_95), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_135), .Y(n_199) );
INVxp33_ASAP7_75t_SL g200 ( .A(n_134), .Y(n_200) );
BUFx10_ASAP7_75t_L g201 ( .A(n_135), .Y(n_201) );
OA22x2_ASAP7_75t_L g202 ( .A1(n_156), .A2(n_109), .B1(n_105), .B2(n_101), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_159), .Y(n_203) );
INVx2_ASAP7_75t_SL g204 ( .A(n_167), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_159), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
INVx3_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_158), .B(n_95), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_158), .B(n_98), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_162), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_163), .B(n_95), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_159), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_146), .B(n_107), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_163), .B(n_91), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_164), .B(n_166), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_159), .Y(n_219) );
AND2x2_ASAP7_75t_L g220 ( .A(n_128), .B(n_77), .Y(n_220) );
INVx3_ASAP7_75t_L g221 ( .A(n_146), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_139), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
AND2x2_ASAP7_75t_SL g224 ( .A(n_144), .B(n_14), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_164), .B(n_16), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_147), .Y(n_226) );
INVx6_ASAP7_75t_L g227 ( .A(n_168), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_136), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_165), .B(n_18), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g231 ( .A1(n_165), .A2(n_19), .B1(n_23), .B2(n_24), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_168), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_168), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_168), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_148), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_166), .B(n_25), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_139), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_188), .A2(n_147), .B1(n_170), .B2(n_149), .C(n_152), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_175), .Y(n_239) );
OR2x6_ASAP7_75t_L g240 ( .A(n_215), .B(n_145), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_184), .B(n_137), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_189), .B(n_143), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_200), .A2(n_140), .B1(n_148), .B2(n_160), .Y(n_243) );
NAND2x1_ASAP7_75t_L g244 ( .A(n_191), .B(n_139), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_208), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_195), .A2(n_129), .B(n_139), .Y(n_246) );
INVx2_ASAP7_75t_SL g247 ( .A(n_194), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_215), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_211), .B(n_130), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_191), .B(n_150), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
INVxp67_ASAP7_75t_SL g252 ( .A(n_191), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_198), .B(n_169), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_221), .Y(n_254) );
INVxp67_ASAP7_75t_L g255 ( .A(n_215), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_237), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_200), .A2(n_141), .B1(n_160), .B2(n_157), .Y(n_257) );
CKINVDCx16_ASAP7_75t_R g258 ( .A(n_182), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_218), .B(n_161), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g260 ( .A1(n_199), .A2(n_130), .B1(n_157), .B2(n_169), .C(n_161), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_221), .Y(n_261) );
AOI21x1_ASAP7_75t_L g262 ( .A1(n_195), .A2(n_192), .B(n_236), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_223), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_197), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_218), .B(n_161), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_235), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_235), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_206), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_207), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_201), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_174), .B(n_26), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_178), .B(n_27), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_201), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_197), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_187), .B(n_36), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_201), .B(n_37), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_226), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_190), .B(n_47), .Y(n_278) );
CKINVDCx6p67_ASAP7_75t_R g279 ( .A(n_224), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_220), .B(n_48), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_204), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_172), .B(n_50), .Y(n_282) );
NAND3xp33_ASAP7_75t_L g283 ( .A(n_185), .B(n_61), .C(n_63), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_216), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_172), .B(n_64), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_216), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_224), .A2(n_65), .B1(n_66), .B2(n_68), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_192), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_198), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_217), .B(n_70), .Y(n_290) );
INVxp67_ASAP7_75t_L g291 ( .A(n_193), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_196), .B(n_71), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_217), .B(n_210), .Y(n_293) );
NOR3x1_ASAP7_75t_L g294 ( .A(n_180), .B(n_228), .C(n_202), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_202), .B(n_177), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_177), .B(n_185), .Y(n_296) );
A2O1A1Ixp33_ASAP7_75t_L g297 ( .A1(n_173), .A2(n_230), .B(n_225), .C(n_237), .Y(n_297) );
INVx2_ASAP7_75t_SL g298 ( .A(n_198), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_198), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_173), .B(n_198), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_222), .B(n_237), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_209), .Y(n_302) );
AOI22x1_ASAP7_75t_L g303 ( .A1(n_222), .A2(n_237), .B1(n_179), .B2(n_181), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_222), .A2(n_213), .B1(n_209), .B2(n_227), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_213), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_231), .B(n_176), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_227), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_176), .B(n_179), .Y(n_308) );
OAI21xp5_ASAP7_75t_SL g309 ( .A1(n_243), .A2(n_181), .B(n_183), .Y(n_309) );
AOI21x1_ASAP7_75t_L g310 ( .A1(n_244), .A2(n_183), .B(n_186), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_291), .B(n_227), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_246), .A2(n_186), .B(n_203), .Y(n_312) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_243), .A2(n_203), .B(n_205), .C(n_212), .Y(n_313) );
AO21x1_ASAP7_75t_L g314 ( .A1(n_246), .A2(n_205), .B(n_212), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_270), .B(n_214), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_270), .B(n_214), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_301), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_249), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_291), .B(n_219), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_266), .Y(n_323) );
OAI22x1_ASAP7_75t_L g324 ( .A1(n_242), .A2(n_219), .B1(n_229), .B2(n_232), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_297), .A2(n_229), .B(n_232), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_306), .A2(n_233), .B(n_234), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_267), .Y(n_328) );
INVxp33_ASAP7_75t_SL g329 ( .A(n_294), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_279), .A2(n_233), .B1(n_234), .B2(n_238), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_263), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_293), .B(n_288), .Y(n_332) );
OAI21xp5_ASAP7_75t_L g333 ( .A1(n_306), .A2(n_296), .B(n_295), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_240), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_264), .B(n_274), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_251), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_273), .B(n_290), .Y(n_337) );
NAND2xp5_ASAP7_75t_SL g338 ( .A(n_273), .B(n_290), .Y(n_338) );
INVx6_ASAP7_75t_L g339 ( .A(n_240), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_275), .A2(n_250), .B(n_241), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_248), .A2(n_255), .B1(n_238), .B2(n_239), .C(n_265), .Y(n_341) );
O2A1O1Ixp33_ASAP7_75t_SL g342 ( .A1(n_292), .A2(n_278), .B(n_280), .C(n_271), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_275), .A2(n_252), .B(n_278), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_248), .A2(n_255), .B1(n_260), .B2(n_277), .Y(n_344) );
O2A1O1Ixp5_ASAP7_75t_SL g345 ( .A1(n_272), .A2(n_276), .B(n_307), .C(n_281), .Y(n_345) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_256), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_259), .B(n_265), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_257), .B(n_259), .Y(n_348) );
AOI21x1_ASAP7_75t_L g349 ( .A1(n_262), .A2(n_292), .B(n_308), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_300), .A2(n_304), .B(n_245), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_300), .A2(n_284), .B(n_254), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_286), .B(n_282), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_268), .B(n_269), .Y(n_353) );
NAND3xp33_ASAP7_75t_SL g354 ( .A(n_287), .B(n_260), .C(n_285), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_261), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_253), .A2(n_298), .B1(n_289), .B2(n_299), .Y(n_356) );
BUFx3_ASAP7_75t_L g357 ( .A(n_302), .Y(n_357) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_256), .A2(n_303), .B(n_305), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_308), .A2(n_283), .B(n_256), .Y(n_359) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_256), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_247), .Y(n_361) );
O2A1O1Ixp5_ASAP7_75t_L g362 ( .A1(n_295), .A2(n_244), .B(n_280), .C(n_276), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g363 ( .A1(n_343), .A2(n_342), .B(n_332), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_341), .A2(n_348), .B1(n_329), .B2(n_330), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
AOI21x1_ASAP7_75t_L g366 ( .A1(n_349), .A2(n_314), .B(n_310), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_347), .B(n_321), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_347), .B(n_319), .Y(n_368) );
AND2x6_ASAP7_75t_L g369 ( .A(n_320), .B(n_346), .Y(n_369) );
INVxp67_ASAP7_75t_SL g370 ( .A(n_317), .Y(n_370) );
NAND3x1_ASAP7_75t_L g371 ( .A(n_318), .B(n_361), .C(n_333), .Y(n_371) );
AOI21x1_ASAP7_75t_L g372 ( .A1(n_312), .A2(n_359), .B(n_358), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_327), .B(n_339), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_334), .B(n_337), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_332), .A2(n_360), .B(n_346), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_346), .A2(n_360), .B(n_340), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_322), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_333), .B(n_344), .Y(n_380) );
OAI22x1_ASAP7_75t_L g381 ( .A1(n_338), .A2(n_335), .B1(n_352), .B2(n_355), .Y(n_381) );
BUFx8_ASAP7_75t_L g382 ( .A(n_335), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_311), .Y(n_383) );
INVx8_ASAP7_75t_L g384 ( .A(n_360), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_322), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_353), .B(n_336), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_309), .A2(n_350), .B(n_313), .C(n_362), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_330), .B(n_351), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_357), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_328), .B(n_324), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_356), .B(n_315), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_354), .B(n_309), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_326), .A2(n_325), .B(n_316), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_345), .Y(n_394) );
AOI21x1_ASAP7_75t_L g395 ( .A1(n_349), .A2(n_314), .B(n_244), .Y(n_395) );
OAI21x1_ASAP7_75t_L g396 ( .A1(n_359), .A2(n_310), .B(n_358), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_379), .B(n_385), .Y(n_397) );
AND2x4_ASAP7_75t_L g398 ( .A(n_365), .B(n_368), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_369), .Y(n_399) );
OAI21x1_ASAP7_75t_L g400 ( .A1(n_366), .A2(n_395), .B(n_396), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_367), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_364), .B(n_386), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
AO31x2_ASAP7_75t_L g404 ( .A1(n_392), .A2(n_387), .A3(n_388), .B(n_394), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_364), .B(n_380), .Y(n_405) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_388), .B(n_372), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_391), .B(n_373), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_391), .B(n_389), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_380), .B(n_383), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_374), .B(n_376), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
OAI21x1_ASAP7_75t_L g412 ( .A1(n_393), .A2(n_378), .B(n_371), .Y(n_412) );
AO21x2_ASAP7_75t_L g413 ( .A1(n_377), .A2(n_390), .B(n_381), .Y(n_413) );
CKINVDCx8_ASAP7_75t_R g414 ( .A(n_384), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_382), .B(n_370), .Y(n_415) );
OAI21x1_ASAP7_75t_L g416 ( .A1(n_369), .A2(n_384), .B(n_382), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
AOI21x1_ASAP7_75t_L g418 ( .A1(n_369), .A2(n_366), .B(n_394), .Y(n_418) );
INVx4_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_387), .A2(n_341), .B(n_255), .Y(n_420) );
BUFx8_ASAP7_75t_L g421 ( .A(n_374), .Y(n_421) );
AO21x1_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_388), .B(n_394), .Y(n_422) );
OAI21x1_ASAP7_75t_L g423 ( .A1(n_366), .A2(n_395), .B(n_396), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_364), .B(n_200), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_379), .B(n_385), .Y(n_425) );
OAI21x1_ASAP7_75t_L g426 ( .A1(n_400), .A2(n_423), .B(n_412), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_397), .B(n_425), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_406), .Y(n_428) );
BUFx4f_ASAP7_75t_SL g429 ( .A(n_421), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_403), .Y(n_430) );
BUFx3_ASAP7_75t_L g431 ( .A(n_414), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_397), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_406), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_399), .Y(n_434) );
AO21x2_ASAP7_75t_L g435 ( .A1(n_422), .A2(n_423), .B(n_400), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_404), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_404), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_404), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_425), .B(n_398), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_398), .B(n_401), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_404), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_412), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_401), .B(n_398), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_422), .A2(n_418), .B(n_420), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_418), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_402), .B(n_407), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_405), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_413), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_402), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_402), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
AOI21x1_ASAP7_75t_L g457 ( .A1(n_399), .A2(n_417), .B(n_408), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_407), .B(n_408), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_408), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_407), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_436), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_427), .B(n_410), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_427), .B(n_410), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_429), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_441), .B(n_410), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_437), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_437), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_453), .B(n_416), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_434), .Y(n_471) );
AO21x1_ASAP7_75t_L g472 ( .A1(n_452), .A2(n_424), .B(n_415), .Y(n_472) );
NOR2x1_ASAP7_75t_L g473 ( .A(n_431), .B(n_419), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_438), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_426), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_441), .B(n_411), .Y(n_476) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_447), .A2(n_426), .B(n_433), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_433), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_438), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_439), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_453), .B(n_411), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_455), .B(n_416), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_440), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_455), .B(n_419), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_443), .B(n_419), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_443), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_451), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_447), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_434), .Y(n_491) );
AO21x2_ASAP7_75t_L g492 ( .A1(n_435), .A2(n_414), .B(n_421), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_442), .B(n_421), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_451), .B(n_450), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_442), .B(n_432), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_450), .B(n_432), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_430), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_448), .B(n_449), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_444), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_452), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_434), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_444), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_448), .B(n_460), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_460), .B(n_458), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_458), .B(n_459), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_459), .B(n_446), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_445), .B(n_431), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_454), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_490), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_490), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_495), .B(n_446), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_495), .B(n_446), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_506), .B(n_456), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_500), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_500), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_473), .B(n_434), .Y(n_518) );
INVx3_ASAP7_75t_R g519 ( .A(n_487), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_508), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_506), .B(n_470), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_503), .B(n_456), .Y(n_522) );
INVx4_ASAP7_75t_L g523 ( .A(n_492), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_503), .B(n_435), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_490), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_505), .B(n_435), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_505), .B(n_457), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_504), .B(n_457), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_504), .B(n_434), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_461), .B(n_494), .Y(n_530) );
OR2x2_ASAP7_75t_L g531 ( .A(n_461), .B(n_494), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_470), .B(n_482), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_489), .B(n_509), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_470), .B(n_482), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_498), .B(n_489), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_498), .B(n_509), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_507), .A2(n_472), .B1(n_493), .B2(n_476), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_508), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_475), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_468), .B(n_480), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_464), .B(n_496), .Y(n_541) );
AND2x4_ASAP7_75t_L g542 ( .A(n_470), .B(n_480), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_472), .A2(n_462), .B1(n_465), .B2(n_467), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_468), .B(n_479), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_464), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_469), .B(n_484), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_469), .B(n_484), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_497), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_497), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_462), .B(n_465), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_474), .B(n_479), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_474), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_478), .B(n_483), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_478), .B(n_483), .Y(n_554) );
AND3x1_ASAP7_75t_L g555 ( .A(n_493), .B(n_473), .C(n_467), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_478), .B(n_485), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_476), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_483), .B(n_485), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_485), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_557), .B(n_487), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_550), .B(n_466), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_536), .B(n_487), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_537), .B(n_496), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_548), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_553), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_536), .B(n_487), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_512), .B(n_488), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_512), .B(n_488), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_548), .Y(n_569) );
NAND4xp25_ASAP7_75t_L g570 ( .A(n_537), .B(n_486), .C(n_481), .D(n_475), .Y(n_570) );
AND3x2_ASAP7_75t_L g571 ( .A(n_555), .B(n_486), .C(n_481), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_549), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_530), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_513), .B(n_488), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_530), .B(n_501), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_531), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_513), .B(n_492), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_535), .B(n_492), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_555), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_529), .B(n_492), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_549), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_529), .B(n_471), .Y(n_583) );
INVx2_ASAP7_75t_SL g584 ( .A(n_531), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_535), .B(n_471), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_541), .B(n_501), .Y(n_586) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_553), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_541), .B(n_501), .Y(n_588) );
INVx2_ASAP7_75t_SL g589 ( .A(n_532), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_533), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_532), .B(n_471), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_533), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_516), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_532), .B(n_501), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_516), .Y(n_595) );
INVxp67_ASAP7_75t_SL g596 ( .A(n_515), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_532), .B(n_534), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_517), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_517), .B(n_499), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_534), .B(n_491), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_534), .B(n_491), .Y(n_601) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_534), .B(n_491), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_520), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_521), .B(n_499), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_520), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_475), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_543), .B(n_475), .C(n_477), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_521), .B(n_522), .Y(n_609) );
NOR2xp67_ASAP7_75t_R g610 ( .A(n_519), .B(n_499), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_521), .B(n_502), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_538), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_554), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_594), .Y(n_614) );
INVxp67_ASAP7_75t_L g615 ( .A(n_573), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_578), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_565), .B(n_526), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_565), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_609), .B(n_526), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_590), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_563), .B(n_524), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_592), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_587), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_576), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_587), .B(n_524), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g626 ( .A(n_579), .B(n_523), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_584), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_597), .B(n_528), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_602), .B(n_522), .Y(n_629) );
AOI322xp5_ASAP7_75t_L g630 ( .A1(n_563), .A2(n_528), .A3(n_527), .B1(n_538), .B2(n_542), .C1(n_545), .C2(n_514), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_602), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_578), .B(n_547), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_579), .A2(n_542), .B1(n_527), .B2(n_518), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_564), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_569), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_572), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_589), .B(n_542), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_561), .B(n_519), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_582), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_593), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_570), .A2(n_514), .B1(n_523), .B2(n_545), .Y(n_641) );
NAND4xp25_ASAP7_75t_L g642 ( .A(n_608), .B(n_523), .C(n_539), .D(n_552), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_595), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_598), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_591), .B(n_566), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_575), .Y(n_646) );
A2O1A1Ixp33_ASAP7_75t_L g647 ( .A1(n_571), .A2(n_547), .B(n_540), .C(n_544), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_562), .B(n_546), .Y(n_648) );
OAI21xp5_ASAP7_75t_L g649 ( .A1(n_577), .A2(n_518), .B(n_523), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_567), .B(n_551), .Y(n_650) );
INVx2_ASAP7_75t_SL g651 ( .A(n_585), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_618), .Y(n_652) );
OAI32xp33_ASAP7_75t_L g653 ( .A1(n_616), .A2(n_577), .A3(n_588), .B1(n_586), .B2(n_581), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_621), .B(n_567), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_635), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_625), .B(n_574), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_636), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_621), .B(n_574), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_616), .B(n_568), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_639), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_640), .Y(n_662) );
AOI22x1_ASAP7_75t_L g663 ( .A1(n_649), .A2(n_571), .B1(n_518), .B2(n_610), .Y(n_663) );
OAI322xp33_ASAP7_75t_L g664 ( .A1(n_632), .A2(n_568), .A3(n_605), .B1(n_613), .B2(n_606), .C1(n_612), .C2(n_604), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_647), .A2(n_596), .B(n_601), .Y(n_665) );
INVxp67_ASAP7_75t_SL g666 ( .A(n_623), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g667 ( .A1(n_641), .A2(n_581), .B1(n_603), .B2(n_580), .C(n_607), .Y(n_667) );
NAND2x1_ASAP7_75t_L g668 ( .A(n_633), .B(n_601), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g669 ( .A1(n_630), .A2(n_560), .B(n_596), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_631), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_629), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_643), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_644), .Y(n_673) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_633), .A2(n_539), .B(n_600), .Y(n_674) );
INVx1_ASAP7_75t_SL g675 ( .A(n_614), .Y(n_675) );
OAI321xp33_ASAP7_75t_L g676 ( .A1(n_669), .A2(n_642), .A3(n_649), .B1(n_615), .B2(n_632), .C(n_638), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_668), .A2(n_626), .B(n_614), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g678 ( .A1(n_653), .A2(n_627), .B(n_646), .C(n_620), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_655), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_675), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g681 ( .A1(n_665), .A2(n_650), .B(n_651), .Y(n_681) );
INVxp67_ASAP7_75t_L g682 ( .A(n_656), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_664), .A2(n_650), .B(n_624), .Y(n_683) );
OAI32xp33_ASAP7_75t_L g684 ( .A1(n_667), .A2(n_617), .A3(n_622), .B1(n_628), .B2(n_645), .Y(n_684) );
AOI322xp5_ASAP7_75t_L g685 ( .A1(n_654), .A2(n_619), .A3(n_648), .B1(n_637), .B2(n_611), .C1(n_583), .C2(n_600), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_652), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_659), .B(n_599), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_660), .B(n_661), .Y(n_688) );
OAI21xp33_ASAP7_75t_L g689 ( .A1(n_674), .A2(n_599), .B(n_539), .Y(n_689) );
OAI321xp33_ASAP7_75t_L g690 ( .A1(n_678), .A2(n_673), .A3(n_672), .B1(n_658), .B2(n_662), .C(n_671), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_677), .A2(n_663), .B(n_666), .Y(n_691) );
OAI21xp5_ASAP7_75t_L g692 ( .A1(n_681), .A2(n_666), .B(n_671), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_684), .A2(n_670), .B1(n_652), .B2(n_657), .C(n_552), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_679), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_682), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_686), .Y(n_696) );
AOI21x1_ASAP7_75t_L g697 ( .A1(n_683), .A2(n_670), .B(n_657), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_693), .B(n_685), .C(n_689), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_690), .B(n_676), .C(n_688), .Y(n_699) );
NOR2x1_ASAP7_75t_L g700 ( .A(n_691), .B(n_680), .Y(n_700) );
AOI211xp5_ASAP7_75t_L g701 ( .A1(n_690), .A2(n_687), .B(n_539), .C(n_546), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_697), .A2(n_559), .B(n_551), .C(n_544), .Y(n_702) );
INVxp67_ASAP7_75t_L g703 ( .A(n_700), .Y(n_703) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_698), .Y(n_704) );
NOR3xp33_ASAP7_75t_L g705 ( .A(n_699), .B(n_695), .C(n_692), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_703), .B(n_694), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_705), .A2(n_701), .B1(n_702), .B2(n_696), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_706), .B(n_704), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_707), .B1(n_559), .B2(n_510), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_709), .Y(n_710) );
AOI211xp5_ASAP7_75t_L g711 ( .A1(n_710), .A2(n_540), .B(n_556), .C(n_558), .Y(n_711) );
OAI21xp5_ASAP7_75t_SL g712 ( .A1(n_711), .A2(n_556), .B(n_558), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_712), .A2(n_525), .B(n_510), .Y(n_713) );
AO21x2_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_525), .B(n_511), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_525), .B1(n_511), .B2(n_510), .Y(n_715) );
endmodule