module real_aes_17124_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_889;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_880;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_0), .Y(n_201) );
AND2x4_ASAP7_75t_L g116 ( .A(n_1), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_2), .B(n_496), .Y(n_495) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_2), .B(n_497), .C(n_505), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_2), .B(n_505), .C(n_510), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g882 ( .A(n_3), .Y(n_882) );
BUFx3_ASAP7_75t_L g267 ( .A(n_4), .Y(n_267) );
INVx1_ASAP7_75t_L g117 ( .A(n_5), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_6), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g109 ( .A(n_7), .B(n_22), .Y(n_109) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_8), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_9), .B(n_156), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g539 ( .A(n_10), .B(n_156), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_11), .B(n_182), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_12), .A2(n_84), .B1(n_152), .B2(n_156), .Y(n_155) );
OAI22x1_ASAP7_75t_L g497 ( .A1(n_13), .A2(n_27), .B1(n_498), .B2(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g499 ( .A(n_13), .Y(n_499) );
OAI21x1_ASAP7_75t_L g145 ( .A1(n_14), .A2(n_38), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_15), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_16), .B(n_193), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_17), .Y(n_551) );
AO32x1_ASAP7_75t_L g143 ( .A1(n_18), .A2(n_144), .A3(n_147), .B1(n_158), .B2(n_162), .Y(n_143) );
AO32x2_ASAP7_75t_L g275 ( .A1(n_18), .A2(n_144), .A3(n_147), .B1(n_158), .B2(n_162), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_19), .B(n_576), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_20), .B(n_162), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_21), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_23), .A2(n_29), .B1(n_516), .B2(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_23), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_24), .A2(n_44), .B1(n_193), .B2(n_194), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_25), .A2(n_92), .B1(n_152), .B2(n_154), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_26), .B(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g498 ( .A(n_27), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_28), .Y(n_555) );
INVx1_ASAP7_75t_L g517 ( .A(n_29), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_30), .B(n_170), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_31), .A2(n_65), .B1(n_154), .B2(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_32), .B(n_156), .Y(n_591) );
INVx2_ASAP7_75t_L g129 ( .A(n_33), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_34), .B(n_157), .Y(n_600) );
INVx1_ASAP7_75t_L g112 ( .A(n_35), .Y(n_112) );
BUFx3_ASAP7_75t_L g880 ( .A(n_35), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_36), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_37), .B(n_558), .Y(n_606) );
AND2x2_ASAP7_75t_L g557 ( .A(n_39), .B(n_558), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_40), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_41), .B(n_202), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_42), .B(n_576), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_43), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_45), .A2(n_104), .B1(n_118), .B2(n_889), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_46), .B(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g253 ( .A1(n_47), .A2(n_78), .B1(n_170), .B2(n_202), .Y(n_253) );
OAI22xp5_ASAP7_75t_SL g513 ( .A1(n_48), .A2(n_514), .B1(n_515), .B2(n_518), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_48), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_49), .B(n_214), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_50), .A2(n_148), .B(n_199), .C(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_51), .A2(n_80), .B1(n_152), .B2(n_156), .Y(n_263) );
INVx1_ASAP7_75t_L g146 ( .A(n_52), .Y(n_146) );
AND2x4_ASAP7_75t_L g160 ( .A(n_53), .B(n_161), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_54), .A2(n_55), .B1(n_154), .B2(n_194), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_56), .B(n_162), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_57), .B(n_558), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_58), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_59), .B(n_154), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_60), .B(n_152), .Y(n_241) );
INVx1_ASAP7_75t_L g161 ( .A(n_61), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_62), .B(n_162), .Y(n_248) );
A2O1A1Ixp33_ASAP7_75t_L g198 ( .A1(n_63), .A2(n_174), .B(n_199), .C(n_200), .Y(n_198) );
NAND3xp33_ASAP7_75t_L g247 ( .A(n_64), .B(n_152), .C(n_246), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_66), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_67), .B(n_162), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_68), .B(n_534), .Y(n_574) );
AND2x2_ASAP7_75t_L g204 ( .A(n_69), .B(n_205), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_70), .Y(n_217) );
NAND3xp33_ASAP7_75t_L g601 ( .A(n_71), .B(n_157), .C(n_193), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_72), .A2(n_95), .B1(n_156), .B2(n_202), .Y(n_255) );
INVx2_ASAP7_75t_L g150 ( .A(n_73), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_74), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_75), .B(n_534), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_76), .B(n_197), .Y(n_563) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_77), .B(n_156), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_79), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_81), .B(n_230), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_82), .Y(n_120) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_83), .A2(n_91), .B1(n_576), .B2(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_85), .B(n_156), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_86), .B(n_246), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g567 ( .A(n_87), .B(n_243), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_88), .B(n_226), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_89), .A2(n_102), .B1(n_154), .B2(n_194), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_90), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_93), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_94), .B(n_182), .Y(n_181) );
NAND2xp33_ASAP7_75t_L g535 ( .A(n_96), .B(n_243), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_97), .B(n_558), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g564 ( .A(n_98), .B(n_197), .C(n_243), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_99), .B(n_534), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_100), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g579 ( .A(n_101), .B(n_576), .Y(n_579) );
BUFx12f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx6_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx11_ASAP7_75t_R g890 ( .A(n_106), .Y(n_890) );
NAND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_109), .Y(n_123) );
NOR2x1_ASAP7_75t_L g888 ( .A(n_109), .B(n_880), .Y(n_888) );
NOR2x1p5_ASAP7_75t_L g110 ( .A(n_111), .B(n_113), .Y(n_110) );
AND3x2_ASAP7_75t_L g122 ( .A(n_111), .B(n_114), .C(n_123), .Y(n_122) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g508 ( .A(n_112), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_114), .Y(n_520) );
BUFx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g874 ( .A(n_115), .Y(n_874) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_124), .Y(n_118) );
INVxp67_ASAP7_75t_L g500 ( .A(n_119), .Y(n_500) );
AOI211xp5_ASAP7_75t_L g501 ( .A1(n_119), .A2(n_133), .B(n_497), .C(n_502), .Y(n_501) );
NOR2xp67_ASAP7_75t_SL g119 ( .A(n_120), .B(n_121), .Y(n_119) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx4_ASAP7_75t_L g496 ( .A(n_122), .Y(n_496) );
AND2x6_ASAP7_75t_SL g506 ( .A(n_123), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_123), .B(n_879), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_511), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_130), .Y(n_125) );
BUFx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g877 ( .A(n_129), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_129), .B(n_886), .Y(n_885) );
OAI21xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_501), .B(n_503), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_494), .Y(n_131) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_132), .A2(n_133), .B1(n_504), .B2(n_509), .Y(n_503) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OA22x2_ASAP7_75t_L g519 ( .A1(n_134), .A2(n_520), .B1(n_521), .B2(n_872), .Y(n_519) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_381), .Y(n_134) );
AND4x1_ASAP7_75t_L g135 ( .A(n_136), .B(n_290), .C(n_328), .D(n_366), .Y(n_135) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_268), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_207), .B(n_218), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_140), .B(n_163), .Y(n_139) );
NAND2xp5_ASAP7_75t_R g339 ( .A(n_140), .B(n_287), .Y(n_339) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g440 ( .A(n_142), .B(n_318), .Y(n_440) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OR2x2_ASAP7_75t_L g209 ( .A(n_143), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g301 ( .A(n_143), .Y(n_301) );
AND2x2_ASAP7_75t_L g315 ( .A(n_143), .B(n_210), .Y(n_315) );
INVx4_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
INVx2_ASAP7_75t_SL g166 ( .A(n_144), .Y(n_166) );
BUFx3_ASAP7_75t_L g211 ( .A(n_144), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_144), .B(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g221 ( .A(n_144), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_144), .B(n_266), .Y(n_265) );
AND2x4_ASAP7_75t_SL g540 ( .A(n_144), .B(n_234), .Y(n_540) );
INVx1_ASAP7_75t_SL g560 ( .A(n_144), .Y(n_560) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B1(n_155), .B2(n_157), .Y(n_147) );
O2A1O1Ixp5_ASAP7_75t_L g223 ( .A1(n_148), .A2(n_224), .B(n_225), .C(n_227), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_148), .A2(n_533), .B(n_535), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_148), .A2(n_566), .B(n_567), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_148), .A2(n_574), .B(n_575), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_148), .A2(n_590), .B(n_591), .Y(n_589) );
BUFx4f_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g246 ( .A(n_149), .Y(n_246) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx8_ASAP7_75t_L g157 ( .A(n_150), .Y(n_157) );
INVx2_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
INVx1_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
INVx2_ASAP7_75t_SL g170 ( .A(n_152), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_152), .B(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_153), .Y(n_154) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_153), .Y(n_156) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_153), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_153), .Y(n_194) );
INVx1_ASAP7_75t_L g199 ( .A(n_153), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_153), .Y(n_202) );
INVx1_ASAP7_75t_L g226 ( .A(n_153), .Y(n_226) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_153), .Y(n_243) );
INVx3_ASAP7_75t_L g534 ( .A(n_153), .Y(n_534) );
INVx1_ASAP7_75t_L g577 ( .A(n_153), .Y(n_577) );
INVx2_ASAP7_75t_L g172 ( .A(n_154), .Y(n_172) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_154), .A2(n_534), .B1(n_555), .B2(n_556), .Y(n_554) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_154), .A2(n_600), .B(n_601), .Y(n_599) );
INVx2_ASAP7_75t_L g613 ( .A(n_154), .Y(n_613) );
INVx3_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_156), .A2(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g605 ( .A(n_156), .Y(n_605) );
INVx6_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_157), .A2(n_241), .B(n_242), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g262 ( .A1(n_157), .A2(n_180), .B1(n_263), .B2(n_264), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_157), .A2(n_593), .B(n_594), .Y(n_592) );
O2A1O1Ixp5_ASAP7_75t_L g621 ( .A1(n_157), .A2(n_225), .B(n_622), .C(n_623), .Y(n_621) );
OAI21x1_ASAP7_75t_L g167 ( .A1(n_158), .A2(n_168), .B(n_176), .Y(n_167) );
INVx2_ASAP7_75t_SL g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_SL g256 ( .A(n_159), .Y(n_256) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_160), .A2(n_211), .A3(n_212), .B(n_216), .Y(n_210) );
BUFx10_ASAP7_75t_L g234 ( .A(n_160), .Y(n_234) );
BUFx10_ASAP7_75t_L g547 ( .A(n_160), .Y(n_547) );
INVx2_ASAP7_75t_L g261 ( .A(n_162), .Y(n_261) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_185), .Y(n_163) );
BUFx2_ASAP7_75t_L g208 ( .A(n_164), .Y(n_208) );
AND2x2_ASAP7_75t_L g273 ( .A(n_164), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g288 ( .A(n_164), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_164), .B(n_210), .Y(n_305) );
INVx3_ASAP7_75t_L g318 ( .A(n_164), .Y(n_318) );
AND2x2_ASAP7_75t_L g353 ( .A(n_164), .B(n_275), .Y(n_353) );
INVx2_ASAP7_75t_L g365 ( .A(n_164), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_164), .Y(n_369) );
INVxp67_ASAP7_75t_L g406 ( .A(n_164), .Y(n_406) );
OR2x2_ASAP7_75t_L g419 ( .A(n_164), .B(n_302), .Y(n_419) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
OAI21x1_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_181), .Y(n_165) );
AOI21x1_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_173), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_172), .A2(n_245), .B(n_247), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_173), .A2(n_180), .B1(n_213), .B2(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_173), .A2(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g553 ( .A(n_174), .Y(n_553) );
BUFx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g231 ( .A(n_175), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_180), .Y(n_176) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_180), .A2(n_253), .B1(n_254), .B2(n_255), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_180), .A2(n_553), .B1(n_612), .B2(n_614), .Y(n_611) );
INVx2_ASAP7_75t_L g188 ( .A(n_182), .Y(n_188) );
NOR2xp67_ASAP7_75t_SL g545 ( .A(n_182), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AO31x2_ASAP7_75t_L g610 ( .A1(n_183), .A2(n_547), .A3(n_611), .B(n_615), .Y(n_610) );
INVx2_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g206 ( .A(n_184), .Y(n_206) );
INVx2_ASAP7_75t_L g238 ( .A(n_184), .Y(n_238) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g271 ( .A(n_186), .Y(n_271) );
INVx1_ASAP7_75t_L g358 ( .A(n_186), .Y(n_358) );
AND2x2_ASAP7_75t_L g373 ( .A(n_186), .B(n_210), .Y(n_373) );
INVx1_ASAP7_75t_L g388 ( .A(n_186), .Y(n_388) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g302 ( .A(n_187), .Y(n_302) );
AOI21x1_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_204), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_198), .B(n_203), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_191), .B(n_196), .Y(n_190) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B1(n_194), .B2(n_195), .Y(n_191) );
INVx2_ASAP7_75t_L g214 ( .A(n_193), .Y(n_214) );
INVx1_ASAP7_75t_L g232 ( .A(n_194), .Y(n_232) );
AOI21x1_ASAP7_75t_L g602 ( .A1(n_196), .A2(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_SL g254 ( .A(n_197), .Y(n_254) );
INVx1_ASAP7_75t_L g538 ( .A(n_199), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_206), .B(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_206), .B(n_616), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_207), .A2(n_477), .B1(n_479), .B2(n_481), .Y(n_476) );
OR2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_208), .B(n_357), .Y(n_434) );
BUFx2_ASAP7_75t_L g448 ( .A(n_208), .Y(n_448) );
AND2x2_ASAP7_75t_L g466 ( .A(n_208), .B(n_322), .Y(n_466) );
INVx2_ASAP7_75t_L g348 ( .A(n_209), .Y(n_348) );
OR2x2_ASAP7_75t_L g364 ( .A(n_209), .B(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g272 ( .A(n_210), .Y(n_272) );
AND2x2_ASAP7_75t_L g357 ( .A(n_210), .B(n_358), .Y(n_357) );
AO31x2_ASAP7_75t_L g251 ( .A1(n_211), .A2(n_252), .A3(n_256), .B(n_257), .Y(n_251) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_249), .Y(n_218) );
OR2x2_ASAP7_75t_L g413 ( .A(n_219), .B(n_370), .Y(n_413) );
OR2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_236), .Y(n_219) );
AND2x2_ASAP7_75t_L g284 ( .A(n_220), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g325 ( .A(n_220), .Y(n_325) );
INVx2_ASAP7_75t_SL g333 ( .A(n_220), .Y(n_333) );
BUFx2_ASAP7_75t_L g345 ( .A(n_220), .Y(n_345) );
OR2x2_ASAP7_75t_L g433 ( .A(n_220), .B(n_251), .Y(n_433) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_235), .Y(n_220) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_221), .A2(n_222), .B(n_235), .Y(n_298) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_221), .A2(n_588), .B(n_595), .Y(n_587) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_221), .A2(n_598), .B(n_606), .Y(n_597) );
OAI21x1_ASAP7_75t_L g652 ( .A1(n_221), .A2(n_588), .B(n_595), .Y(n_652) );
OA21x2_ASAP7_75t_L g655 ( .A1(n_221), .A2(n_598), .B(n_606), .Y(n_655) );
OAI21x1_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_228), .B(n_234), .Y(n_222) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_231), .B1(n_232), .B2(n_233), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_230), .A2(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_231), .A2(n_537), .B1(n_538), .B2(n_539), .Y(n_536) );
OAI21x1_ASAP7_75t_L g239 ( .A1(n_234), .A2(n_240), .B(n_244), .Y(n_239) );
AOI31xp67_ASAP7_75t_L g260 ( .A1(n_234), .A2(n_261), .A3(n_262), .B(n_265), .Y(n_260) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_234), .A2(n_562), .B(n_565), .Y(n_561) );
OAI21x1_ASAP7_75t_L g572 ( .A1(n_234), .A2(n_573), .B(n_578), .Y(n_572) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_234), .A2(n_589), .B(n_592), .Y(n_588) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_234), .A2(n_599), .B(n_602), .Y(n_598) );
OAI21x1_ASAP7_75t_L g620 ( .A1(n_234), .A2(n_621), .B(n_624), .Y(n_620) );
AND2x2_ASAP7_75t_L g277 ( .A(n_236), .B(n_259), .Y(n_277) );
AND2x2_ASAP7_75t_L g313 ( .A(n_236), .B(n_298), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_239), .B(n_248), .Y(n_236) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_237), .A2(n_239), .B(n_248), .Y(n_283) );
OAI21xp33_ASAP7_75t_SL g571 ( .A1(n_237), .A2(n_572), .B(n_581), .Y(n_571) );
OAI21x1_ASAP7_75t_L g619 ( .A1(n_237), .A2(n_620), .B(n_628), .Y(n_619) );
OAI21x1_ASAP7_75t_L g643 ( .A1(n_237), .A2(n_572), .B(n_581), .Y(n_643) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_237), .A2(n_620), .B(n_628), .Y(n_703) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g558 ( .A(n_238), .Y(n_558) );
INVx2_ASAP7_75t_L g627 ( .A(n_243), .Y(n_627) );
INVx1_ASAP7_75t_L g351 ( .A(n_249), .Y(n_351) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_250), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g457 ( .A(n_250), .B(n_437), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_250), .B(n_280), .Y(n_481) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_259), .Y(n_250) );
INVx1_ASAP7_75t_L g285 ( .A(n_251), .Y(n_285) );
INVx2_ASAP7_75t_L g295 ( .A(n_251), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_251), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g324 ( .A(n_251), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g338 ( .A(n_251), .B(n_298), .Y(n_338) );
OR2x2_ASAP7_75t_L g370 ( .A(n_251), .B(n_310), .Y(n_370) );
INVx1_ASAP7_75t_L g454 ( .A(n_251), .Y(n_454) );
AND2x2_ASAP7_75t_L g297 ( .A(n_259), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g335 ( .A(n_259), .Y(n_335) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g311 ( .A(n_260), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_267), .Y(n_266) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_276), .B1(n_278), .B2(n_286), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g415 ( .A(n_271), .Y(n_415) );
INVx1_ASAP7_75t_L g289 ( .A(n_272), .Y(n_289) );
AND2x4_ASAP7_75t_L g322 ( .A(n_272), .B(n_275), .Y(n_322) );
AND2x2_ASAP7_75t_L g431 ( .A(n_272), .B(n_302), .Y(n_431) );
AND2x2_ASAP7_75t_L g483 ( .A(n_273), .B(n_357), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_273), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g337 ( .A(n_277), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g470 ( .A(n_277), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_284), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_280), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g389 ( .A(n_280), .Y(n_389) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g455 ( .A(n_281), .Y(n_455) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g342 ( .A(n_282), .Y(n_342) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g327 ( .A(n_283), .B(n_311), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_284), .B(n_326), .Y(n_442) );
AND2x2_ASAP7_75t_L g334 ( .A(n_285), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx1_ASAP7_75t_L g474 ( .A(n_289), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_299), .B1(n_306), .B2(n_314), .C(n_319), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
AND2x2_ASAP7_75t_L g392 ( .A(n_293), .B(n_313), .Y(n_392) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_294), .B(n_313), .Y(n_361) );
OR2x2_ASAP7_75t_L g376 ( .A(n_294), .B(n_327), .Y(n_376) );
INVx2_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g341 ( .A(n_295), .B(n_342), .Y(n_341) );
INVxp67_ASAP7_75t_L g452 ( .A(n_297), .Y(n_452) );
INVx1_ASAP7_75t_L g412 ( .A(n_298), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
AND2x2_ASAP7_75t_L g472 ( .A(n_300), .B(n_473), .Y(n_472) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g426 ( .A(n_301), .B(n_388), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_302), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g347 ( .A(n_302), .Y(n_347) );
INVx1_ASAP7_75t_L g399 ( .A(n_302), .Y(n_399) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_307), .A2(n_333), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g362 ( .A(n_309), .B(n_345), .Y(n_362) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_309), .Y(n_402) );
AND2x2_ASAP7_75t_L g486 ( .A(n_309), .B(n_423), .Y(n_486) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g493 ( .A(n_312), .B(n_410), .Y(n_493) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
INVx2_ASAP7_75t_SL g394 ( .A(n_315), .Y(n_394) );
AND2x2_ASAP7_75t_L g398 ( .A(n_315), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g458 ( .A(n_315), .B(n_318), .Y(n_458) );
AND2x2_ASAP7_75t_L g480 ( .A(n_315), .B(n_405), .Y(n_480) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g377 ( .A(n_318), .B(n_322), .Y(n_377) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g371 ( .A(n_322), .B(n_347), .Y(n_371) );
AND2x2_ASAP7_75t_L g404 ( .A(n_322), .B(n_405), .Y(n_404) );
INVx3_ASAP7_75t_L g421 ( .A(n_322), .Y(n_421) );
INVx1_ASAP7_75t_L g490 ( .A(n_323), .Y(n_490) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
AND2x4_ASAP7_75t_L g354 ( .A(n_324), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g396 ( .A(n_326), .B(n_345), .Y(n_396) );
AND2x2_ASAP7_75t_L g422 ( .A(n_326), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g432 ( .A(n_327), .B(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_329), .B(n_349), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_336), .B(n_339), .C(n_340), .Y(n_329) );
INVx2_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_332), .B(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_333), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_333), .B(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_334), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g355 ( .A(n_335), .B(n_342), .Y(n_355) );
INVx1_ASAP7_75t_L g410 ( .A(n_335), .Y(n_410) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B(n_346), .Y(n_340) );
NAND2x1p5_ASAP7_75t_L g411 ( .A(n_342), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g423 ( .A(n_345), .Y(n_423) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x4_ASAP7_75t_L g447 ( .A(n_348), .B(n_415), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_359), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_352), .B(n_354), .C(n_356), .Y(n_350) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g414 ( .A(n_353), .B(n_415), .Y(n_414) );
BUFx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OAI21xp5_ASAP7_75t_SL g359 ( .A1(n_360), .A2(n_362), .B(n_363), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_365), .Y(n_374) );
OR2x2_ASAP7_75t_L g393 ( .A(n_365), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g475 ( .A(n_365), .Y(n_475) );
AOI222xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B1(n_372), .B2(n_375), .C1(n_377), .C2(n_378), .Y(n_366) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_368), .B(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_369), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g380 ( .A(n_370), .Y(n_380) );
INVx1_ASAP7_75t_L g478 ( .A(n_370), .Y(n_478) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_373), .B(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g456 ( .A(n_373), .Y(n_456) );
AND2x4_ASAP7_75t_L g463 ( .A(n_373), .B(n_440), .Y(n_463) );
INVx2_ASAP7_75t_L g492 ( .A(n_373), .Y(n_492) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI22xp33_ASAP7_75t_L g428 ( .A1(n_376), .A2(n_429), .B1(n_432), .B2(n_434), .Y(n_428) );
AOI211xp5_ASAP7_75t_L g482 ( .A1(n_378), .A2(n_483), .B(n_484), .C(n_488), .Y(n_482) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NOR2xp67_ASAP7_75t_SL g381 ( .A(n_382), .B(n_443), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_400), .C(n_407), .D(n_427), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_389), .B(n_390), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_393), .B1(n_395), .B2(n_397), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_394), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_395), .B(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g405 ( .A(n_399), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g430 ( .A(n_406), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_414), .B1(n_416), .B2(n_422), .C(n_424), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_413), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_409), .B(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
AND2x2_ASAP7_75t_L g462 ( .A(n_410), .B(n_437), .Y(n_462) );
INVx2_ASAP7_75t_L g437 ( .A(n_411), .Y(n_437) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
NAND2x1_ASAP7_75t_SL g417 ( .A(n_418), .B(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g487 ( .A(n_418), .Y(n_487) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g489 ( .A(n_426), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_435), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx1_ASAP7_75t_L g471 ( .A(n_433), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B1(n_441), .B2(n_442), .Y(n_435) );
AND2x2_ASAP7_75t_L g468 ( .A(n_437), .B(n_454), .Y(n_468) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g449 ( .A(n_442), .Y(n_449) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_459), .C(n_482), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_449), .B1(n_450), .B2(n_456), .C1(n_457), .C2(n_458), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_446), .B(n_448), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AOI211xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_463), .B(n_464), .C(n_476), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_467), .B1(n_469), .B2(n_472), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B1(n_491), .B2(n_493), .Y(n_488) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_497), .B(n_500), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_495), .Y(n_502) );
INVx1_ASAP7_75t_L g510 ( .A(n_497), .Y(n_510) );
BUFx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AOI21xp33_ASAP7_75t_SL g511 ( .A1(n_512), .A2(n_875), .B(n_881), .Y(n_511) );
XNOR2x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_752), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_523), .B(n_660), .C(n_711), .Y(n_522) );
OAI211xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_582), .B(n_629), .C(n_647), .Y(n_523) );
NAND3x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_541), .C(n_569), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g720 ( .A(n_526), .B(n_699), .Y(n_720) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND3x2_ASAP7_75t_L g640 ( .A(n_527), .B(n_641), .C(n_645), .Y(n_640) );
AND2x2_ASAP7_75t_L g675 ( .A(n_527), .B(n_659), .Y(n_675) );
AND2x2_ASAP7_75t_L g681 ( .A(n_527), .B(n_677), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_527), .B(n_645), .Y(n_822) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g724 ( .A(n_528), .B(n_645), .Y(n_724) );
AND2x2_ASAP7_75t_L g735 ( .A(n_528), .B(n_689), .Y(n_735) );
BUFx2_ASAP7_75t_L g741 ( .A(n_528), .Y(n_741) );
NAND2x1_ASAP7_75t_L g757 ( .A(n_528), .B(n_758), .Y(n_757) );
OR2x2_ASAP7_75t_L g763 ( .A(n_528), .B(n_764), .Y(n_763) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g657 ( .A(n_529), .Y(n_657) );
AND2x2_ASAP7_75t_L g688 ( .A(n_529), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g708 ( .A(n_529), .B(n_644), .Y(n_708) );
INVx1_ASAP7_75t_L g779 ( .A(n_529), .Y(n_779) );
AND2x4_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
OAI21x1_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_536), .B(n_540), .Y(n_531) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OR2x6_ASAP7_75t_L g756 ( .A(n_542), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g658 ( .A(n_543), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_543), .B(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_559), .Y(n_543) );
INVx2_ASAP7_75t_L g646 ( .A(n_544), .Y(n_646) );
INVx1_ASAP7_75t_L g700 ( .A(n_544), .Y(n_700) );
AOI21x1_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B(n_557), .Y(n_544) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g644 ( .A(n_559), .Y(n_644) );
INVx2_ASAP7_75t_L g678 ( .A(n_559), .Y(n_678) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_561), .B(n_568), .Y(n_559) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_570), .A2(n_860), .B(n_864), .Y(n_859) );
BUFx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g699 ( .A(n_571), .B(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_607), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_SL g855 ( .A(n_584), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp67_ASAP7_75t_L g585 ( .A(n_586), .B(n_596), .Y(n_585) );
INVx3_ASAP7_75t_L g637 ( .A(n_586), .Y(n_637) );
AND2x2_ASAP7_75t_L g784 ( .A(n_586), .B(n_597), .Y(n_784) );
BUFx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g673 ( .A(n_587), .Y(n_673) );
AND2x4_ASAP7_75t_L g638 ( .A(n_596), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g697 ( .A(n_597), .Y(n_697) );
AND2x2_ASAP7_75t_L g714 ( .A(n_597), .B(n_610), .Y(n_714) );
AND2x2_ASAP7_75t_L g826 ( .A(n_597), .B(n_703), .Y(n_826) );
AND2x2_ASAP7_75t_L g848 ( .A(n_597), .B(n_618), .Y(n_848) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_609), .B(n_617), .Y(n_608) );
INVx1_ASAP7_75t_L g668 ( .A(n_609), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_609), .B(n_858), .Y(n_857) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
OR2x2_ASAP7_75t_L g654 ( .A(n_610), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g672 ( .A(n_610), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g726 ( .A(n_610), .B(n_652), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_610), .B(n_655), .Y(n_768) );
OR2x2_ASAP7_75t_L g838 ( .A(n_610), .B(n_652), .Y(n_838) );
INVx1_ASAP7_75t_L g666 ( .A(n_617), .Y(n_666) );
AND2x4_ASAP7_75t_L g684 ( .A(n_617), .B(n_638), .Y(n_684) );
AND2x2_ASAP7_75t_L g830 ( .A(n_617), .B(n_672), .Y(n_830) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx3_ASAP7_75t_L g632 ( .A(n_618), .Y(n_632) );
AND2x2_ASAP7_75t_L g692 ( .A(n_618), .B(n_651), .Y(n_692) );
INVx1_ASAP7_75t_L g745 ( .A(n_618), .Y(n_745) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_618), .Y(n_783) );
AND2x2_ASAP7_75t_L g786 ( .A(n_618), .B(n_655), .Y(n_786) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_618), .Y(n_796) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI21xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_633), .B(n_640), .Y(n_629) );
AND2x2_ASAP7_75t_L g828 ( .A(n_630), .B(n_733), .Y(n_828) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g695 ( .A(n_631), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_631), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_632), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g775 ( .A(n_632), .B(n_638), .Y(n_775) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_637), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g773 ( .A(n_637), .B(n_714), .Y(n_773) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_637), .Y(n_804) );
INVx2_ASAP7_75t_L g738 ( .A(n_638), .Y(n_738) );
AND2x2_ASAP7_75t_L g867 ( .A(n_639), .B(n_652), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_640), .A2(n_722), .B1(n_723), .B2(n_725), .C(n_727), .Y(n_721) );
AND2x2_ASAP7_75t_L g662 ( .A(n_641), .B(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g723 ( .A(n_641), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx2_ASAP7_75t_L g659 ( .A(n_642), .Y(n_659) );
OR2x2_ASAP7_75t_L g792 ( .A(n_642), .B(n_677), .Y(n_792) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g689 ( .A(n_643), .Y(n_689) );
INVxp67_ASAP7_75t_L g719 ( .A(n_644), .Y(n_719) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g663 ( .A(n_646), .Y(n_663) );
AND2x2_ASAP7_75t_L g676 ( .A(n_646), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g683 ( .A(n_646), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_656), .Y(n_647) );
AND2x2_ASAP7_75t_L g806 ( .A(n_648), .B(n_807), .Y(n_806) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g733 ( .A(n_650), .B(n_714), .Y(n_733) );
HB1xp67_ASAP7_75t_L g863 ( .A(n_650), .Y(n_863) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g691 ( .A(n_653), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g841 ( .A(n_653), .Y(n_841) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g729 ( .A(n_654), .Y(n_729) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_654), .Y(n_803) );
AND2x2_ASAP7_75t_L g702 ( .A(n_655), .B(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_656), .B(n_828), .Y(n_827) );
AND2x4_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
AND2x2_ASAP7_75t_L g698 ( .A(n_657), .B(n_699), .Y(n_698) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_658), .A2(n_680), .B(n_684), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g660 ( .A(n_661), .B(n_679), .C(n_685), .D(n_693), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_664), .B(n_669), .Y(n_661) );
INVx2_ASAP7_75t_L g750 ( .A(n_663), .Y(n_750) );
AND2x2_ASAP7_75t_L g761 ( .A(n_663), .B(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_L g771 ( .A(n_663), .B(n_688), .Y(n_771) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g847 ( .A(n_668), .B(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_674), .Y(n_669) );
INVxp67_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI33xp33_ASAP7_75t_L g817 ( .A1(n_671), .A2(n_708), .A3(n_818), .B1(n_820), .B2(n_823), .B3(n_824), .Y(n_817) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g850 ( .A(n_672), .B(n_702), .Y(n_850) );
BUFx2_ASAP7_75t_L g705 ( .A(n_673), .Y(n_705) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_676), .B(n_688), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_677), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_678), .Y(n_731) );
INVx1_ASAP7_75t_L g764 ( .A(n_678), .Y(n_764) );
AND2x2_ASAP7_75t_L g778 ( .A(n_678), .B(n_779), .Y(n_778) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
AND2x2_ASAP7_75t_L g749 ( .A(n_681), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_SL g801 ( .A(n_681), .Y(n_801) );
INVx1_ASAP7_75t_L g811 ( .A(n_682), .Y(n_811) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g687 ( .A(n_683), .Y(n_687) );
INVx1_ASAP7_75t_L g793 ( .A(n_683), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_690), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
OR2x2_ASAP7_75t_L g776 ( .A(n_687), .B(n_777), .Y(n_776) );
AND2x2_ASAP7_75t_L g747 ( .A(n_688), .B(n_731), .Y(n_747) );
AND2x2_ASAP7_75t_L g710 ( .A(n_689), .B(n_700), .Y(n_710) );
INVx2_ASAP7_75t_L g758 ( .A(n_689), .Y(n_758) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g751 ( .A(n_692), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_698), .B1(n_701), .B2(n_706), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_696), .Y(n_869) );
AOI221xp5_ASAP7_75t_L g780 ( .A1(n_698), .A2(n_781), .B1(n_785), .B2(n_787), .C(n_789), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_699), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g835 ( .A(n_699), .Y(n_835) );
AND2x2_ASAP7_75t_L g854 ( .A(n_699), .B(n_778), .Y(n_854) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g823 ( .A(n_702), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_702), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g809 ( .A(n_703), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_704), .B(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g797 ( .A(n_704), .B(n_738), .Y(n_797) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g851 ( .A1(n_706), .A2(n_852), .B1(n_854), .B2(n_855), .Y(n_851) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_709), .Y(n_707) );
OR2x2_ASAP7_75t_L g868 ( .A(n_709), .B(n_763), .Y(n_868) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g816 ( .A(n_710), .B(n_778), .Y(n_816) );
OAI211xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_715), .B(n_721), .C(n_736), .Y(n_711) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_714), .Y(n_722) );
AND2x2_ASAP7_75t_L g795 ( .A(n_714), .B(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
NAND2x1p5_ASAP7_75t_L g717 ( .A(n_718), .B(n_720), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g788 ( .A(n_720), .Y(n_788) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_726), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g785 ( .A(n_726), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g819 ( .A(n_726), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_726), .B(n_833), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_730), .B1(n_732), .B2(n_734), .Y(n_727) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI21xp33_ASAP7_75t_SL g736 ( .A1(n_737), .A2(n_739), .B(n_742), .Y(n_736) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_746), .B1(n_748), .B2(n_751), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_744), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AOI211xp5_ASAP7_75t_SL g829 ( .A1(n_747), .A2(n_830), .B(n_831), .C(n_839), .Y(n_829) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g844 ( .A(n_750), .B(n_778), .Y(n_844) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_812), .C(n_842), .Y(n_752) );
NAND3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_780), .C(n_800), .Y(n_753) );
O2A1O1Ixp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_759), .B(n_765), .C(n_769), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp33_ASAP7_75t_SL g831 ( .A1(n_757), .A2(n_832), .B1(n_834), .B2(n_836), .Y(n_831) );
INVx1_ASAP7_75t_SL g821 ( .A(n_758), .Y(n_821) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
OR2x2_ASAP7_75t_L g834 ( .A(n_763), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_772), .B1(n_774), .B2(n_776), .Y(n_769) );
NAND2xp33_ASAP7_75t_SL g787 ( .A(n_770), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g853 ( .A(n_775), .Y(n_853) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g807 ( .A(n_778), .B(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_782), .B(n_816), .Y(n_815) );
AND2x4_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g858 ( .A(n_783), .Y(n_858) );
INVx1_ASAP7_75t_L g833 ( .A(n_786), .Y(n_833) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_794), .B1(n_797), .B2(n_798), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NOR2x1p5_ASAP7_75t_SL g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx1_ASAP7_75t_L g799 ( .A(n_792), .Y(n_799) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g805 ( .A(n_796), .Y(n_805) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B(n_806), .C(n_810), .Y(n_800) );
NOR3x1_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .C(n_805), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_807), .B(n_862), .Y(n_861) );
AND2x2_ASAP7_75t_L g866 ( .A(n_808), .B(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND3xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_827), .C(n_829), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_814), .B(n_817), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
BUFx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp67_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
INVx1_ASAP7_75t_L g871 ( .A(n_840), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_851), .C(n_859), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVxp67_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVxp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVxp67_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVxp67_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_868), .B1(n_869), .B2(n_870), .Y(n_864) );
INVx2_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx4_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g887 ( .A(n_874), .B(n_888), .Y(n_887) );
BUFx6f_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
AND2x6_ASAP7_75t_SL g876 ( .A(n_877), .B(n_878), .Y(n_876) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .Y(n_881) );
INVx5_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
BUFx10_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_890), .Y(n_889) );
endmodule