module real_jpeg_18779_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_288;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_184;
wire n_164;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx3_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_0),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_1),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_1),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_1),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_2),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_7),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_3),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_4),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_4),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_109),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

AOI31xp33_ASAP7_75t_SL g47 ( 
.A1(n_7),
.A2(n_48),
.A3(n_52),
.B(n_56),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_7),
.B(n_85),
.Y(n_84)
);

NAND2x1_ASAP7_75t_SL g95 ( 
.A(n_7),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_7),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_7),
.B(n_82),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_7),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_7),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_25),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_8),
.B(n_72),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_8),
.B(n_102),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_8),
.Y(n_124)
);

NAND2x1_ASAP7_75t_SL g143 ( 
.A(n_8),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_8),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_9),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_9),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_9),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_9),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_9),
.B(n_68),
.Y(n_223)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_10),
.Y(n_126)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_10),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_11),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_11),
.B(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_13),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_13),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_13),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_13),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_13),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_13),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_13),
.B(n_263),
.Y(n_262)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

BUFx8_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_184),
.B1(n_287),
.B2(n_288),
.Y(n_17)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_18),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_182),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_138),
.Y(n_19)
);

NOR2x1_ASAP7_75t_L g183 ( 
.A(n_20),
.B(n_138),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_74),
.C(n_114),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_21),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_46),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_22),
.B(n_47),
.C(n_61),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_33),
.C(n_40),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_23),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_24),
.B(n_28),
.Y(n_222)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_24),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_24),
.A2(n_247),
.B1(n_248),
.B2(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_31),
.Y(n_205)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_34),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_274)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_61),
.Y(n_46)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_50),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_56),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_56),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_62),
.B(n_67),
.C(n_71),
.Y(n_181)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_71),
.B(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_71),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_74),
.B(n_114),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_89),
.C(n_106),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_75),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_81),
.C(n_84),
.Y(n_136)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_78),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_88),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_81),
.B(n_236),
.C(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_81),
.A2(n_88),
.B1(n_238),
.B2(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_90),
.B(n_107),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_95),
.C(n_100),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_91),
.A2(n_100),
.B1(n_101),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_91),
.Y(n_229)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2x2_ASAP7_75t_L g227 ( 
.A(n_95),
.B(n_228),
.Y(n_227)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_100),
.A2(n_101),
.B1(n_162),
.B2(n_167),
.Y(n_161)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_135),
.Y(n_114)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_127),
.C(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B1(n_133),
.B2(n_134),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_123),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_137),
.C(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_154),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

XNOR2x1_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_150),
.Y(n_141)
);

XNOR2x2_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_168),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_181),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_173),
.B1(n_179),
.B2(n_180),
.Y(n_169)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_170),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_184),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_282),
.B(n_286),
.Y(n_185)
);

AOI21x1_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_268),
.B(n_281),
.Y(n_186)
);

OAI21x1_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_230),
.B(n_267),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_218),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_189),
.B(n_218),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_197),
.C(n_206),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_190),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_196),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_196),
.C(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_198),
.B1(n_206),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_199),
.B(n_203),
.Y(n_237)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_206)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_212),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_216),
.Y(n_220)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_213),
.Y(n_250)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_262),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_219),
.B(n_225),
.C(n_227),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_222),
.C(n_223),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

AOI21x1_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_241),
.B(n_266),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_235),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_237),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_251),
.B(n_265),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_261),
.B(n_264),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_259),
.Y(n_264)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_280),
.Y(n_268)
);

NOR2x1p5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_280),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_277),
.B2(n_278),
.Y(n_269)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_276),
.C(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_284),
.Y(n_286)
);


endmodule