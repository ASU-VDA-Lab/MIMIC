module fake_jpeg_1619_n_486 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_486);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_486;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_0),
.B(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_33),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_60),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_61),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_22),
.B(n_12),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_91),
.Y(n_115)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_69),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_16),
.Y(n_70)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_74),
.Y(n_157)
);

BUFx12f_ASAP7_75t_SL g75 ( 
.A(n_26),
.Y(n_75)
);

BUFx2_ASAP7_75t_R g151 ( 
.A(n_75),
.Y(n_151)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_80),
.Y(n_133)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_82),
.Y(n_153)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_85),
.Y(n_163)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_22),
.B(n_10),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_100),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_14),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_94),
.Y(n_123)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_10),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_16),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx6_ASAP7_75t_SL g150 ( 
.A(n_95),
.Y(n_150)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_18),
.B(n_28),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_102),
.Y(n_127)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_23),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_16),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_25),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_18),
.B(n_10),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_37),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_47),
.B1(n_38),
.B2(n_28),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_105),
.A2(n_110),
.B1(n_113),
.B2(n_124),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_53),
.A2(n_47),
.B1(n_48),
.B2(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_21),
.B1(n_47),
.B2(n_44),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_55),
.A2(n_48),
.B1(n_34),
.B2(n_39),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_62),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_70),
.B1(n_43),
.B2(n_36),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_73),
.B(n_35),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_134),
.B(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_17),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_141),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_88),
.B(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_145),
.B(n_0),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_84),
.B(n_20),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_37),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_59),
.Y(n_181)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_104),
.B(n_43),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_166),
.B(n_179),
.Y(n_232)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_194),
.B1(n_195),
.B2(n_203),
.Y(n_229)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_146),
.Y(n_169)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_169),
.Y(n_234)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_170),
.Y(n_240)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_112),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_171),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_60),
.B1(n_76),
.B2(n_77),
.Y(n_173)
);

AO22x2_ASAP7_75t_SL g247 ( 
.A1(n_173),
.A2(n_178),
.B1(n_199),
.B2(n_200),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_177),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_113),
.A2(n_63),
.B1(n_71),
.B2(n_72),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_31),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_119),
.Y(n_180)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_188),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_106),
.B(n_30),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_182),
.B(n_190),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_114),
.A2(n_21),
.B1(n_36),
.B2(n_25),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_183),
.A2(n_201),
.B1(n_207),
.B2(n_210),
.Y(n_230)
);

NAND2x2_ASAP7_75t_SL g185 ( 
.A(n_141),
.B(n_16),
.Y(n_185)
);

OAI22x1_ASAP7_75t_R g233 ( 
.A1(n_185),
.A2(n_125),
.B1(n_133),
.B2(n_129),
.Y(n_233)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_114),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_120),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_108),
.B(n_99),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_193),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_123),
.B(n_94),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_101),
.B1(n_100),
.B2(n_82),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_128),
.B1(n_144),
.B2(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_138),
.B(n_95),
.C(n_78),
.Y(n_197)
);

OAI32xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_208),
.A3(n_149),
.B1(n_40),
.B2(n_107),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_162),
.A2(n_81),
.B1(n_50),
.B2(n_80),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_95),
.B1(n_80),
.B2(n_40),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_123),
.A2(n_16),
.B1(n_40),
.B2(n_42),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_160),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_122),
.A2(n_40),
.B1(n_42),
.B2(n_27),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_204),
.Y(n_214)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_117),
.A2(n_40),
.B1(n_27),
.B2(n_3),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_143),
.B(n_1),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_150),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_126),
.Y(n_211)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_212),
.B(n_238),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_165),
.B(n_111),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_225),
.B(n_210),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_175),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_185),
.A2(n_133),
.B(n_129),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_231),
.A2(n_237),
.B(n_245),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_R g267 ( 
.A(n_233),
.B(n_190),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_185),
.A2(n_158),
.B(n_125),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_172),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_184),
.A2(n_126),
.B1(n_118),
.B2(n_112),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_244),
.A2(n_178),
.B1(n_173),
.B2(n_199),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_185),
.A2(n_140),
.B(n_109),
.Y(n_245)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_181),
.B1(n_166),
.B2(n_174),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_249),
.A2(n_251),
.B1(n_260),
.B2(n_262),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_250),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_220),
.A2(n_181),
.B1(n_208),
.B2(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_218),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_224),
.Y(n_253)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_254),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_216),
.B(n_228),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_257),
.A2(n_243),
.B(n_247),
.Y(n_293)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_258),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_182),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_259),
.B(n_261),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_220),
.A2(n_175),
.B1(n_192),
.B2(n_179),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_232),
.B(n_189),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_193),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_263),
.Y(n_283)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_197),
.C(n_193),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_265),
.B(n_206),
.C(n_169),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_270),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_268),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_269),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_223),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_235),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_271),
.A2(n_213),
.B1(n_204),
.B2(n_243),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_216),
.A2(n_170),
.B(n_177),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_274),
.A2(n_188),
.B(n_240),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_229),
.A2(n_200),
.B1(n_196),
.B2(n_122),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_247),
.B1(n_240),
.B2(n_219),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_167),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_276),
.B(n_223),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_233),
.B(n_244),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_278),
.A2(n_274),
.B1(n_270),
.B2(n_254),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_247),
.B1(n_230),
.B2(n_233),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_285),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_215),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_280),
.B(n_263),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_284),
.A2(n_267),
.B1(n_276),
.B2(n_262),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_286),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_293),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_205),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_296),
.C(n_303),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_239),
.B(n_235),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_295),
.A2(n_273),
.B(n_250),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_297),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_239),
.B1(n_242),
.B2(n_186),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_298),
.A2(n_263),
.B1(n_264),
.B2(n_248),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_272),
.Y(n_299)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_187),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_251),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_309),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_260),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_332),
.C(n_283),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_261),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_310),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_332),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_290),
.B(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_314),
.B(n_318),
.Y(n_342)
);

XNOR2x1_ASAP7_75t_L g316 ( 
.A(n_303),
.B(n_263),
.Y(n_316)
);

XNOR2x1_ASAP7_75t_L g334 ( 
.A(n_316),
.B(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_321),
.B1(n_324),
.B2(n_330),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_287),
.A2(n_275),
.B1(n_249),
.B2(n_256),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_322),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_287),
.A2(n_275),
.B1(n_257),
.B2(n_255),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_285),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_302),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_213),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_326),
.B(n_271),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_327),
.A2(n_286),
.B1(n_279),
.B2(n_278),
.Y(n_337)
);

AOI221xp5_ASAP7_75t_L g328 ( 
.A1(n_291),
.A2(n_252),
.B1(n_253),
.B2(n_268),
.C(n_274),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_325),
.Y(n_339)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_288),
.Y(n_329)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_329),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_291),
.A2(n_264),
.B1(n_258),
.B2(n_271),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_331),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_191),
.C(n_209),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_334),
.B(n_335),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_307),
.B(n_290),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_343),
.C(n_353),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_337),
.A2(n_339),
.B1(n_350),
.B2(n_357),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_307),
.B(n_283),
.CI(n_295),
.CON(n_338),
.SN(n_338)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_311),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_293),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_340),
.B(n_341),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_316),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_302),
.C(n_281),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_313),
.B(n_324),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_347),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_348),
.B(n_359),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_284),
.B1(n_278),
.B2(n_281),
.Y(n_350)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_289),
.C(n_278),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_354),
.B(n_330),
.Y(n_363)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_313),
.A2(n_298),
.B1(n_305),
.B2(n_300),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_315),
.B(n_318),
.C(n_317),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_358),
.B(n_301),
.C(n_304),
.Y(n_378)
);

XOR2x2_ASAP7_75t_SL g359 ( 
.A(n_311),
.B(n_305),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_352),
.A2(n_317),
.B1(n_315),
.B2(n_323),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_361),
.A2(n_374),
.B1(n_356),
.B2(n_347),
.Y(n_387)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_378),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_300),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_367),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_368),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_359),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_370),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_344),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_345),
.Y(n_371)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_371),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_337),
.A2(n_323),
.B1(n_329),
.B2(n_331),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_322),
.Y(n_375)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_375),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_350),
.A2(n_304),
.B1(n_301),
.B2(n_292),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_376),
.A2(n_382),
.B1(n_383),
.B2(n_333),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_349),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_217),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_292),
.C(n_242),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_381),
.C(n_384),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_335),
.B(n_236),
.C(n_234),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_357),
.A2(n_297),
.B1(n_171),
.B2(n_234),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_348),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_236),
.C(n_221),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_364),
.A2(n_340),
.B(n_353),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_386),
.A2(n_398),
.B(n_402),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_388),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_362),
.A2(n_356),
.B1(n_347),
.B2(n_341),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_360),
.A2(n_338),
.B1(n_334),
.B2(n_154),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_365),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_375),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_362),
.Y(n_412)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_373),
.A2(n_338),
.B(n_153),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_372),
.B(n_221),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_403),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_217),
.C(n_164),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_384),
.C(n_381),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_373),
.A2(n_153),
.B(n_156),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_372),
.B(n_211),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_156),
.B(n_109),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_404),
.A2(n_371),
.B(n_376),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_401),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_407),
.B(n_411),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_408),
.B(n_417),
.Y(n_431)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_409),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_399),
.B(n_378),
.C(n_366),
.Y(n_411)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_412),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_366),
.C(n_380),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_423),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_416),
.A2(n_404),
.B1(n_405),
.B2(n_400),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_365),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_397),
.B(n_380),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_424),
.Y(n_438)
);

AOI22xp33_ASAP7_75t_SL g421 ( 
.A1(n_406),
.A2(n_374),
.B1(n_394),
.B2(n_371),
.Y(n_421)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_421),
.Y(n_440)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_386),
.B(n_377),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_385),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_R g427 ( 
.A(n_425),
.B(n_394),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_427),
.B(n_428),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_390),
.C(n_393),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_418),
.A2(n_398),
.B(n_387),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_430),
.A2(n_434),
.B(n_414),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_391),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_135),
.C(n_2),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_415),
.B(n_390),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_433),
.B(n_436),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_414),
.A2(n_402),
.B(n_392),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_420),
.B(n_403),
.C(n_408),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_437),
.A2(n_439),
.B1(n_409),
.B2(n_425),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_422),
.A2(n_385),
.B1(n_154),
.B2(n_118),
.Y(n_439)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_442),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_429),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_443),
.B(n_447),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_444),
.B(n_451),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_441),
.A2(n_416),
.B(n_424),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_445),
.B(n_449),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_435),
.A2(n_419),
.B(n_413),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_426),
.B(n_410),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_448),
.B(n_450),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_440),
.A2(n_410),
.B(n_131),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_430),
.A2(n_131),
.B(n_135),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_434),
.A2(n_1),
.B(n_2),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_453),
.B(n_455),
.Y(n_464)
);

NOR2x1_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_1),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_454),
.A2(n_437),
.B(n_439),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_2),
.C(n_3),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_460),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_431),
.C(n_436),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_465),
.Y(n_470)
);

INVx11_ASAP7_75t_L g463 ( 
.A(n_452),
.Y(n_463)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_463),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_431),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_432),
.C(n_438),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_461),
.Y(n_472)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_457),
.Y(n_469)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_469),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_456),
.A2(n_454),
.B(n_3),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_471),
.A2(n_464),
.B(n_458),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_472),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_459),
.B(n_2),
.Y(n_473)
);

O2A1O1Ixp33_ASAP7_75t_SL g477 ( 
.A1(n_473),
.A2(n_460),
.B(n_4),
.C(n_5),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_474),
.B(n_477),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_470),
.A2(n_462),
.B(n_463),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_476),
.A2(n_467),
.B(n_5),
.Y(n_481)
);

O2A1O1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_475),
.A2(n_468),
.B(n_467),
.C(n_466),
.Y(n_479)
);

OAI321xp33_ASAP7_75t_L g483 ( 
.A1(n_479),
.A2(n_481),
.A3(n_3),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_483)
);

AOI321xp33_ASAP7_75t_L g482 ( 
.A1(n_480),
.A2(n_478),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_482),
.B(n_483),
.C(n_6),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_484),
.A2(n_9),
.B(n_480),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_485),
.Y(n_486)
);


endmodule