module fake_netlist_1_2162_n_32 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_7), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
BUFx6f_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
AOI21xp5_ASAP7_75t_L g17 ( .A1(n_11), .A2(n_5), .B(n_6), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_13), .B(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_15), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_14), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_14), .Y(n_21) );
INVx3_ASAP7_75t_L g22 ( .A(n_19), .Y(n_22) );
BUFx10_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_22), .B(n_18), .Y(n_24) );
O2A1O1Ixp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_22), .B(n_17), .C(n_21), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_0), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_9), .B1(n_23), .B2(n_3), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_3), .Y(n_28) );
XOR2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_4), .Y(n_29) );
INVxp67_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
AOI21xp5_ASAP7_75t_L g31 ( .A1(n_30), .A2(n_25), .B(n_23), .Y(n_31) );
OR2x2_ASAP7_75t_L g32 ( .A(n_31), .B(n_29), .Y(n_32) );
endmodule