module fake_jpeg_5986_n_336 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_37),
.B(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_40),
.B1(n_34),
.B2(n_33),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_13),
.CON(n_40),
.SN(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_48),
.Y(n_80)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_51),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_53),
.Y(n_90)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g100 ( 
.A(n_55),
.Y(n_100)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g104 ( 
.A(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_22),
.B1(n_34),
.B2(n_20),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_62),
.B1(n_88),
.B2(n_96),
.Y(n_109)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_57),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_59),
.B(n_63),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_61),
.A2(n_98),
.B1(n_1),
.B2(n_2),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_36),
.B1(n_32),
.B2(n_23),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_65),
.Y(n_132)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_17),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_19),
.Y(n_106)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_81),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_48),
.A2(n_18),
.B1(n_35),
.B2(n_32),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_72),
.A2(n_75),
.B1(n_84),
.B2(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_52),
.A2(n_18),
.B1(n_35),
.B2(n_32),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_29),
.B1(n_28),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_92),
.B1(n_95),
.B2(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_89),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_39),
.A2(n_35),
.B1(n_18),
.B2(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_36),
.B1(n_20),
.B2(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_44),
.A2(n_23),
.B1(n_20),
.B2(n_16),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_43),
.B(n_28),
.Y(n_91)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_24),
.B1(n_15),
.B2(n_16),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_42),
.A2(n_16),
.B1(n_31),
.B2(n_30),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_33),
.B1(n_31),
.B2(n_27),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_45),
.A2(n_19),
.B1(n_17),
.B2(n_24),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_106),
.B(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_24),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_110),
.B(n_120),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_104),
.Y(n_111)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_113),
.A2(n_6),
.B(n_7),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_55),
.B1(n_49),
.B2(n_24),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_1),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_121),
.A2(n_123),
.B1(n_7),
.B2(n_8),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_71),
.A2(n_55),
.B1(n_49),
.B2(n_6),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_95),
.A2(n_77),
.B1(n_88),
.B2(n_76),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_128),
.B1(n_87),
.B2(n_85),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_49),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_3),
.Y(n_131)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_136),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_69),
.B(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_106),
.Y(n_144)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_3),
.Y(n_137)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_8),
.B(n_9),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_3),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_138),
.A2(n_134),
.B(n_110),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_59),
.B1(n_105),
.B2(n_76),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_142),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_103),
.B1(n_89),
.B2(n_93),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_143),
.A2(n_158),
.B1(n_169),
.B2(n_107),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_144),
.B(n_133),
.Y(n_202)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_146),
.B(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_90),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_161),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_102),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_152),
.Y(n_203)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_79),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_166),
.B1(n_170),
.B2(n_135),
.Y(n_206)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_79),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_164),
.C(n_119),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_155),
.A2(n_112),
.B(n_116),
.Y(n_205)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_156),
.B(n_159),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_68),
.B1(n_73),
.B2(n_64),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_124),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_160),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_120),
.B(n_82),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_80),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_165),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_125),
.B(n_78),
.C(n_60),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_5),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_119),
.A2(n_94),
.B1(n_67),
.B2(n_60),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_127),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_111),
.B(n_67),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_173),
.B(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_122),
.B(n_8),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_175),
.B(n_176),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_193),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_181),
.A2(n_198),
.B1(n_206),
.B2(n_151),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_149),
.A2(n_131),
.B(n_137),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_182),
.A2(n_188),
.B(n_162),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_140),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_184),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_186),
.A2(n_194),
.B1(n_195),
.B2(n_204),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_163),
.A2(n_139),
.B1(n_118),
.B2(n_112),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_207),
.B1(n_213),
.B2(n_214),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_126),
.Y(n_192)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_192),
.Y(n_222)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_126),
.Y(n_196)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_164),
.B(n_127),
.C(n_129),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_211),
.C(n_140),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_154),
.A2(n_135),
.B1(n_108),
.B2(n_118),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_140),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_159),
.B(n_156),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_152),
.A2(n_108),
.B1(n_136),
.B2(n_107),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_174),
.B(n_116),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_209),
.Y(n_221)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_153),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_141),
.B(n_116),
.C(n_107),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_150),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_141),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_237),
.Y(n_244)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_241),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_218),
.A2(n_234),
.B(n_238),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_233),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_151),
.B1(n_169),
.B2(n_146),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_181),
.A2(n_206),
.B1(n_195),
.B2(n_183),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_147),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_232),
.C(n_236),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_180),
.B(n_172),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_145),
.B1(n_162),
.B2(n_160),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_145),
.B(n_10),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_235),
.B(n_242),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_196),
.A2(n_9),
.B(n_11),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_178),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_222),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_204),
.B(n_160),
.C(n_9),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_199),
.C(n_177),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_187),
.A2(n_12),
.B1(n_194),
.B2(n_203),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_180),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_203),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_250),
.C(n_255),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_248),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_239),
.B(n_191),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_261),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_211),
.Y(n_250)
);

OAI32xp33_ASAP7_75t_L g251 ( 
.A1(n_229),
.A2(n_190),
.A3(n_192),
.B1(n_188),
.B2(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_189),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_222),
.B(n_193),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_256),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_218),
.B(n_182),
.C(n_188),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_229),
.B(n_208),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_185),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_227),
.B(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_259),
.B(n_265),
.C(n_245),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_235),
.B(n_191),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_262),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_263),
.A2(n_233),
.B(n_242),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_217),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_177),
.C(n_200),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_228),
.B1(n_220),
.B2(n_221),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_274),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_228),
.B1(n_220),
.B2(n_221),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_241),
.B1(n_226),
.B2(n_234),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_280),
.B1(n_256),
.B2(n_260),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_284),
.C(n_277),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_251),
.A2(n_243),
.B1(n_240),
.B2(n_231),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_283),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_247),
.A2(n_232),
.B1(n_238),
.B2(n_223),
.Y(n_281)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_255),
.A2(n_12),
.B1(n_200),
.B2(n_267),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_12),
.C(n_265),
.Y(n_284)
);

FAx1_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_244),
.CI(n_267),
.CON(n_287),
.SN(n_287)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_287),
.A2(n_289),
.B(n_283),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_244),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_291),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_250),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_294),
.B(n_279),
.Y(n_301)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_295),
.B(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_246),
.Y(n_297)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_297),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_284),
.C(n_282),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_299),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_259),
.C(n_254),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_271),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_268),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_305),
.C(n_311),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_275),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_307),
.B(n_286),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_263),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_304),
.B(n_309),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_280),
.B1(n_272),
.B2(n_271),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_268),
.B(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_300),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_303),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_294),
.C(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_318),
.C(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_320),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_288),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_291),
.C(n_299),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_281),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_315),
.B(n_269),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_326),
.Y(n_328)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_302),
.B(n_312),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_310),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_324),
.B(n_311),
.C(n_290),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_330),
.C(n_269),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_329),
.A2(n_325),
.A3(n_323),
.B1(n_328),
.B2(n_313),
.C1(n_258),
.C2(n_287),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_276),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_331),
.B(n_332),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_307),
.C(n_329),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_285),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);


endmodule