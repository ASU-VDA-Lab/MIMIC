module fake_jpeg_20679_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

BUFx2_ASAP7_75t_SL g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_7),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_21),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_21),
.B1(n_16),
.B2(n_24),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_49),
.B1(n_26),
.B2(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_40),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_16),
.B1(n_24),
.B2(n_25),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_50),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_56),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_36),
.B1(n_24),
.B2(n_37),
.Y(n_55)
);

AO21x2_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_58),
.B(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_28),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_34),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_57),
.A2(n_44),
.B(n_51),
.Y(n_77)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_49),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_66),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_18),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_70),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_43),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_2),
.C(n_3),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_15),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_0),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_5),
.C(n_8),
.Y(n_87)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_81),
.B(n_82),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_44),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_59),
.C(n_65),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_57),
.A2(n_3),
.B(n_5),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_57),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_55),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_5),
.B(n_7),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_91),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_97),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_60),
.B1(n_55),
.B2(n_58),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_96),
.B(n_98),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_60),
.B1(n_73),
.B2(n_66),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_92),
.Y(n_107)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_85),
.B(n_77),
.C(n_78),
.D(n_80),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_95),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_88),
.C(n_79),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_95),
.C(n_86),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_99),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_109),
.C(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_104),
.C(n_100),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_113),
.B(n_114),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_103),
.A2(n_102),
.B1(n_78),
.B2(n_89),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_103),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_106),
.A3(n_78),
.B1(n_105),
.B2(n_89),
.C1(n_72),
.C2(n_11),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_118),
.B(n_115),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_123),
.Y(n_124)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_106),
.B(n_10),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_9),
.C(n_118),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_124),
.A2(n_121),
.B1(n_59),
.B2(n_10),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_126),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_127),
.Y(n_129)
);


endmodule