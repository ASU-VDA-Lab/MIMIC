module fake_jpeg_10707_n_563 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_563);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_563;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_7),
.B(n_3),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_1),
.Y(n_55)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_56),
.Y(n_60)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_61),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_63),
.B(n_98),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_42),
.B(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_65),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_66),
.B(n_69),
.Y(n_131)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_67),
.Y(n_170)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_70),
.Y(n_154)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_72),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_0),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_73),
.B(n_108),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_74),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_75),
.B(n_78),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_79),
.Y(n_173)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

INVx6_ASAP7_75t_SL g82 ( 
.A(n_38),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_88),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_30),
.Y(n_89)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_53),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_90),
.B(n_92),
.Y(n_161)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_53),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_40),
.Y(n_93)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_95),
.B(n_112),
.Y(n_162)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_37),
.B(n_15),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_99),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_102),
.Y(n_209)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_103),
.Y(n_203)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_104),
.Y(n_187)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_106),
.Y(n_201)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_22),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_20),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_114),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_20),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_13),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_115),
.B(n_116),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_13),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_118),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_34),
.B(n_13),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_23),
.Y(n_120)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_120),
.Y(n_207)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_19),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_121),
.B(n_123),
.Y(n_210)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_122),
.B(n_126),
.Y(n_168)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_25),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_23),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_124),
.B(n_125),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_31),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_41),
.B1(n_36),
.B2(n_32),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_130),
.A2(n_151),
.B1(n_155),
.B2(n_159),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_32),
.B1(n_41),
.B2(n_36),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_136),
.A2(n_138),
.B1(n_158),
.B2(n_64),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_73),
.A2(n_41),
.B1(n_32),
.B2(n_36),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_73),
.A2(n_51),
.B1(n_58),
.B2(n_35),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_144),
.A2(n_148),
.B(n_152),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_93),
.A2(n_43),
.B1(n_25),
.B2(n_49),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_79),
.A2(n_51),
.B1(n_32),
.B2(n_55),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_25),
.B1(n_49),
.B2(n_43),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_96),
.A2(n_51),
.B1(n_43),
.B2(n_49),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_82),
.B(n_29),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_157),
.B(n_74),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_24),
.B1(n_50),
.B2(n_48),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_97),
.A2(n_29),
.B1(n_50),
.B2(n_48),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_83),
.B(n_35),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_160),
.B(n_169),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_59),
.B(n_55),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_86),
.B(n_29),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_174),
.B(n_177),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_52),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_77),
.A2(n_85),
.B1(n_91),
.B2(n_121),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_178),
.A2(n_180),
.B1(n_181),
.B2(n_199),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_99),
.A2(n_47),
.B1(n_44),
.B2(n_28),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_124),
.A2(n_52),
.B1(n_34),
.B2(n_44),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_87),
.B(n_12),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_186),
.B(n_188),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_87),
.B(n_47),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_61),
.B(n_28),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_193),
.B(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_67),
.B(n_26),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_106),
.B(n_26),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_197),
.B(n_198),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_84),
.B(n_24),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_62),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_107),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_123),
.B1(n_88),
.B2(n_117),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_110),
.B(n_1),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_206),
.B(n_208),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_72),
.B(n_4),
.Y(n_208)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_5),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_212),
.B(n_223),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_103),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_213),
.B(n_233),
.Y(n_288)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_168),
.Y(n_214)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_214),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_215),
.Y(n_295)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_219),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_220),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_221),
.A2(n_248),
.B1(n_239),
.B2(n_190),
.Y(n_312)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_129),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_222),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_5),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_136),
.A2(n_81),
.B1(n_111),
.B2(n_109),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_224),
.Y(n_308)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_185),
.Y(n_225)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_225),
.Y(n_322)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_157),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_239),
.Y(n_283)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_228),
.Y(n_331)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_229),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_144),
.B(n_6),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_231),
.B(n_234),
.Y(n_301)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_187),
.Y(n_232)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_232),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_131),
.B(n_125),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_127),
.B(n_8),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_8),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_235),
.B(n_240),
.Y(n_311)
);

INVx4_ASAP7_75t_SL g236 ( 
.A(n_176),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_241),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_162),
.B(n_108),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_238),
.B(n_258),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_157),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_156),
.B(n_8),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_141),
.Y(n_242)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g244 ( 
.A(n_128),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_244),
.B(n_263),
.Y(n_329)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_167),
.Y(n_247)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_167),
.A2(n_70),
.B1(n_101),
.B2(n_100),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_249),
.A2(n_140),
.B1(n_171),
.B2(n_166),
.Y(n_324)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_250),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_251),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_133),
.B(n_139),
.C(n_138),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_252),
.B(n_257),
.C(n_272),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_170),
.Y(n_253)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_253),
.Y(n_325)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_143),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_260),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_161),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_255),
.B(n_256),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_180),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g257 ( 
.A(n_147),
.B(n_102),
.C(n_60),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_209),
.B(n_8),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_135),
.B(n_10),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_259),
.B(n_281),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_158),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_154),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_264),
.Y(n_300)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_145),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_265),
.B(n_274),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_150),
.B(n_10),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_266),
.B(n_267),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_150),
.B(n_153),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_271),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_189),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_270),
.Y(n_323)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_192),
.Y(n_271)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_201),
.B(n_89),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_210),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_273),
.B(n_275),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_191),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_202),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_134),
.B(n_11),
.Y(n_277)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_277),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_159),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_280),
.Y(n_290)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_134),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_170),
.B(n_11),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_227),
.A2(n_178),
.B1(n_210),
.B2(n_152),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_285),
.A2(n_269),
.B1(n_241),
.B2(n_243),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_230),
.A2(n_148),
.B(n_205),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_292),
.A2(n_305),
.B(n_316),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_201),
.C(n_196),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_296),
.B(n_307),
.C(n_313),
.Y(n_339)
);

OA21x2_ASAP7_75t_L g297 ( 
.A1(n_231),
.A2(n_155),
.B(n_203),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_297),
.A2(n_274),
.B(n_265),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_212),
.B(n_149),
.CI(n_203),
.CON(n_304),
.SN(n_304)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_304),
.B(n_244),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_190),
.B(n_149),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_191),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_312),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g313 ( 
.A(n_218),
.B(n_234),
.C(n_223),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_241),
.A2(n_60),
.B(n_207),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_259),
.B(n_171),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_336),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_324),
.A2(n_328),
.B1(n_154),
.B2(n_183),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_237),
.B(n_102),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_236),
.C(n_265),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_249),
.A2(n_140),
.B1(n_166),
.B2(n_164),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_279),
.B(n_164),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_318),
.B(n_235),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_337),
.B(n_338),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_291),
.B(n_261),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_252),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_355),
.C(n_364),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_342),
.B(n_344),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_302),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_343),
.B(n_348),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_308),
.A2(n_272),
.B1(n_216),
.B2(n_173),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_345),
.A2(n_347),
.B1(n_369),
.B2(n_375),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_297),
.A2(n_272),
.B1(n_173),
.B2(n_274),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g348 ( 
.A(n_298),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_240),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_349),
.B(n_351),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_286),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_225),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_352),
.A2(n_373),
.B1(n_319),
.B2(n_289),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_300),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_362),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_336),
.B(n_228),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_360),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_313),
.B(n_232),
.Y(n_355)
);

AOI21xp33_ASAP7_75t_L g399 ( 
.A1(n_356),
.A2(n_372),
.B(n_377),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_329),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_357),
.B(n_359),
.Y(n_408)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_321),
.Y(n_358)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_358),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_247),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_315),
.B(n_263),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_290),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_363),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_280),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_315),
.B(n_271),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_283),
.C(n_296),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_311),
.B(n_211),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_371),
.Y(n_397)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_282),
.Y(n_367)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_295),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_297),
.A2(n_146),
.B1(n_254),
.B2(n_175),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_222),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_314),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_317),
.B(n_219),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_292),
.A2(n_183),
.B1(n_175),
.B2(n_146),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_305),
.A2(n_290),
.B(n_287),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_374),
.A2(n_376),
.B(n_316),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_301),
.A2(n_172),
.B1(n_179),
.B2(n_262),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_298),
.A2(n_246),
.B(n_245),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_325),
.A2(n_250),
.B1(n_253),
.B2(n_220),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_SL g378 ( 
.A1(n_325),
.A2(n_172),
.B1(n_179),
.B2(n_215),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_SL g392 ( 
.A(n_378),
.B(n_329),
.C(n_319),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_342),
.A2(n_324),
.B1(n_328),
.B2(n_301),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_379),
.B(n_396),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_380),
.B(n_341),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g381 ( 
.A(n_339),
.B(n_311),
.C(n_286),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_401),
.C(n_364),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_339),
.B(n_327),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_391),
.B(n_370),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_392),
.A2(n_366),
.B(n_344),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_393),
.Y(n_441)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_394),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_346),
.A2(n_320),
.B1(n_304),
.B2(n_303),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_346),
.A2(n_304),
.B1(n_289),
.B2(n_295),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_398),
.A2(n_334),
.B1(n_309),
.B2(n_368),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_373),
.A2(n_352),
.B1(n_358),
.B2(n_340),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_400),
.A2(n_404),
.B1(n_347),
.B2(n_369),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_351),
.B(n_330),
.C(n_329),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_359),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_411),
.Y(n_422)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_367),
.Y(n_403)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_403),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_340),
.A2(n_282),
.B1(n_284),
.B2(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_284),
.Y(n_405)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_405),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_337),
.B(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_360),
.B(n_294),
.Y(n_409)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_409),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_375),
.Y(n_412)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_412),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_414),
.B(n_421),
.C(n_430),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_417),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_416),
.Y(n_448)
);

XOR2x2_ASAP7_75t_SL g417 ( 
.A(n_396),
.B(n_356),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_410),
.A2(n_366),
.B(n_374),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_418),
.A2(n_393),
.B(n_408),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_419),
.A2(n_423),
.B1(n_443),
.B2(n_379),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_420),
.A2(n_434),
.B(n_413),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_385),
.B(n_349),
.C(n_355),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_410),
.A2(n_345),
.B1(n_363),
.B2(n_350),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_383),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_397),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_428),
.B(n_431),
.Y(n_467)
);

OAI211xp5_ASAP7_75t_L g429 ( 
.A1(n_387),
.A2(n_371),
.B(n_353),
.C(n_357),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_429),
.B(n_437),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_385),
.B(n_370),
.C(n_376),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_397),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_404),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_433),
.B(n_440),
.Y(n_469)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_395),
.B(n_334),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_411),
.B(n_343),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_438),
.A2(n_412),
.B1(n_394),
.B2(n_413),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_388),
.B(n_310),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g447 ( 
.A(n_439),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_386),
.B(n_310),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_400),
.A2(n_368),
.B1(n_242),
.B2(n_251),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_444),
.A2(n_432),
.B1(n_416),
.B2(n_443),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_441),
.A2(n_398),
.B1(n_399),
.B2(n_407),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_446),
.A2(n_463),
.B1(n_465),
.B2(n_438),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_414),
.B(n_382),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_453),
.C(n_456),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_425),
.A2(n_382),
.B1(n_383),
.B2(n_395),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_451),
.A2(n_464),
.B1(n_427),
.B2(n_442),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_460),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_421),
.B(n_380),
.C(n_381),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_422),
.Y(n_455)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_455),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_415),
.B(n_391),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_428),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_457),
.B(n_461),
.Y(n_475)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_401),
.C(n_406),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_462),
.C(n_468),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_420),
.A2(n_384),
.B(n_392),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_424),
.B(n_386),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_425),
.A2(n_405),
.B1(n_409),
.B2(n_403),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_419),
.A2(n_390),
.B1(n_389),
.B2(n_334),
.Y(n_465)
);

A2O1A1O1Ixp25_ASAP7_75t_L g466 ( 
.A1(n_418),
.A2(n_417),
.B(n_435),
.C(n_436),
.D(n_427),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_466),
.B(n_434),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_390),
.C(n_299),
.Y(n_468)
);

OA22x2_ASAP7_75t_L g471 ( 
.A1(n_463),
.A2(n_431),
.B1(n_433),
.B2(n_416),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_471),
.B(n_472),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_477),
.A2(n_479),
.B1(n_491),
.B2(n_468),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_442),
.Y(n_478)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_478),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_447),
.A2(n_435),
.B1(n_436),
.B2(n_432),
.Y(n_482)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_482),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_426),
.C(n_294),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_483),
.B(n_490),
.C(n_449),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g486 ( 
.A(n_470),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_488),
.Y(n_495)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_464),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_487),
.B(n_489),
.Y(n_496)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_469),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_451),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_445),
.B(n_299),
.C(n_306),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_434),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_491),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_492),
.A2(n_452),
.B(n_450),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_453),
.B(n_306),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_460),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_481),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_498),
.A2(n_484),
.B1(n_488),
.B2(n_471),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_483),
.B(n_456),
.C(n_459),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_503),
.Y(n_522)
);

INVx13_ASAP7_75t_L g501 ( 
.A(n_480),
.Y(n_501)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_501),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_444),
.Y(n_502)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_502),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_504),
.A2(n_484),
.B(n_475),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_454),
.C(n_462),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_505),
.B(n_507),
.C(n_508),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_474),
.B(n_454),
.C(n_461),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_474),
.B(n_446),
.C(n_466),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_481),
.B(n_293),
.C(n_333),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_497),
.C(n_499),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_509),
.B(n_479),
.Y(n_514)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_514),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_506),
.B(n_495),
.Y(n_516)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_516),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_517),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_519),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_495),
.B(n_473),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_520),
.A2(n_502),
.B1(n_504),
.B2(n_494),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_510),
.B(n_471),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_523),
.Y(n_536)
);

FAx1_ASAP7_75t_SL g524 ( 
.A(n_508),
.B(n_485),
.CI(n_471),
.CON(n_524),
.SN(n_524)
);

BUFx24_ASAP7_75t_SL g534 ( 
.A(n_524),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_496),
.B(n_477),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g531 ( 
.A1(n_525),
.A2(n_515),
.B1(n_514),
.B2(n_516),
.Y(n_531)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_528),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_520),
.B(n_485),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_523),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_531),
.A2(n_533),
.B1(n_526),
.B2(n_535),
.Y(n_543)
);

OAI21xp33_ASAP7_75t_L g532 ( 
.A1(n_521),
.A2(n_494),
.B(n_503),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_532),
.B(n_512),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_525),
.A2(n_494),
.B1(n_500),
.B2(n_507),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_522),
.A2(n_511),
.B1(n_505),
.B2(n_501),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_537),
.B(n_518),
.Y(n_545)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_534),
.B(n_524),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_538),
.B(n_541),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_SL g539 ( 
.A1(n_529),
.A2(n_517),
.B(n_513),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_539),
.A2(n_532),
.B(n_309),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_540),
.B(n_546),
.Y(n_549)
);

FAx1_ASAP7_75t_SL g541 ( 
.A(n_529),
.B(n_513),
.CI(n_524),
.CON(n_541),
.SN(n_541)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_543),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_545),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_322),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_536),
.C(n_530),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_548),
.B(n_550),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_293),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_553),
.B(n_333),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_554),
.B(n_557),
.Y(n_559)
);

OAI31xp33_ASAP7_75t_SL g555 ( 
.A1(n_551),
.A2(n_538),
.A3(n_541),
.B(n_331),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g558 ( 
.A1(n_555),
.A2(n_552),
.B(n_553),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_549),
.B(n_538),
.Y(n_557)
);

BUFx24_ASAP7_75t_SL g560 ( 
.A(n_558),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_556),
.B1(n_547),
.B2(n_559),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_538),
.B(n_322),
.Y(n_562)
);

AO21x1_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_331),
.B(n_11),
.Y(n_563)
);


endmodule