module fake_jpeg_23315_n_32 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_32);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_19),
.Y(n_20)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_17),
.B(n_8),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_21),
.A2(n_22),
.B(n_1),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_2),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_26),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_10),
.B1(n_3),
.B2(n_4),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_22),
.B1(n_2),
.B2(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_25),
.Y(n_30)
);

A2O1A1O1Ixp25_ASAP7_75t_L g31 ( 
.A1(n_30),
.A2(n_29),
.B(n_27),
.C(n_12),
.D(n_13),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_5),
.B(n_11),
.C(n_15),
.Y(n_32)
);


endmodule