module fake_netlist_1_4488_n_566 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_566);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_566;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_61), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_46), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_33), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_28), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_24), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_9), .Y(n_86) );
CKINVDCx16_ASAP7_75t_R g87 ( .A(n_22), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_57), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_29), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_75), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_39), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_40), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_48), .Y(n_93) );
CKINVDCx16_ASAP7_75t_R g94 ( .A(n_47), .Y(n_94) );
BUFx2_ASAP7_75t_L g95 ( .A(n_41), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_36), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_8), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_3), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_73), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_21), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_58), .Y(n_101) );
INVx2_ASAP7_75t_SL g102 ( .A(n_69), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_64), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
INVxp33_ASAP7_75t_L g105 ( .A(n_66), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_63), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_30), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_54), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_19), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_18), .Y(n_113) );
CKINVDCx16_ASAP7_75t_R g114 ( .A(n_79), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_4), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_42), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_44), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_81), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_95), .B(n_0), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_90), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_95), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_113), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_88), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_102), .B(n_0), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_104), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
OA21x2_ASAP7_75t_L g133 ( .A1(n_91), .A2(n_32), .B(n_77), .Y(n_133) );
NAND2xp5_ASAP7_75t_SL g134 ( .A(n_102), .B(n_84), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_87), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_91), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_94), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_92), .Y(n_140) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_86), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_127), .B(n_114), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_125), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_127), .B(n_80), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_131), .B(n_105), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_119), .B(n_80), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_118), .Y(n_148) );
OR2x2_ASAP7_75t_L g149 ( .A(n_131), .B(n_86), .Y(n_149) );
INVx4_ASAP7_75t_L g150 ( .A(n_118), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_125), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_119), .B(n_107), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_122), .Y(n_153) );
INVxp33_ASAP7_75t_L g154 ( .A(n_134), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g156 ( .A(n_120), .B(n_111), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_120), .B(n_106), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g159 ( .A1(n_121), .A2(n_129), .B1(n_140), .B2(n_139), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
BUFx4f_ASAP7_75t_L g161 ( .A(n_121), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
INVx4_ASAP7_75t_L g163 ( .A(n_118), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_124), .B(n_107), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_124), .B(n_98), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_129), .B(n_132), .Y(n_166) );
OAI22xp33_ASAP7_75t_L g167 ( .A1(n_141), .A2(n_115), .B1(n_97), .B2(n_108), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_132), .B(n_115), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_161), .B(n_83), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_149), .B(n_137), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_161), .B(n_83), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_161), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_166), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_166), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_166), .Y(n_175) );
NAND2xp33_ASAP7_75t_SL g176 ( .A(n_153), .B(n_123), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_166), .A2(n_140), .B1(n_139), .B2(n_137), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_153), .B(n_130), .Y(n_178) );
AND2x4_ASAP7_75t_SL g179 ( .A(n_145), .B(n_128), .Y(n_179) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_168), .A2(n_141), .B1(n_125), .B2(n_111), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_161), .B(n_93), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_159), .B(n_93), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_145), .A2(n_101), .B1(n_112), .B2(n_116), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g186 ( .A(n_168), .B(n_133), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_157), .B(n_101), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_143), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_158), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_151), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_168), .Y(n_196) );
AND2x2_ASAP7_75t_SL g197 ( .A(n_168), .B(n_133), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_149), .B(n_126), .Y(n_199) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_146), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_147), .B(n_126), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_165), .Y(n_202) );
BUFx4f_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
OR2x6_ASAP7_75t_L g204 ( .A(n_187), .B(n_162), .Y(n_204) );
CKINVDCx12_ASAP7_75t_R g205 ( .A(n_187), .Y(n_205) );
CKINVDCx10_ASAP7_75t_R g206 ( .A(n_179), .Y(n_206) );
INVx3_ASAP7_75t_SL g207 ( .A(n_179), .Y(n_207) );
NAND2x1_ASAP7_75t_L g208 ( .A(n_174), .B(n_150), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_170), .B(n_144), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_180), .B(n_142), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_173), .Y(n_211) );
AND2x2_ASAP7_75t_L g212 ( .A(n_170), .B(n_162), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_173), .Y(n_213) );
AOI221x1_ASAP7_75t_L g214 ( .A1(n_185), .A2(n_146), .B1(n_118), .B2(n_136), .C(n_117), .Y(n_214) );
OR2x6_ASAP7_75t_L g215 ( .A(n_196), .B(n_152), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_196), .Y(n_216) );
BUFx12f_ASAP7_75t_L g217 ( .A(n_199), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_203), .Y(n_218) );
BUFx4f_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_174), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_178), .B(n_156), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_197), .A2(n_185), .B(n_200), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_197), .A2(n_146), .B(n_164), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_203), .B(n_126), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_177), .B(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_175), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_197), .A2(n_146), .B(n_164), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_185), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_177), .B(n_146), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_190), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_202), .B(n_154), .Y(n_235) );
CKINVDCx6p67_ASAP7_75t_R g236 ( .A(n_202), .Y(n_236) );
AOI22xp33_ASAP7_75t_SL g237 ( .A1(n_203), .A2(n_167), .B1(n_126), .B2(n_133), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_192), .A2(n_112), .B(n_116), .C(n_117), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_209), .B(n_175), .Y(n_239) );
OAI21x1_ASAP7_75t_SL g240 ( .A1(n_233), .A2(n_194), .B(n_193), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_223), .A2(n_186), .B(n_193), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_214), .A2(n_186), .B(n_192), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_209), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_219), .A2(n_176), .B1(n_181), .B2(n_199), .Y(n_244) );
INVx5_ASAP7_75t_L g245 ( .A(n_224), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_225), .A2(n_186), .B(n_194), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_219), .B(n_199), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_226), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_204), .B(n_184), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_204), .Y(n_250) );
NOR2xp33_ASAP7_75t_SL g251 ( .A(n_207), .B(n_172), .Y(n_251) );
OAI21x1_ASAP7_75t_L g252 ( .A1(n_230), .A2(n_198), .B(n_148), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_209), .B(n_172), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_222), .A2(n_181), .B(n_189), .C(n_201), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_232), .A2(n_198), .B(n_160), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_204), .B(n_183), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_212), .A2(n_182), .B1(n_169), .B2(n_171), .C(n_100), .Y(n_257) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_232), .A2(n_148), .B(n_160), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g259 ( .A1(n_210), .A2(n_82), .B1(n_99), .B2(n_103), .C(n_109), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_233), .A2(n_160), .B(n_195), .Y(n_260) );
OR2x2_ASAP7_75t_L g261 ( .A(n_207), .B(n_188), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_235), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_206), .Y(n_264) );
OA21x2_ASAP7_75t_L g265 ( .A1(n_238), .A2(n_110), .B(n_195), .Y(n_265) );
OAI21x1_ASAP7_75t_SL g266 ( .A1(n_234), .A2(n_191), .B(n_188), .Y(n_266) );
AO21x2_ASAP7_75t_L g267 ( .A1(n_238), .A2(n_191), .B(n_200), .Y(n_267) );
AOI221xp5_ASAP7_75t_L g268 ( .A1(n_259), .A2(n_227), .B1(n_211), .B2(n_213), .C(n_229), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_240), .A2(n_231), .B(n_224), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_240), .A2(n_231), .B(n_224), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_249), .A2(n_217), .B1(n_215), .B2(n_236), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_262), .B(n_215), .Y(n_272) );
AOI22xp33_ASAP7_75t_SL g273 ( .A1(n_251), .A2(n_217), .B1(n_205), .B2(n_218), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_244), .A2(n_215), .B1(n_236), .B2(n_216), .Y(n_274) );
OAI332xp33_ASAP7_75t_L g275 ( .A1(n_263), .A2(n_264), .A3(n_243), .B1(n_256), .B2(n_261), .B3(n_262), .C1(n_205), .C2(n_228), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_252), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_267), .A2(n_237), .B(n_216), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_254), .A2(n_231), .B(n_224), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_226), .B(n_208), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_252), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_246), .A2(n_150), .B(n_163), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_265), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_250), .B(n_221), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_248), .B(n_231), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_246), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_260), .Y(n_288) );
AOI21x1_ASAP7_75t_L g289 ( .A1(n_255), .A2(n_200), .B(n_185), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_253), .B(n_221), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_253), .A2(n_221), .B1(n_220), .B2(n_200), .Y(n_291) );
BUFx2_ASAP7_75t_L g292 ( .A(n_287), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_276), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_277), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_272), .B(n_267), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_272), .B(n_267), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_277), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
NOR2x1_ASAP7_75t_SL g299 ( .A(n_286), .B(n_245), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_287), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_282), .Y(n_301) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_290), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_281), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_290), .B(n_247), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_275), .B(n_239), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_275), .B(n_239), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_284), .B(n_248), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_288), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_286), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_290), .B(n_247), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
BUFx3_ASAP7_75t_L g316 ( .A(n_312), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_298), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_294), .B(n_278), .Y(n_318) );
AND2x2_ASAP7_75t_L g319 ( .A(n_296), .B(n_278), .Y(n_319) );
NAND3xp33_ASAP7_75t_SL g320 ( .A(n_313), .B(n_273), .C(n_271), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_292), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_294), .B(n_278), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_297), .Y(n_325) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_300), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_296), .B(n_288), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_295), .B(n_286), .Y(n_329) );
AOI33xp33_ASAP7_75t_L g330 ( .A1(n_304), .A2(n_274), .A3(n_239), .B1(n_96), .B2(n_268), .B3(n_253), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_295), .B(n_286), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_306), .A2(n_290), .B1(n_286), .B2(n_291), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_309), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_297), .B(n_283), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_308), .A2(n_314), .B1(n_304), .B2(n_302), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_301), .B(n_283), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_301), .B(n_307), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_307), .B(n_241), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_311), .B(n_241), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_314), .B(n_261), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_311), .B(n_258), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
NOR3xp33_ASAP7_75t_L g344 ( .A(n_312), .B(n_257), .C(n_163), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_312), .B(n_289), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_317), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_326), .B(n_310), .Y(n_347) );
INVxp67_ASAP7_75t_L g348 ( .A(n_334), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_338), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_338), .B(n_310), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_329), .B(n_305), .Y(n_351) );
OA21x2_ASAP7_75t_L g352 ( .A1(n_318), .A2(n_305), .B(n_289), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_328), .B(n_303), .Y(n_353) );
INVx3_ASAP7_75t_L g354 ( .A(n_345), .Y(n_354) );
OAI33xp33_ASAP7_75t_L g355 ( .A1(n_325), .A2(n_2), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_328), .B(n_303), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_336), .B(n_299), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_319), .B(n_293), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_319), .B(n_293), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_322), .B(n_245), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_322), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_335), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_327), .B(n_245), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_320), .B(n_6), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_337), .B(n_299), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_345), .B(n_280), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_337), .B(n_258), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
AOI21xp5_ASAP7_75t_SL g373 ( .A1(n_321), .A2(n_270), .B(n_269), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_323), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_323), .Y(n_376) );
INVx6_ASAP7_75t_L g377 ( .A(n_316), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_333), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_329), .B(n_136), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_336), .B(n_7), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_344), .A2(n_332), .B1(n_331), .B2(n_316), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_333), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_331), .B(n_136), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_315), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_339), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_339), .B(n_136), .Y(n_387) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_343), .B(n_279), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_340), .B(n_315), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_136), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g391 ( .A(n_366), .B(n_330), .C(n_318), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_349), .B(n_340), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_348), .B(n_332), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_372), .B(n_343), .Y(n_394) );
INVx1_ASAP7_75t_SL g395 ( .A(n_377), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_364), .B(n_324), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_346), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_357), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_361), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_364), .B(n_324), .Y(n_403) );
NOR2x1_ASAP7_75t_L g404 ( .A(n_365), .B(n_316), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_389), .B(n_345), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_386), .B(n_315), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_386), .B(n_315), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_347), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_389), .B(n_342), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_359), .B(n_342), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_369), .B(n_341), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_359), .B(n_136), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_360), .B(n_8), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_360), .B(n_9), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_367), .B(n_10), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_353), .B(n_242), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_367), .B(n_10), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_351), .B(n_11), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_353), .B(n_242), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_380), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_356), .B(n_280), .Y(n_423) );
INVx4_ASAP7_75t_L g424 ( .A(n_362), .Y(n_424) );
NAND2x1_ASAP7_75t_L g425 ( .A(n_377), .B(n_266), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_356), .B(n_12), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_387), .B(n_12), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_380), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_354), .Y(n_429) );
NOR2x1_ASAP7_75t_SL g430 ( .A(n_358), .B(n_245), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_384), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_354), .B(n_13), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_351), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_354), .B(n_13), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_374), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_374), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_375), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_387), .B(n_14), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_381), .B(n_14), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_363), .B(n_15), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_371), .B(n_15), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_382), .B(n_16), .Y(n_443) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_390), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_409), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_441), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_417), .B(n_370), .Y(n_447) );
AOI21xp33_ASAP7_75t_L g448 ( .A1(n_443), .A2(n_390), .B(n_371), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_398), .Y(n_449) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_391), .A2(n_362), .B(n_373), .Y(n_450) );
OAI31xp33_ASAP7_75t_L g451 ( .A1(n_416), .A2(n_362), .A3(n_369), .B(n_371), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_430), .A2(n_373), .B(n_355), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_434), .B(n_376), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_397), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_413), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_424), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_R g457 ( .A1(n_419), .A2(n_385), .B(n_379), .C(n_368), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_393), .B(n_370), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_394), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g461 ( .A1(n_393), .A2(n_377), .B1(n_388), .B2(n_383), .C(n_375), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_405), .B(n_369), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_424), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_436), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g465 ( .A1(n_440), .A2(n_383), .B(n_378), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_437), .Y(n_466) );
BUFx3_ASAP7_75t_L g467 ( .A(n_424), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_397), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_441), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_413), .B(n_378), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_438), .Y(n_471) );
AOI22x1_ASAP7_75t_SL g472 ( .A1(n_395), .A2(n_377), .B1(n_376), .B2(n_379), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_412), .A2(n_368), .B1(n_385), .B2(n_352), .Y(n_473) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_440), .A2(n_352), .B(n_16), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_410), .B(n_352), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_408), .B(n_352), .Y(n_476) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_414), .B(n_163), .C(n_150), .D(n_220), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_406), .Y(n_478) );
NAND2xp33_ASAP7_75t_L g479 ( .A(n_404), .B(n_245), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_407), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_410), .B(n_163), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_426), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_425), .A2(n_266), .B(n_260), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_392), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_411), .B(n_150), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_429), .B(n_200), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_396), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_403), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_411), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
OAI221xp5_ASAP7_75t_SL g491 ( .A1(n_451), .A2(n_420), .B1(n_415), .B2(n_426), .C(n_439), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_478), .Y(n_492) );
NOR3xp33_ASAP7_75t_L g493 ( .A(n_450), .B(n_427), .C(n_442), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_446), .A2(n_412), .B1(n_405), .B2(n_435), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_460), .B(n_444), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_474), .B(n_442), .C(n_435), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_467), .A2(n_433), .B1(n_429), .B2(n_423), .Y(n_498) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_475), .A2(n_399), .B(n_400), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_487), .B(n_399), .Y(n_500) );
INVxp67_ASAP7_75t_L g501 ( .A(n_446), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_447), .B(n_423), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_488), .B(n_432), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_467), .B(n_429), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_466), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_469), .A2(n_431), .B1(n_428), .B2(n_422), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_454), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_471), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_476), .A2(n_401), .B(n_400), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_449), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_458), .B(n_401), .Y(n_512) );
OA22x2_ASAP7_75t_L g513 ( .A1(n_456), .A2(n_421), .B1(n_418), .B2(n_23), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_463), .A2(n_421), .B1(n_418), .B2(n_25), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_459), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_453), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_480), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_454), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_473), .B(n_17), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_468), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_489), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_500), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_500), .Y(n_523) );
AOI211xp5_ASAP7_75t_L g524 ( .A1(n_491), .A2(n_465), .B(n_457), .C(n_461), .Y(n_524) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_513), .A2(n_469), .B1(n_482), .B2(n_479), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_499), .Y(n_526) );
AOI322xp5_ASAP7_75t_L g527 ( .A1(n_501), .A2(n_476), .A3(n_484), .B1(n_490), .B2(n_462), .C1(n_448), .C2(n_455), .Y(n_527) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_519), .B(n_479), .Y(n_528) );
AND2x4_ASAP7_75t_SL g529 ( .A(n_493), .B(n_468), .Y(n_529) );
OAI221xp5_ASAP7_75t_L g530 ( .A1(n_495), .A2(n_452), .B1(n_477), .B2(n_470), .C(n_481), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_513), .A2(n_485), .B1(n_472), .B2(n_486), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_497), .A2(n_486), .B1(n_483), .B2(n_27), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_496), .A2(n_20), .B(n_26), .C(n_31), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_492), .Y(n_534) );
OAI22xp33_ASAP7_75t_R g535 ( .A1(n_502), .A2(n_34), .B1(n_35), .B2(n_37), .Y(n_535) );
NOR4xp25_ASAP7_75t_L g536 ( .A(n_510), .B(n_38), .C(n_43), .D(n_45), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_507), .B(n_49), .Y(n_537) );
OAI211xp5_ASAP7_75t_L g538 ( .A1(n_505), .A2(n_51), .B(n_52), .C(n_56), .Y(n_538) );
OAI31xp33_ASAP7_75t_L g539 ( .A1(n_498), .A2(n_59), .A3(n_60), .B(n_62), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_512), .B(n_65), .Y(n_540) );
NOR3xp33_ASAP7_75t_SL g541 ( .A(n_531), .B(n_530), .C(n_514), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_524), .B(n_510), .C(n_494), .Y(n_542) );
BUFx2_ASAP7_75t_L g543 ( .A(n_528), .Y(n_543) );
AOI221x1_ASAP7_75t_L g544 ( .A1(n_537), .A2(n_498), .B1(n_509), .B2(n_515), .C(n_511), .Y(n_544) );
INVx1_ASAP7_75t_SL g545 ( .A(n_529), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_525), .A2(n_516), .B(n_517), .C(n_504), .Y(n_546) );
NAND4xp25_ASAP7_75t_L g547 ( .A(n_525), .B(n_506), .C(n_503), .D(n_521), .Y(n_547) );
AOI211xp5_ASAP7_75t_SL g548 ( .A1(n_532), .A2(n_520), .B(n_518), .C(n_508), .Y(n_548) );
AOI21xp33_ASAP7_75t_SL g549 ( .A1(n_536), .A2(n_499), .B(n_68), .Y(n_549) );
AOI211xp5_ASAP7_75t_L g550 ( .A1(n_535), .A2(n_67), .B(n_70), .C(n_71), .Y(n_550) );
AND4x1_ASAP7_75t_L g551 ( .A(n_541), .B(n_539), .C(n_533), .D(n_534), .Y(n_551) );
AOI221xp5_ASAP7_75t_L g552 ( .A1(n_543), .A2(n_523), .B1(n_522), .B2(n_526), .C(n_527), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_545), .B(n_540), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_548), .B(n_538), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g555 ( .A(n_542), .B(n_72), .C(n_74), .Y(n_555) );
OR4x2_ASAP7_75t_L g556 ( .A(n_551), .B(n_546), .C(n_547), .D(n_544), .Y(n_556) );
NAND3xp33_ASAP7_75t_SL g557 ( .A(n_552), .B(n_549), .C(n_550), .Y(n_557) );
NOR3xp33_ASAP7_75t_L g558 ( .A(n_555), .B(n_76), .C(n_78), .Y(n_558) );
AO22x2_ASAP7_75t_L g559 ( .A1(n_557), .A2(n_553), .B1(n_554), .B2(n_556), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_558), .Y(n_560) );
AND2x2_ASAP7_75t_SL g561 ( .A(n_560), .B(n_559), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_559), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_561), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_563), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_564), .Y(n_565) );
OA21x2_ASAP7_75t_L g566 ( .A1(n_565), .A2(n_562), .B(n_561), .Y(n_566) );
endmodule