module fake_jpeg_15075_n_71 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_71);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

HAxp5_ASAP7_75t_SL g11 ( 
.A(n_6),
.B(n_8),
.CON(n_11),
.SN(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_4),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_19),
.B(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_22),
.A2(n_24),
.B1(n_26),
.B2(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_21),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_15),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_32),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_18),
.C(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_33),
.B(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_11),
.B1(n_16),
.B2(n_18),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_40),
.B1(n_24),
.B2(n_17),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_20),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_27),
.A2(n_3),
.B1(n_28),
.B2(n_21),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_19),
.A2(n_23),
.B1(n_17),
.B2(n_13),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_51),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_32),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_30),
.A2(n_39),
.B1(n_37),
.B2(n_29),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_49),
.A2(n_37),
.B1(n_44),
.B2(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_56),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_40),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_57),
.B(n_58),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_60),
.B(n_63),
.Y(n_66)
);

AND2x4_ASAP7_75t_SL g62 ( 
.A(n_57),
.B(n_49),
.Y(n_62)
);

XOR2x2_ASAP7_75t_SL g65 ( 
.A(n_62),
.B(n_56),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_62),
.B(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_45),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

OAI321xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_65),
.A3(n_64),
.B1(n_66),
.B2(n_55),
.C(n_47),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_50),
.CI(n_68),
.CON(n_71),
.SN(n_71)
);


endmodule