module fake_jpeg_11716_n_156 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_156);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_SL g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_2),
.B(n_4),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_43),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_38),
.B(n_41),
.Y(n_85)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_39),
.Y(n_91)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_55),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_13),
.A2(n_4),
.B1(n_18),
.B2(n_29),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_60),
.B(n_49),
.Y(n_83)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_32),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_50),
.B(n_61),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_29),
.A2(n_18),
.B1(n_27),
.B2(n_16),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_48),
.B1(n_42),
.B2(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_22),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_21),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_14),
.B(n_16),
.C(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_20),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_31),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_31),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_26),
.B(n_45),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_91),
.C(n_68),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_64),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_70),
.B(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_89),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_65),
.B1(n_67),
.B2(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_36),
.B(n_50),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_63),
.C(n_73),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_98),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_82),
.A2(n_81),
.B1(n_83),
.B2(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_119)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_SL g125 ( 
.A(n_99),
.B(n_111),
.C(n_103),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_79),
.B1(n_78),
.B2(n_66),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_100),
.A2(n_102),
.B1(n_112),
.B2(n_101),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_78),
.B1(n_67),
.B2(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_91),
.B1(n_87),
.B2(n_74),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_108),
.A2(n_112),
.B(n_93),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_82),
.B1(n_86),
.B2(n_51),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_86),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_110),
.B(n_109),
.C(n_105),
.Y(n_118)
);

FAx1_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_96),
.CI(n_94),
.CON(n_113),
.SN(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_116),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_125),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_124),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_126),
.A2(n_119),
.B1(n_118),
.B2(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_131),
.Y(n_137)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_115),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_126),
.B1(n_121),
.B2(n_123),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_113),
.A2(n_122),
.B(n_119),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_130),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_136),
.Y(n_141)
);

NOR2xp67_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_121),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_125),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_128),
.C(n_134),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_133),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_148),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_146),
.B(n_121),
.C(n_137),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_149),
.B(n_150),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_147),
.B(n_140),
.Y(n_150)
);

NAND2x1_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_145),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_152),
.A2(n_129),
.B1(n_143),
.B2(n_149),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_134),
.B(n_153),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);


endmodule