module fake_jpeg_16722_n_277 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_16),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_7),
.B(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_21),
.Y(n_38)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_41),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_28),
.B(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_21),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_33),
.B1(n_34),
.B2(n_17),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_45),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_17),
.B1(n_27),
.B2(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_17),
.B1(n_27),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_51),
.B1(n_59),
.B2(n_35),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_41),
.A2(n_18),
.B1(n_24),
.B2(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_32),
.B1(n_18),
.B2(n_19),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_38),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_62),
.Y(n_84)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_29),
.B1(n_30),
.B2(n_25),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_30),
.B1(n_20),
.B2(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_60),
.A2(n_20),
.B1(n_29),
.B2(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_21),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_70),
.B1(n_88),
.B2(n_50),
.Y(n_92)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_46),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_87),
.B(n_0),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_85),
.Y(n_101)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_64),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_21),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_58),
.B(n_37),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_44),
.A2(n_29),
.B1(n_1),
.B2(n_5),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_31),
.B1(n_22),
.B2(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_58),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_65),
.Y(n_105)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_73),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_48),
.B1(n_63),
.B2(n_53),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_93),
.A2(n_95),
.B1(n_79),
.B2(n_72),
.Y(n_131)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_99),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_63),
.B1(n_53),
.B2(n_49),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_71),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_108),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_107),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_81),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_86),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_81),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_90),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_90),
.B(n_23),
.C(n_79),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_115),
.B(n_85),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_120),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_89),
.B1(n_80),
.B2(n_88),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_123),
.B1(n_95),
.B2(n_135),
.Y(n_151)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_79),
.B(n_72),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_124),
.A2(n_139),
.B(n_94),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g126 ( 
.A1(n_101),
.A2(n_44),
.B(n_36),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_100),
.B(n_113),
.Y(n_163)
);

XNOR2x1_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_84),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_97),
.C(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_109),
.B1(n_86),
.B2(n_83),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_133),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_104),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_103),
.A2(n_76),
.B(n_39),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_151),
.A2(n_169),
.B1(n_132),
.B2(n_134),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_105),
.C(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_112),
.C(n_108),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_31),
.B(n_1),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_98),
.Y(n_158)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_72),
.B1(n_109),
.B2(n_69),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_164),
.B1(n_167),
.B2(n_141),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_163),
.A2(n_165),
.B(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_123),
.A2(n_109),
.B1(n_65),
.B2(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_111),
.Y(n_168)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_168),
.B(n_126),
.CI(n_124),
.CON(n_181),
.SN(n_181)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_123),
.A2(n_83),
.B1(n_61),
.B2(n_102),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_171),
.B(n_186),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_158),
.A2(n_124),
.B(n_137),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_177),
.B(n_178),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_165),
.A2(n_124),
.B(n_116),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_179),
.A2(n_184),
.B1(n_185),
.B2(n_187),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_159),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_124),
.B1(n_126),
.B2(n_133),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_120),
.B1(n_102),
.B2(n_125),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_168),
.A2(n_102),
.B1(n_141),
.B2(n_130),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_152),
.B1(n_149),
.B2(n_160),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_142),
.A2(n_12),
.B(n_1),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_154),
.B1(n_146),
.B2(n_6),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_148),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_198),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_142),
.C(n_153),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_199),
.C(n_204),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_189),
.B(n_147),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_163),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_201),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_163),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_199),
.Y(n_223)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_207),
.Y(n_215)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_167),
.B1(n_164),
.B2(n_154),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_211),
.B1(n_185),
.B2(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_214),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_172),
.A2(n_157),
.B1(n_155),
.B2(n_150),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_143),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_191),
.B(n_179),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_217),
.A2(n_9),
.B(n_5),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_195),
.A2(n_173),
.B1(n_175),
.B2(n_170),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_219),
.A2(n_221),
.B1(n_231),
.B2(n_0),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_208),
.B1(n_213),
.B2(n_212),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_227),
.Y(n_242)
);

INVx13_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_225),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_39),
.B(n_23),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_181),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_181),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_198),
.C(n_204),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_183),
.B1(n_188),
.B2(n_150),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_234),
.C(n_235),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_202),
.C(n_210),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_194),
.C(n_61),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_243),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_222),
.B(n_228),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_241),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_15),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_220),
.C(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_215),
.B(n_9),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_236),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_217),
.B(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_250),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_234),
.A2(n_220),
.B1(n_231),
.B2(n_229),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_226),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_236),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_257),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_246),
.A2(n_240),
.B(n_242),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_242),
.B(n_232),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_260),
.C(n_9),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_259),
.B(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_230),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_249),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g269 ( 
.A1(n_263),
.A2(n_268),
.A3(n_11),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_247),
.B(n_252),
.Y(n_264)
);

NAND3xp33_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_12),
.C(n_13),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_7),
.C(n_11),
.Y(n_270)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_270),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_272),
.B1(n_13),
.B2(n_14),
.Y(n_273)
);

AOI321xp33_ASAP7_75t_SL g272 ( 
.A1(n_266),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_0),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_264),
.B(n_274),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_265),
.C(n_15),
.Y(n_277)
);


endmodule