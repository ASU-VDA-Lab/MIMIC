module fake_ibex_170_n_1009 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_181, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_182, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_1009);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_182;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_1009;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_992;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_926;
wire n_328;
wire n_372;
wire n_341;
wire n_293;
wire n_418;
wire n_256;
wire n_510;
wire n_193;
wire n_845;
wire n_947;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_994;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_909;
wire n_545;
wire n_862;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_991;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_996;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_698;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_708;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_196;
wire n_327;
wire n_326;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_497;
wire n_243;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_989;
wire n_373;
wire n_854;
wire n_1008;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_987;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_281;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_490;
wire n_407;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_1001;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_543;
wire n_420;
wire n_483;
wire n_580;
wire n_769;
wire n_487;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_993;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_999;
wire n_560;
wire n_429;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_1004;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_433;
wire n_439;
wire n_704;
wire n_949;
wire n_1007;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_1006;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_998;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_918;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_567;
wire n_548;
wire n_516;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_986;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_990;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_712;
wire n_451;
wire n_702;
wire n_971;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_1002;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_320;
wire n_285;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_997;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_588;
wire n_212;
wire n_513;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_1005;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_450;
wire n_302;
wire n_443;
wire n_686;
wire n_985;
wire n_572;
wire n_867;
wire n_983;
wire n_1003;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_921;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_995;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_1000;
wire n_364;
wire n_687;
wire n_895;
wire n_988;
wire n_298;
wire n_231;
wire n_202;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_71),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_58),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_86),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_2),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_57),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_23),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_22),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_148),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_64),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_68),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_100),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_43),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_62),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_130),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_76),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_81),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_96),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_14),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_10),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_27),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_137),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_22),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_141),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_134),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_67),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_42),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_66),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_179),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_170),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_19),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_45),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_29),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_102),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_10),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g235 ( 
.A(n_89),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_129),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_119),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_160),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_44),
.Y(n_239)
);

BUFx8_ASAP7_75t_SL g240 ( 
.A(n_46),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_120),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_65),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_79),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_92),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_94),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_97),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_132),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_146),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_38),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_23),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_55),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_82),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_98),
.B(n_56),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_108),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_153),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_L g260 ( 
.A(n_90),
.B(n_19),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_113),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_41),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_133),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_99),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_53),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_74),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_59),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_128),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_145),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_85),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_84),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_0),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_38),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_88),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_93),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_110),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_40),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_33),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_3),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_39),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_111),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_63),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_73),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_34),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_L g285 ( 
.A(n_17),
.B(n_163),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_20),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_171),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_61),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_95),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_117),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_70),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_112),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_180),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_15),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_121),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_174),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g297 ( 
.A(n_24),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_138),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_11),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_8),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_101),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_83),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_80),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_169),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_91),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_175),
.Y(n_306)
);

INVx5_ASAP7_75t_L g307 ( 
.A(n_191),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_201),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_235),
.B(n_0),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_235),
.B(n_1),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_279),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_200),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_286),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

NOR2x1_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_1),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_185),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_201),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_186),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_191),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_284),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_200),
.B(n_2),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_187),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_191),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_189),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_216),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_298),
.B(n_3),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_240),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_194),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_193),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_197),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_274),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_216),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_198),
.Y(n_339)
);

BUFx8_ASAP7_75t_L g340 ( 
.A(n_257),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

INVx6_ASAP7_75t_L g342 ( 
.A(n_274),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_242),
.Y(n_343)
);

BUFx12f_ASAP7_75t_L g344 ( 
.A(n_183),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_270),
.Y(n_345)
);

NAND2xp33_ASAP7_75t_L g346 ( 
.A(n_288),
.B(n_290),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_270),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_288),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_291),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_291),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_288),
.Y(n_351)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_246),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_246),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_199),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_203),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_204),
.Y(n_356)
);

AND2x4_ASAP7_75t_L g357 ( 
.A(n_208),
.B(n_5),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_240),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_205),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_209),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_210),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_290),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_196),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_212),
.B(n_263),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_290),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_218),
.Y(n_366)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_217),
.B(n_6),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_219),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_222),
.B(n_7),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

INVx5_ASAP7_75t_L g371 ( 
.A(n_290),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_238),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_194),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_231),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_239),
.Y(n_375)
);

BUFx8_ASAP7_75t_L g376 ( 
.A(n_295),
.Y(n_376)
);

BUFx12f_ASAP7_75t_L g377 ( 
.A(n_184),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_243),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_244),
.Y(n_379)
);

OA21x2_ASAP7_75t_L g380 ( 
.A1(n_245),
.A2(n_87),
.B(n_178),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_214),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_295),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_249),
.B(n_16),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_332),
.B(n_190),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_SL g385 ( 
.A(n_311),
.B(n_207),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_316),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_342),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

INVx8_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_357),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_323),
.B(n_248),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_323),
.B(n_251),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_332),
.B(n_215),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

INVxp33_ASAP7_75t_SL g398 ( 
.A(n_364),
.Y(n_398)
);

BUFx6f_ASAP7_75t_SL g399 ( 
.A(n_357),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_363),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_341),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_341),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_363),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_330),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_367),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_310),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_316),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_332),
.B(n_229),
.Y(n_412)
);

AND3x2_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_297),
.C(n_256),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_336),
.B(n_342),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_336),
.B(n_234),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_309),
.B(n_272),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_310),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_313),
.Y(n_420)
);

NAND2xp33_ASAP7_75t_SL g421 ( 
.A(n_311),
.B(n_312),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_316),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_369),
.A2(n_278),
.B1(n_280),
.B2(n_277),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_321),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_323),
.B(n_252),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_321),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_315),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_321),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_315),
.Y(n_430)
);

NAND2xp33_ASAP7_75t_L g431 ( 
.A(n_318),
.B(n_295),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_321),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_309),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_369),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_322),
.B(n_250),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_308),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_318),
.B(n_259),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_308),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_L g439 ( 
.A(n_320),
.B(n_295),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_325),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_L g441 ( 
.A1(n_331),
.A2(n_220),
.B1(n_214),
.B2(n_207),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_376),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_325),
.Y(n_443)
);

AOI22xp33_ASAP7_75t_L g444 ( 
.A1(n_333),
.A2(n_294),
.B1(n_300),
.B2(n_299),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_325),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_342),
.B(n_324),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_319),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_344),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_353),
.B(n_261),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_324),
.B(n_266),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_326),
.B(n_188),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_326),
.B(n_267),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_319),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_330),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_353),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_325),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_358),
.B(n_262),
.Y(n_457)
);

BUFx6f_ASAP7_75t_SL g458 ( 
.A(n_335),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_343),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_343),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_325),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_335),
.B(n_339),
.Y(n_462)
);

OR2x6_ASAP7_75t_L g463 ( 
.A(n_373),
.B(n_260),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_339),
.B(n_271),
.Y(n_464)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_353),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_328),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_355),
.B(n_192),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_356),
.B(n_275),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_328),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_337),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_337),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_338),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_338),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_358),
.B(n_306),
.Y(n_474)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_329),
.B(n_224),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_356),
.B(n_372),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_372),
.B(n_285),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g478 ( 
.A1(n_354),
.A2(n_282),
.B1(n_289),
.B2(n_293),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_377),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_354),
.B(n_195),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_345),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g482 ( 
.A(n_373),
.B(n_264),
.C(n_206),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_345),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_347),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_347),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_343),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_349),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_348),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_377),
.B(n_220),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_359),
.B(n_360),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_349),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_348),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_359),
.B(n_202),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_352),
.B(n_211),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_340),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_350),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_340),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_348),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_350),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_446),
.B(n_340),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g503 ( 
.A(n_417),
.B(n_331),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_486),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_442),
.Y(n_506)
);

NAND2xp33_ASAP7_75t_L g507 ( 
.A(n_449),
.B(n_213),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_384),
.B(n_340),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_479),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_317),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_446),
.B(n_314),
.Y(n_512)
);

O2A1O1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_434),
.A2(n_383),
.B(n_374),
.C(n_368),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_486),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_413),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_451),
.B(n_467),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_395),
.B(n_360),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_458),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_402),
.B(n_221),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_414),
.B(n_314),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_459),
.Y(n_522)
);

A2O1A1Ixp33_ASAP7_75t_L g523 ( 
.A1(n_476),
.A2(n_408),
.B(n_409),
.C(n_421),
.Y(n_523)
);

BUFx6f_ASAP7_75t_SL g524 ( 
.A(n_448),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_412),
.B(n_361),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_414),
.B(n_352),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_401),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_458),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_435),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_416),
.B(n_366),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_421),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_462),
.B(n_370),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_399),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_460),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_462),
.B(n_375),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_391),
.B(n_223),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_465),
.B(n_375),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_465),
.B(n_391),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_491),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_444),
.B(n_378),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_415),
.A2(n_379),
.B1(n_317),
.B2(n_381),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_489),
.B(n_381),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_493),
.B(n_379),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_460),
.Y(n_546)
);

AOI22xp33_ASAP7_75t_L g547 ( 
.A1(n_415),
.A2(n_380),
.B1(n_376),
.B2(n_224),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g548 ( 
.A1(n_392),
.A2(n_425),
.B(n_393),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_449),
.B(n_225),
.Y(n_549)
);

AO221x1_ASAP7_75t_L g550 ( 
.A1(n_441),
.A2(n_281),
.B1(n_232),
.B2(n_376),
.C(n_365),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_398),
.B(n_226),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_401),
.B(n_232),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_398),
.A2(n_281),
.B1(n_227),
.B2(n_276),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_423),
.B(n_388),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_399),
.B(n_228),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_457),
.B(n_230),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_474),
.B(n_233),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_392),
.B(n_237),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_499),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_477),
.B(n_247),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_477),
.B(n_253),
.Y(n_561)
);

AOI33xp33_ASAP7_75t_L g562 ( 
.A1(n_478),
.A2(n_477),
.A3(n_410),
.B1(n_418),
.B2(n_430),
.B3(n_419),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g563 ( 
.A(n_475),
.B(n_380),
.C(n_296),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

BUFx5_ASAP7_75t_L g565 ( 
.A(n_449),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_494),
.B(n_254),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_437),
.B(n_450),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_437),
.B(n_255),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_406),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_420),
.B(n_258),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_495),
.A2(n_302),
.B1(n_265),
.B2(n_268),
.Y(n_571)
);

NOR2x1p5_ASAP7_75t_L g572 ( 
.A(n_454),
.B(n_269),
.Y(n_572)
);

O2A1O1Ixp5_ASAP7_75t_L g573 ( 
.A1(n_452),
.A2(n_380),
.B(n_346),
.C(n_371),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_427),
.A2(n_380),
.B1(n_382),
.B2(n_351),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_438),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_490),
.Y(n_576)
);

O2A1O1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_464),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_468),
.B(n_283),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_495),
.B(n_287),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_475),
.B(n_18),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_466),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_480),
.B(n_292),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_469),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_470),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_385),
.B(n_21),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_385),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_471),
.B(n_301),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_472),
.B(n_303),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_473),
.B(n_304),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_481),
.B(n_305),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_483),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_484),
.B(n_307),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_485),
.B(n_24),
.Y(n_595)
);

O2A1O1Ixp5_ASAP7_75t_L g596 ( 
.A1(n_490),
.A2(n_371),
.B(n_362),
.C(n_307),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_487),
.Y(n_597)
);

AO22x1_ASAP7_75t_L g598 ( 
.A1(n_527),
.A2(n_482),
.B1(n_463),
.B2(n_496),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_524),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_517),
.A2(n_439),
.B(n_431),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_529),
.A2(n_463),
.B1(n_480),
.B2(n_407),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_588),
.A2(n_531),
.B1(n_500),
.B2(n_501),
.Y(n_602)
);

OAI22x1_ASAP7_75t_L g603 ( 
.A1(n_552),
.A2(n_463),
.B1(n_26),
.B2(n_28),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_542),
.B(n_25),
.Y(n_604)
);

AOI221xp5_ASAP7_75t_L g605 ( 
.A1(n_513),
.A2(n_389),
.B1(n_404),
.B2(n_403),
.C(n_400),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_519),
.B(n_25),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_501),
.Y(n_607)
);

AO21x1_ASAP7_75t_L g608 ( 
.A1(n_577),
.A2(n_394),
.B(n_386),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_504),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g610 ( 
.A(n_500),
.B(n_396),
.C(n_394),
.Y(n_610)
);

INVxp67_ASAP7_75t_SL g611 ( 
.A(n_504),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_R g612 ( 
.A(n_569),
.B(n_26),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_540),
.A2(n_397),
.B(n_400),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_524),
.Y(n_614)
);

AOI21xp33_ASAP7_75t_L g615 ( 
.A1(n_551),
.A2(n_508),
.B(n_503),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_588),
.A2(n_531),
.B1(n_511),
.B2(n_567),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_511),
.B(n_28),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_573),
.A2(n_403),
.B(n_498),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_556),
.B(n_29),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_506),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_575),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_526),
.A2(n_521),
.B(n_512),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_553),
.B(n_30),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_580),
.B(n_30),
.Y(n_624)
);

AO21x1_ASAP7_75t_L g625 ( 
.A1(n_577),
.A2(n_525),
.B(n_502),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_557),
.B(n_31),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_523),
.B(n_31),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_595),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_518),
.B(n_32),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_539),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_519),
.B(n_32),
.Y(n_631)
);

AO22x1_ASAP7_75t_L g632 ( 
.A1(n_528),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_632)
);

BUFx4f_ASAP7_75t_L g633 ( 
.A(n_587),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_506),
.Y(n_634)
);

AOI21x1_ASAP7_75t_L g635 ( 
.A1(n_548),
.A2(n_492),
.B(n_488),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_564),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_530),
.B(n_35),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_562),
.B(n_36),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_560),
.B(n_36),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_510),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_528),
.B(n_37),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_506),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_547),
.A2(n_307),
.B1(n_362),
.B2(n_371),
.Y(n_643)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_513),
.A2(n_382),
.B(n_362),
.C(n_371),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_509),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_579),
.B(n_37),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_538),
.A2(n_461),
.B(n_456),
.Y(n_647)
);

NOR2x1_ASAP7_75t_L g648 ( 
.A(n_533),
.B(n_456),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_597),
.B(n_39),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_563),
.A2(n_574),
.B(n_536),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_583),
.B(n_586),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_561),
.B(n_40),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_593),
.B(n_582),
.Y(n_653)
);

CKINVDCx10_ASAP7_75t_R g654 ( 
.A(n_544),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_594),
.A2(n_532),
.B(n_514),
.Y(n_655)
);

O2A1O1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_581),
.A2(n_445),
.B(n_443),
.C(n_440),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_547),
.A2(n_509),
.B1(n_543),
.B2(n_585),
.Y(n_657)
);

NAND2x1p5_ASAP7_75t_L g658 ( 
.A(n_533),
.B(n_307),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_545),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_554),
.B(n_558),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_571),
.Y(n_661)
);

NOR2x1_ASAP7_75t_L g662 ( 
.A(n_572),
.B(n_445),
.Y(n_662)
);

A2O1A1Ixp33_ASAP7_75t_L g663 ( 
.A1(n_576),
.A2(n_382),
.B(n_362),
.C(n_371),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g664 ( 
.A1(n_574),
.A2(n_443),
.B(n_440),
.Y(n_664)
);

OAI22x1_ASAP7_75t_L g665 ( 
.A1(n_550),
.A2(n_371),
.B1(n_362),
.B2(n_49),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_515),
.B(n_47),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_543),
.B(n_48),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_555),
.B(n_51),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_SL g669 ( 
.A1(n_566),
.A2(n_432),
.B(n_429),
.C(n_426),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_584),
.B(n_52),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_568),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_505),
.A2(n_424),
.B(n_422),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_590),
.A2(n_592),
.B(n_516),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_520),
.B(n_54),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_522),
.A2(n_428),
.B(n_411),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_534),
.A2(n_535),
.B(n_546),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_570),
.B(n_537),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_559),
.Y(n_679)
);

BUFx12f_ASAP7_75t_L g680 ( 
.A(n_589),
.Y(n_680)
);

INVx6_ASAP7_75t_L g681 ( 
.A(n_565),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_591),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_578),
.Y(n_683)
);

AOI211x1_ASAP7_75t_L g684 ( 
.A1(n_625),
.A2(n_596),
.B(n_549),
.C(n_507),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_616),
.B(n_565),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_615),
.B(n_565),
.Y(n_686)
);

AO22x2_ASAP7_75t_L g687 ( 
.A1(n_657),
.A2(n_565),
.B1(n_60),
.B2(n_69),
.Y(n_687)
);

OA22x2_ASAP7_75t_L g688 ( 
.A1(n_641),
.A2(n_631),
.B1(n_606),
.B2(n_603),
.Y(n_688)
);

INVx4_ASAP7_75t_SL g689 ( 
.A(n_641),
.Y(n_689)
);

NAND3xp33_ASAP7_75t_SL g690 ( 
.A(n_612),
.B(n_72),
.C(n_75),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_640),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_673),
.A2(n_387),
.B(n_78),
.Y(n_692)
);

BUFx2_ASAP7_75t_SL g693 ( 
.A(n_620),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_634),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_636),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_651),
.A2(n_103),
.B(n_104),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_646),
.Y(n_697)
);

OAI22xp5_ASAP7_75t_L g698 ( 
.A1(n_633),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_660),
.A2(n_109),
.B(n_115),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_628),
.B(n_118),
.Y(n_700)
);

AOI21xp33_ASAP7_75t_L g701 ( 
.A1(n_661),
.A2(n_123),
.B(n_124),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_602),
.B(n_126),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_599),
.Y(n_703)
);

OA21x2_ASAP7_75t_L g704 ( 
.A1(n_664),
.A2(n_135),
.B(n_136),
.Y(n_704)
);

A2O1A1Ixp33_ASAP7_75t_L g705 ( 
.A1(n_627),
.A2(n_139),
.B(n_140),
.C(n_142),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_620),
.B(n_144),
.Y(n_706)
);

AOI21xp5_ASAP7_75t_L g707 ( 
.A1(n_613),
.A2(n_653),
.B(n_672),
.Y(n_707)
);

AO32x2_ASAP7_75t_L g708 ( 
.A1(n_643),
.A2(n_147),
.A3(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_598),
.B(n_155),
.C(n_156),
.Y(n_709)
);

OAI21x1_ASAP7_75t_L g710 ( 
.A1(n_676),
.A2(n_157),
.B(n_158),
.Y(n_710)
);

OAI221xp5_ASAP7_75t_L g711 ( 
.A1(n_601),
.A2(n_182),
.B1(n_164),
.B2(n_166),
.C(n_167),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_604),
.A2(n_172),
.B1(n_637),
.B2(n_629),
.Y(n_712)
);

NOR2x1_ASAP7_75t_R g713 ( 
.A(n_614),
.B(n_680),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_654),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_623),
.B(n_631),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_606),
.B(n_624),
.Y(n_716)
);

OAI21x1_ASAP7_75t_SL g717 ( 
.A1(n_638),
.A2(n_668),
.B(n_649),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_671),
.B(n_617),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_659),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_619),
.B(n_626),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_620),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_683),
.B(n_678),
.Y(n_722)
);

NOR2xp33_ASAP7_75t_L g723 ( 
.A(n_682),
.B(n_652),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_674),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_621),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_658),
.Y(n_726)
);

OAI21xp5_ASAP7_75t_L g727 ( 
.A1(n_656),
.A2(n_600),
.B(n_647),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_632),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_667),
.B(n_639),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_610),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_662),
.B(n_611),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_648),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_645),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_642),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_609),
.B(n_645),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_645),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_679),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_609),
.B(n_666),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_605),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_670),
.A2(n_675),
.B(n_669),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_663),
.A2(n_681),
.B(n_679),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_681),
.B(n_531),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_635),
.A2(n_655),
.B(n_618),
.Y(n_743)
);

AO31x2_ASAP7_75t_L g744 ( 
.A1(n_608),
.A2(n_625),
.A3(n_644),
.B(n_665),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_616),
.B(n_531),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_633),
.A2(n_630),
.B1(n_651),
.B2(n_653),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_607),
.Y(n_747)
);

OAI21x1_ASAP7_75t_L g748 ( 
.A1(n_635),
.A2(n_655),
.B(n_618),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_616),
.B(n_531),
.Y(n_749)
);

OA21x2_ASAP7_75t_L g750 ( 
.A1(n_650),
.A2(n_574),
.B(n_573),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_640),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_616),
.B(n_531),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_616),
.B(n_531),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_636),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_616),
.B(n_531),
.Y(n_755)
);

INVx3_ASAP7_75t_L g756 ( 
.A(n_645),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_616),
.B(n_531),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_622),
.A2(n_650),
.B(n_523),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_635),
.A2(n_655),
.B(n_618),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_665),
.B(n_533),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_644),
.B(n_547),
.C(n_563),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_616),
.B(n_531),
.Y(n_762)
);

OAI21x1_ASAP7_75t_SL g763 ( 
.A1(n_651),
.A2(n_638),
.B(n_677),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_616),
.B(n_531),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_673),
.A2(n_622),
.B(n_517),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_673),
.A2(n_622),
.B(n_517),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_607),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_657),
.A2(n_421),
.B1(n_550),
.B2(n_661),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_616),
.B(n_531),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_640),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_616),
.B(n_531),
.Y(n_771)
);

AO31x2_ASAP7_75t_L g772 ( 
.A1(n_608),
.A2(n_625),
.A3(n_644),
.B(n_665),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_634),
.Y(n_773)
);

AO31x2_ASAP7_75t_L g774 ( 
.A1(n_608),
.A2(n_625),
.A3(n_644),
.B(n_665),
.Y(n_774)
);

A2O1A1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_673),
.A2(n_615),
.B(n_525),
.C(n_508),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_747),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_751),
.Y(n_777)
);

HB1xp67_ASAP7_75t_L g778 ( 
.A(n_747),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_695),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_691),
.B(n_703),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_754),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_767),
.B(n_715),
.Y(n_782)
);

NAND2x1p5_ASAP7_75t_L g783 ( 
.A(n_726),
.B(n_733),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_758),
.A2(n_761),
.B(n_739),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_725),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_728),
.Y(n_786)
);

BUFx3_ASAP7_75t_L g787 ( 
.A(n_770),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_714),
.Y(n_788)
);

AO32x2_ASAP7_75t_L g789 ( 
.A1(n_746),
.A2(n_698),
.A3(n_712),
.B1(n_744),
.B2(n_772),
.Y(n_789)
);

INVx8_ASAP7_75t_L g790 ( 
.A(n_694),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_689),
.Y(n_791)
);

OAI21xp5_ASAP7_75t_L g792 ( 
.A1(n_758),
.A2(n_761),
.B(n_707),
.Y(n_792)
);

OAI21xp5_ASAP7_75t_L g793 ( 
.A1(n_768),
.A2(n_686),
.B(n_727),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_730),
.Y(n_794)
);

INVx2_ASAP7_75t_SL g795 ( 
.A(n_689),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_693),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_688),
.A2(n_729),
.B1(n_716),
.B2(n_720),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_697),
.A2(n_718),
.B1(n_722),
.B2(n_723),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_724),
.B(n_760),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_768),
.A2(n_687),
.B1(n_749),
.B2(n_745),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_737),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_SL g802 ( 
.A1(n_705),
.A2(n_701),
.B(n_706),
.C(n_690),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_736),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_752),
.B(n_755),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_753),
.B(n_764),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_721),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_717),
.A2(n_750),
.B(n_692),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_735),
.B(n_757),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_685),
.A2(n_762),
.B(n_771),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_732),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_769),
.B(n_756),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_700),
.Y(n_812)
);

OAI221xp5_ASAP7_75t_SL g813 ( 
.A1(n_711),
.A2(n_709),
.B1(n_702),
.B2(n_738),
.C(n_731),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_742),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_744),
.B(n_774),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_744),
.Y(n_816)
);

INVx2_ASAP7_75t_SL g817 ( 
.A(n_734),
.Y(n_817)
);

AO31x2_ASAP7_75t_L g818 ( 
.A1(n_699),
.A2(n_774),
.A3(n_772),
.B(n_696),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_773),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_710),
.A2(n_741),
.B(n_740),
.Y(n_820)
);

OAI211xp5_ASAP7_75t_L g821 ( 
.A1(n_684),
.A2(n_704),
.B(n_708),
.C(n_713),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_713),
.B(n_684),
.Y(n_822)
);

AOI222xp33_ASAP7_75t_L g823 ( 
.A1(n_708),
.A2(n_373),
.B1(n_381),
.B2(n_441),
.C1(n_543),
.C2(n_689),
.Y(n_823)
);

A2O1A1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_775),
.A2(n_768),
.B(n_766),
.C(n_765),
.Y(n_824)
);

AOI221xp5_ASAP7_75t_L g825 ( 
.A1(n_754),
.A2(n_615),
.B1(n_441),
.B2(n_543),
.C(n_513),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_775),
.A2(n_766),
.B(n_765),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_747),
.Y(n_827)
);

BUFx4f_ASAP7_75t_L g828 ( 
.A(n_691),
.Y(n_828)
);

BUFx2_ASAP7_75t_L g829 ( 
.A(n_751),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_695),
.Y(n_830)
);

OA21x2_ASAP7_75t_L g831 ( 
.A1(n_743),
.A2(n_759),
.B(n_748),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_695),
.Y(n_832)
);

BUFx2_ASAP7_75t_L g833 ( 
.A(n_751),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_747),
.B(n_527),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_739),
.B(n_719),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_695),
.Y(n_836)
);

OAI21x1_ASAP7_75t_SL g837 ( 
.A1(n_746),
.A2(n_763),
.B(n_717),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_695),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_726),
.B(n_620),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_693),
.B(n_641),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_786),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_831),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_776),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_825),
.A2(n_824),
.B(n_813),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_781),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_825),
.B(n_835),
.Y(n_846)
);

BUFx2_ASAP7_75t_SL g847 ( 
.A(n_791),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_808),
.B(n_811),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_785),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_840),
.A2(n_797),
.B1(n_798),
.B2(n_800),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_816),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_796),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_778),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_835),
.B(n_804),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_788),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_839),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_794),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_826),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_840),
.A2(n_800),
.B1(n_827),
.B2(n_804),
.Y(n_859)
);

CKINVDCx11_ASAP7_75t_R g860 ( 
.A(n_829),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_840),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_790),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_837),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_779),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_830),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_806),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_832),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_839),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_836),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_790),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_819),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_823),
.A2(n_805),
.B1(n_822),
.B2(n_814),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_822),
.B(n_799),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_782),
.B(n_838),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_809),
.B(n_784),
.Y(n_875)
);

AO21x2_ASAP7_75t_L g876 ( 
.A1(n_807),
.A2(n_792),
.B(n_820),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_777),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_834),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_809),
.B(n_784),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_790),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_L g881 ( 
.A1(n_823),
.A2(n_812),
.B1(n_828),
.B2(n_799),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_815),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_783),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_815),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_793),
.B(n_803),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_842),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_843),
.Y(n_887)
);

INVxp67_ASAP7_75t_L g888 ( 
.A(n_843),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_851),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_882),
.B(n_884),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_875),
.B(n_792),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_853),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_875),
.B(n_879),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_871),
.Y(n_894)
);

INVx4_ASAP7_75t_R g895 ( 
.A(n_856),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_879),
.B(n_789),
.Y(n_896)
);

BUFx12f_ASAP7_75t_L g897 ( 
.A(n_877),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_874),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_874),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_850),
.A2(n_833),
.B1(n_795),
.B2(n_810),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_858),
.B(n_818),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_846),
.B(n_854),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_885),
.B(n_821),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_866),
.B(n_787),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_871),
.Y(n_905)
);

INVxp67_ASAP7_75t_L g906 ( 
.A(n_859),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_904),
.B(n_860),
.Y(n_907)
);

NAND2x1_ASAP7_75t_L g908 ( 
.A(n_895),
.B(n_873),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_889),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_893),
.B(n_876),
.Y(n_910)
);

NOR2xp67_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_861),
.Y(n_911)
);

INVxp67_ASAP7_75t_SL g912 ( 
.A(n_905),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_897),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_893),
.B(n_876),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_898),
.B(n_841),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_899),
.B(n_893),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_891),
.B(n_876),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_890),
.B(n_863),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_891),
.B(n_848),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_892),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_887),
.B(n_857),
.Y(n_921)
);

NAND2x1_ASAP7_75t_L g922 ( 
.A(n_895),
.B(n_873),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_886),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_896),
.B(n_848),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_897),
.B(n_828),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_905),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_894),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_887),
.B(n_873),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_896),
.B(n_848),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_902),
.B(n_845),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_910),
.B(n_896),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_918),
.B(n_890),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_916),
.B(n_910),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_926),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_920),
.B(n_890),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_914),
.B(n_901),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_923),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_909),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_927),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_930),
.B(n_888),
.Y(n_940)
);

NAND2xp33_ASAP7_75t_L g941 ( 
.A(n_913),
.B(n_900),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_915),
.B(n_888),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_914),
.B(n_903),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_917),
.B(n_903),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_917),
.B(n_924),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_919),
.B(n_906),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_933),
.B(n_921),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_932),
.A2(n_911),
.B1(n_922),
.B2(n_908),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_937),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_936),
.B(n_924),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_938),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_938),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_942),
.B(n_907),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_945),
.B(n_929),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_933),
.B(n_921),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_943),
.B(n_927),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_941),
.A2(n_872),
.B1(n_906),
.B2(n_881),
.Y(n_957)
);

OR2x2_ASAP7_75t_L g958 ( 
.A(n_943),
.B(n_912),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_945),
.B(n_936),
.Y(n_959)
);

AOI222xp33_ASAP7_75t_L g960 ( 
.A1(n_941),
.A2(n_844),
.B1(n_902),
.B2(n_925),
.C1(n_878),
.C2(n_845),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_947),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_953),
.B(n_946),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_949),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_955),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_959),
.B(n_931),
.Y(n_965)
);

NOR4xp25_ASAP7_75t_L g966 ( 
.A(n_956),
.B(n_849),
.C(n_940),
.D(n_934),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_951),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_952),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_958),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_950),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_960),
.A2(n_932),
.B1(n_935),
.B2(n_872),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_963),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_962),
.A2(n_948),
.B(n_908),
.C(n_922),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_966),
.A2(n_960),
.B(n_939),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_970),
.B(n_931),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_971),
.A2(n_957),
.B(n_894),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_974),
.A2(n_962),
.B(n_969),
.C(n_852),
.Y(n_977)
);

OAI221xp5_ASAP7_75t_L g978 ( 
.A1(n_973),
.A2(n_957),
.B1(n_964),
.B2(n_961),
.C(n_968),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_976),
.A2(n_967),
.B1(n_965),
.B2(n_963),
.C(n_954),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_979),
.B(n_975),
.Y(n_980)
);

NAND4xp75_ASAP7_75t_L g981 ( 
.A(n_977),
.B(n_780),
.C(n_852),
.D(n_847),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_981),
.B(n_972),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_980),
.B(n_978),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_982),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_983),
.B(n_877),
.Y(n_985)
);

XOR2xp5_ASAP7_75t_L g986 ( 
.A(n_984),
.B(n_855),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_985),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_986),
.Y(n_988)
);

OR2x6_ASAP7_75t_L g989 ( 
.A(n_987),
.B(n_847),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_986),
.B(n_877),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_988),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_989),
.Y(n_992)
);

XOR2x2_ASAP7_75t_L g993 ( 
.A(n_990),
.B(n_877),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_988),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_989),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_995),
.A2(n_868),
.B1(n_856),
.B2(n_883),
.Y(n_996)
);

OAI22x1_ASAP7_75t_L g997 ( 
.A1(n_991),
.A2(n_783),
.B1(n_862),
.B2(n_870),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_L g998 ( 
.A(n_994),
.B(n_991),
.C(n_992),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_993),
.B(n_849),
.Y(n_999)
);

OA21x2_ASAP7_75t_L g1000 ( 
.A1(n_994),
.A2(n_862),
.B(n_870),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_991),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_995),
.B(n_857),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_1001),
.A2(n_868),
.B1(n_880),
.B2(n_944),
.Y(n_1003)
);

OA22x2_ASAP7_75t_L g1004 ( 
.A1(n_997),
.A2(n_880),
.B1(n_873),
.B2(n_928),
.Y(n_1004)
);

AO221x1_ASAP7_75t_L g1005 ( 
.A1(n_996),
.A2(n_880),
.B1(n_869),
.B2(n_867),
.C(n_864),
.Y(n_1005)
);

OAI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_1003),
.A2(n_998),
.B1(n_1000),
.B2(n_1002),
.C(n_999),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_1006),
.B(n_1005),
.Y(n_1007)
);

OA22x2_ASAP7_75t_L g1008 ( 
.A1(n_1007),
.A2(n_1004),
.B1(n_801),
.B2(n_865),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_1008),
.A2(n_802),
.B(n_817),
.Y(n_1009)
);


endmodule