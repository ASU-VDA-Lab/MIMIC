module fake_jpeg_20821_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_37;
wire n_29;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

OR2x2_ASAP7_75t_SL g8 ( 
.A(n_3),
.B(n_4),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx16_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_SL g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_15),
.B(n_16),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2xp33_ASAP7_75t_SL g26 ( 
.A(n_18),
.B(n_20),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_21),
.B1(n_12),
.B2(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_9),
.A2(n_5),
.B1(n_6),
.B2(n_0),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_10),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_10),
.B(n_11),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_30),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_11),
.B(n_13),
.Y(n_24)
);

XOR2x1_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_15),
.B(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_27),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_37),
.Y(n_42)
);

AO21x1_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_17),
.B(n_22),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_29),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_26),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_41),
.A2(n_36),
.B1(n_31),
.B2(n_14),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.C(n_45),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_40),
.C(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_47),
.Y(n_50)
);


endmodule