module fake_jpeg_3609_n_241 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_241);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_241;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_8),
.B(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_39),
.B(n_46),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_21),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_25),
.B(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_23),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_30),
.B1(n_16),
.B2(n_38),
.Y(n_71)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_55),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_34),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx9p33_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_63),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_21),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_18),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_71),
.A2(n_68),
.B1(n_65),
.B2(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_72),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_17),
.B1(n_32),
.B2(n_22),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_90),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_16),
.B1(n_30),
.B2(n_38),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_99),
.B1(n_57),
.B2(n_54),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_50),
.A2(n_32),
.B1(n_22),
.B2(n_19),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_94),
.B(n_97),
.Y(n_120)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_42),
.B(n_19),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_28),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_12),
.C(n_13),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_18),
.B1(n_17),
.B2(n_35),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_40),
.B(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_101),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_35),
.B1(n_5),
.B2(n_6),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_47),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_53),
.B1(n_60),
.B2(n_40),
.Y(n_102)
);

NAND2xp33_ASAP7_75t_R g149 ( 
.A(n_102),
.B(n_111),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_89),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_112),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_75),
.B(n_53),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_106),
.B(n_109),
.C(n_79),
.Y(n_138)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_44),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_114),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_60),
.C(n_45),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_4),
.Y(n_111)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_10),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_119),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_118),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_10),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_65),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_121),
.B(n_66),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_11),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_103),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_124),
.Y(n_141)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_85),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_85),
.B(n_87),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_131),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_100),
.B1(n_70),
.B2(n_77),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_74),
.A2(n_96),
.B1(n_79),
.B2(n_84),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_130),
.A2(n_96),
.B1(n_68),
.B2(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_104),
.B1(n_120),
.B2(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_140),
.B1(n_143),
.B2(n_156),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_136),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_86),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_132),
.C(n_129),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_158),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_114),
.B1(n_112),
.B2(n_104),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_111),
.B(n_109),
.CI(n_113),
.CON(n_146),
.SN(n_146)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_146),
.B(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_108),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_150),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_115),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_152),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_155),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_110),
.A2(n_84),
.B1(n_88),
.B2(n_70),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_77),
.B1(n_100),
.B2(n_69),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_69),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_119),
.A2(n_116),
.B1(n_102),
.B2(n_128),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_171),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_106),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_168),
.B(n_178),
.C(n_180),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_176),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_143),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_179),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_147),
.A2(n_128),
.B(n_124),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_172),
.B(n_154),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_181),
.B(n_192),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_158),
.B1(n_133),
.B2(n_140),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_182),
.A2(n_188),
.B1(n_175),
.B2(n_160),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_160),
.A2(n_153),
.B1(n_152),
.B2(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_190),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_177),
.A2(n_156),
.B1(n_137),
.B2(n_148),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_176),
.B(n_141),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g194 ( 
.A1(n_162),
.A2(n_128),
.B(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_194),
.B(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_175),
.B(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_146),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_160),
.C(n_168),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_190),
.C(n_183),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_207),
.B1(n_208),
.B2(n_188),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_203),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_162),
.B1(n_163),
.B2(n_167),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_180),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

AOI221xp5_ASAP7_75t_L g210 ( 
.A1(n_196),
.A2(n_163),
.B1(n_167),
.B2(n_166),
.C(n_161),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g218 ( 
.A(n_210),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_213),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_187),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_197),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_216),
.B(n_208),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_182),
.B1(n_165),
.B2(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_200),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_221),
.B(n_226),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_209),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_223),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_202),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_191),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_202),
.B1(n_219),
.B2(n_204),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_SL g235 ( 
.A1(n_228),
.A2(n_230),
.B(n_231),
.Y(n_235)
);

OAI321xp33_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_227),
.A3(n_225),
.B1(n_207),
.B2(n_193),
.C(n_222),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_205),
.B1(n_199),
.B2(n_165),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_233),
.B(n_234),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_SL g233 ( 
.A1(n_227),
.A2(n_178),
.B(n_189),
.C(n_223),
.Y(n_233)
);

AOI322xp5_ASAP7_75t_L g234 ( 
.A1(n_231),
.A2(n_212),
.A3(n_159),
.B1(n_191),
.B2(n_171),
.C1(n_170),
.C2(n_164),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_179),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_237),
.B(n_146),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_236),
.B1(n_102),
.B2(n_169),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_239),
.A2(n_169),
.B(n_118),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_169),
.Y(n_241)
);


endmodule