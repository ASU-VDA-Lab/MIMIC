module fake_jpeg_10385_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_20),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_38),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_43),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_19),
.B1(n_31),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_45),
.A2(n_51),
.B1(n_57),
.B2(n_16),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_66),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_63),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_19),
.B1(n_31),
.B2(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_59),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_30),
.B1(n_18),
.B2(n_29),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_60),
.B1(n_16),
.B2(n_1),
.Y(n_82)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_62),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_34),
.A2(n_23),
.B1(n_17),
.B2(n_21),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_35),
.A2(n_30),
.B1(n_22),
.B2(n_23),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_28),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_21),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_77),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_88),
.Y(n_89)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_83),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_36),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_47),
.C(n_49),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_82),
.A2(n_46),
.B1(n_64),
.B2(n_50),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_43),
.B1(n_35),
.B2(n_4),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_50),
.B1(n_26),
.B2(n_55),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_14),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_86),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_0),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_92),
.B(n_70),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_48),
.B1(n_64),
.B2(n_63),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_93),
.A2(n_94),
.B1(n_111),
.B2(n_50),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_64),
.B1(n_46),
.B2(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_102),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_47),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_106),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_105),
.A2(n_69),
.B1(n_80),
.B2(n_6),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_36),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_40),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_40),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_76),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_40),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_43),
.B1(n_39),
.B2(n_58),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_103),
.B(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_123),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_74),
.B1(n_77),
.B2(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

A2O1A1O1Ixp25_ASAP7_75t_L g116 ( 
.A1(n_104),
.A2(n_76),
.B(n_72),
.C(n_85),
.D(n_86),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_101),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_118),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_102),
.B(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_126),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_127),
.A2(n_128),
.B(n_132),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_70),
.B(n_4),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_100),
.B(n_91),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_89),
.B(n_2),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_80),
.B1(n_5),
.B2(n_6),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_149),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_106),
.C(n_99),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_141),
.B(n_145),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_94),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_112),
.C(n_93),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_146),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_101),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_109),
.B(n_97),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_123),
.B(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_120),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_152),
.B1(n_98),
.B2(n_96),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_119),
.B1(n_91),
.B2(n_132),
.Y(n_158)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_148),
.A2(n_126),
.B(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_165),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_167),
.B(n_2),
.Y(n_181)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_160),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_139),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_161),
.B(n_5),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_147),
.A2(n_117),
.B1(n_115),
.B2(n_113),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_162),
.A2(n_163),
.B1(n_171),
.B2(n_98),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_147),
.A2(n_133),
.B1(n_116),
.B2(n_130),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_166),
.B1(n_154),
.B2(n_136),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_156),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_140),
.B1(n_139),
.B2(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_175),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_155),
.B1(n_143),
.B2(n_154),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_169),
.B(n_138),
.C(n_146),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_179),
.C(n_184),
.Y(n_197)
);

AOI221xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_181),
.B1(n_183),
.B2(n_187),
.C(n_167),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_92),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_186),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_166),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_165),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_191),
.B(n_159),
.Y(n_201)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_193),
.Y(n_208)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_194),
.B(n_183),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_174),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_199),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_171),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_160),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_185),
.B(n_178),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_189),
.A2(n_157),
.B1(n_170),
.B2(n_175),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_202),
.A2(n_168),
.B1(n_96),
.B2(n_8),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_186),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_204),
.B(n_192),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_205),
.B(n_211),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_184),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_197),
.C(n_199),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_13),
.Y(n_218)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_200),
.B(n_203),
.C(n_202),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_204),
.B1(n_208),
.B2(n_206),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_210),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_197),
.Y(n_214)
);

OAI21x1_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_215),
.B(n_212),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_6),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_220),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_222),
.A2(n_223),
.B(n_217),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_7),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_216),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_226),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_213),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_227),
.A2(n_220),
.B(n_8),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_228),
.A3(n_229),
.B1(n_9),
.B2(n_11),
.C1(n_7),
.C2(n_13),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_8),
.B(n_9),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_232),
.A2(n_9),
.B(n_12),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_12),
.Y(n_234)
);


endmodule