module fake_jpeg_10593_n_62 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx2_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_36),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_6),
.B(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_11),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_25),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_41),
.Y(n_54)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_37),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_49),
.Y(n_52)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_20),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_47),
.B1(n_43),
.B2(n_40),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_52),
.Y(n_58)
);

MAJx2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_54),
.C(n_55),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_59),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_50),
.C(n_51),
.Y(n_61)
);

MAJx2_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_50),
.C(n_53),
.Y(n_62)
);


endmodule