module fake_jpeg_2800_n_230 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

BUFx16f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_13),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_82),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_68),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_85),
.A2(n_61),
.B1(n_64),
.B2(n_78),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_92),
.B1(n_83),
.B2(n_67),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_64),
.B1(n_77),
.B2(n_62),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_97),
.B(n_100),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_65),
.B1(n_77),
.B2(n_70),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_99),
.A2(n_65),
.B1(n_87),
.B2(n_86),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_60),
.Y(n_100)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_105),
.B1(n_96),
.B2(n_67),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_70),
.B1(n_62),
.B2(n_76),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_66),
.B1(n_59),
.B2(n_74),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_58),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_57),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_98),
.B(n_57),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_109),
.B(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_113),
.Y(n_122)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_118),
.Y(n_134)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_119),
.Y(n_129)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_94),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_59),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_106),
.A2(n_72),
.B1(n_63),
.B2(n_56),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_131),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_151)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_137),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_83),
.B1(n_94),
.B2(n_75),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_141),
.B1(n_142),
.B2(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_50),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_9),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_75),
.B1(n_71),
.B2(n_55),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_138),
.A2(n_102),
.B1(n_114),
.B2(n_107),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_71),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.C(n_0),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_55),
.C(n_73),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_73),
.B1(n_53),
.B2(n_2),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_73),
.B(n_53),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_5),
.B(n_6),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_111),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_144),
.B(n_162),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_158),
.B1(n_136),
.B2(n_122),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_166),
.Y(n_186)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_37),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_123),
.A2(n_116),
.B1(n_3),
.B2(n_4),
.Y(n_149)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_159),
.B(n_165),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_151),
.B(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_1),
.B(n_5),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_155),
.A2(n_14),
.B(n_16),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_141),
.B(n_132),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_49),
.B1(n_47),
.B2(n_44),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_10),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_125),
.A2(n_10),
.B(n_11),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_126),
.B(n_15),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_133),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_12),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_167),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_181),
.B1(n_182),
.B2(n_165),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_130),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_190),
.C(n_158),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_189),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_179),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_177),
.B(n_164),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_26),
.B1(n_39),
.B2(n_36),
.Y(n_181)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_145),
.A2(n_168),
.B(n_156),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_163),
.A2(n_41),
.B(n_35),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_184),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_14),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_148),
.B(n_33),
.C(n_31),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_199),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_184),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_182),
.A2(n_149),
.B1(n_159),
.B2(n_155),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_198),
.B1(n_200),
.B2(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_187),
.C(n_172),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_169),
.C(n_188),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_197),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_151),
.B1(n_19),
.B2(n_20),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_17),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_193),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_19),
.B1(n_23),
.B2(n_24),
.Y(n_203)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_210),
.C(n_191),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_195),
.Y(n_208)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_169),
.C(n_190),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_186),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_175),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_211),
.A2(n_194),
.B1(n_176),
.B2(n_199),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_175),
.B1(n_205),
.B2(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_214),
.B(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_216),
.B(n_218),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_217),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_221),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_224),
.A2(n_220),
.B(n_210),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_225),
.A2(n_209),
.B(n_216),
.Y(n_226)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_215),
.CI(n_204),
.CON(n_227),
.SN(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_181),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_228),
.A2(n_227),
.B(n_29),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_23),
.Y(n_230)
);


endmodule