module fake_jpeg_26091_n_35 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

AOI22xp33_ASAP7_75t_SL g8 ( 
.A1(n_6),
.A2(n_4),
.B1(n_0),
.B2(n_2),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_13),
.A2(n_16),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_2),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_9),
.B(n_3),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_23),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_17),
.C(n_16),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_25),
.B(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

MAJx2_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_16),
.C(n_8),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_3),
.Y(n_31)
);

AOI31xp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_30),
.A3(n_29),
.B(n_15),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_27),
.A2(n_5),
.B(n_11),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_5),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_34),
.B(n_32),
.Y(n_35)
);


endmodule