module fake_jpeg_5703_n_50 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_50);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_50;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx5_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx6_ASAP7_75t_SL g8 ( 
.A(n_1),
.Y(n_8)
);

INVx11_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx6_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_0),
.B(n_6),
.C(n_8),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_0),
.C(n_6),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_12),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

AND2x6_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_15),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_31),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_15),
.B(n_10),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_33),
.B(n_31),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_19),
.A2(n_9),
.B1(n_12),
.B2(n_22),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_29),
.B1(n_32),
.B2(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_40),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_40),
.C(n_39),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_43),
.B(n_37),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

AOI211xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_44),
.B(n_48),
.C(n_45),
.Y(n_50)
);


endmodule