module fake_aes_1007_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NAND2xp5_ASAP7_75t_L g13 ( .A(n_5), .B(n_9), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_12), .Y(n_14) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_6), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
BUFx6f_ASAP7_75t_L g19 ( .A(n_1), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_17), .B(n_0), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_15), .B(n_0), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
OAI221xp5_ASAP7_75t_SL g24 ( .A1(n_23), .A2(n_20), .B1(n_21), .B2(n_13), .C(n_19), .Y(n_24) );
AOI211x1_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_1), .B(n_2), .C(n_19), .Y(n_25) );
AOI211x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_2), .B(n_16), .C(n_14), .Y(n_26) );
XNOR2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_3), .Y(n_27) );
OAI22x1_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_18), .B1(n_7), .B2(n_8), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
endmodule