module fake_jpeg_23307_n_335 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_335);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_335;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_24),
.Y(n_61)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_41),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_17),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_48),
.B(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_18),
.B1(n_26),
.B2(n_23),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_52),
.A2(n_56),
.B1(n_72),
.B2(n_74),
.Y(n_93)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_53),
.B(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_34),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_61),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_34),
.Y(n_66)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_30),
.B1(n_20),
.B2(n_17),
.Y(n_112)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_31),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_73),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_36),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_31),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_27),
.B1(n_32),
.B2(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_25),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_91),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_52),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_80),
.A2(n_105),
.B1(n_54),
.B2(n_20),
.Y(n_121)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_82),
.Y(n_140)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_49),
.B1(n_66),
.B2(n_62),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_83),
.A2(n_86),
.B1(n_101),
.B2(n_10),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_19),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_84),
.B(n_95),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_19),
.B1(n_29),
.B2(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_87),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_25),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_44),
.C(n_43),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_17),
.C(n_28),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_44),
.Y(n_95)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_66),
.A2(n_29),
.B1(n_35),
.B2(n_30),
.Y(n_101)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_40),
.B1(n_72),
.B2(n_51),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_57),
.B(n_74),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_110),
.Y(n_128)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_112),
.A2(n_63),
.B1(n_64),
.B2(n_54),
.Y(n_116)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_113),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_114),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_123),
.B1(n_127),
.B2(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_137),
.C(n_78),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_28),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_92),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_76),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_142),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_94),
.B(n_5),
.C(n_6),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_91),
.A2(n_5),
.B(n_6),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_8),
.B(n_11),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_76),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_80),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_102),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_97),
.Y(n_154)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_147),
.B(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_115),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_152),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_SL g204 ( 
.A(n_149),
.B(n_159),
.C(n_171),
.Y(n_204)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_157),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_77),
.B(n_95),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_151),
.A2(n_153),
.B(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_89),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_89),
.B(n_112),
.Y(n_153)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_138),
.A2(n_127),
.B(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_156),
.Y(n_211)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_115),
.B(n_89),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_128),
.A2(n_93),
.B(n_79),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_85),
.Y(n_161)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_121),
.A2(n_111),
.B(n_113),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_164),
.A2(n_168),
.B(n_173),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_142),
.B(n_90),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_136),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_167),
.B(n_172),
.Y(n_205)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_122),
.B(n_81),
.Y(n_168)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_96),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_131),
.A2(n_114),
.B(n_88),
.C(n_107),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_100),
.B(n_99),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_103),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_177),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_134),
.Y(n_176)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_12),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_180),
.B(n_200),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_125),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_185),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_126),
.C(n_125),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_203),
.C(n_206),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_172),
.A2(n_98),
.B1(n_135),
.B2(n_126),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_210),
.B1(n_165),
.B2(n_163),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_146),
.A2(n_130),
.B1(n_133),
.B2(n_124),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_157),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_146),
.A2(n_130),
.B1(n_133),
.B2(n_124),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_120),
.B1(n_117),
.B2(n_87),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_196),
.Y(n_222)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_198),
.A2(n_178),
.B(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_82),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_168),
.B(n_120),
.C(n_129),
.Y(n_206)
);

A2O1A1Ixp33_ASAP7_75t_SL g207 ( 
.A1(n_164),
.A2(n_104),
.B(n_106),
.C(n_14),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_207),
.A2(n_151),
.B(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_209),
.B(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_159),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_209),
.A2(n_174),
.B1(n_177),
.B2(n_166),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_212),
.A2(n_214),
.B1(n_227),
.B2(n_232),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_233),
.B1(n_234),
.B2(n_182),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_204),
.A2(n_166),
.B1(n_145),
.B2(n_171),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_224),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_216),
.A2(n_220),
.B(n_221),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_150),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_204),
.B(n_145),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_237),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_158),
.Y(n_223)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_189),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_226),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_188),
.A2(n_149),
.B1(n_168),
.B2(n_147),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_155),
.Y(n_228)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_228),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_208),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_236),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_176),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_188),
.A2(n_168),
.B1(n_173),
.B2(n_155),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_205),
.A2(n_193),
.B1(n_206),
.B2(n_210),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_235),
.A2(n_198),
.B(n_199),
.Y(n_244)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_192),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_162),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_162),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_239),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_202),
.B(n_193),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_240),
.A2(n_221),
.B1(n_213),
.B2(n_225),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_241),
.A2(n_214),
.B1(n_212),
.B2(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_184),
.C(n_202),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_243),
.C(n_234),
.Y(n_274)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_182),
.B(n_196),
.C(n_207),
.D(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_244),
.B(n_251),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_249),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_233),
.B(n_207),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_254),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_218),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_256),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_228),
.A2(n_207),
.B(n_211),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

INVx13_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_255),
.B(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_267),
.Y(n_290)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_218),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_271),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_223),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_247),
.B(n_237),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_280),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_222),
.C(n_230),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_243),
.C(n_240),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_279),
.B1(n_252),
.B2(n_222),
.Y(n_284)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_257),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_288),
.C(n_270),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_284),
.A2(n_281),
.B1(n_263),
.B2(n_267),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_249),
.B(n_253),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_286),
.A2(n_245),
.B(n_195),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_247),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_291),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_249),
.A3(n_232),
.B1(n_244),
.B2(n_259),
.C1(n_254),
.C2(n_256),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_275),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_278),
.A2(n_259),
.B1(n_245),
.B2(n_246),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_296),
.A2(n_279),
.B1(n_271),
.B2(n_272),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_304),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_302),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_283),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_301),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_277),
.C(n_265),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_295),
.A2(n_281),
.B(n_266),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_307),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_308),
.B1(n_284),
.B2(n_290),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_270),
.C(n_274),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_289),
.A2(n_262),
.B(n_194),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_289),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_298),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_194),
.B1(n_276),
.B2(n_282),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_294),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_316),
.B(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_276),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_314),
.A2(n_285),
.A3(n_276),
.B1(n_303),
.B2(n_307),
.C1(n_304),
.C2(n_306),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_323),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_282),
.B1(n_179),
.B2(n_288),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_324),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_235),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g324 ( 
.A1(n_314),
.A2(n_197),
.A3(n_179),
.B1(n_157),
.B2(n_169),
.C1(n_15),
.C2(n_12),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_325),
.B(n_316),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_329),
.B(n_328),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_312),
.B(n_320),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_331),
.C(n_327),
.Y(n_332)
);

OAI21x1_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_328),
.B(n_323),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_169),
.CI(n_15),
.CON(n_334),
.SN(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_308),
.Y(n_335)
);


endmodule