module real_jpeg_6418_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_0),
.Y(n_132)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_0),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_1),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_1),
.B(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_4),
.B(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_4),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_4),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_4),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_4),
.B(n_328),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_4),
.B(n_98),
.Y(n_359)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_6),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_6),
.Y(n_211)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_6),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g301 ( 
.A(n_6),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_7),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_7),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_7),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_7),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_7),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_7),
.B(n_241),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_7),
.B(n_262),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_8),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_8),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_8),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_8),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_9),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_9),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_9),
.B(n_163),
.Y(n_162)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_9),
.B(n_51),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_9),
.B(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_9),
.B(n_33),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_10),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_10),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_10),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_10),
.B(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_10),
.B(n_284),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_10),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_10),
.B(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_11),
.Y(n_113)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_11),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_12),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_12),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_12),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_12),
.B(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_12),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_12),
.B(n_185),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_12),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_12),
.B(n_308),
.Y(n_358)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_14),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_15),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_15),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_15),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_15),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_15),
.B(n_56),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_15),
.B(n_244),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_16),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_16),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_16),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_16),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_16),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_16),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_16),
.B(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_17),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_17),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_17),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_17),
.Y(n_322)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_191),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_190),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_148),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_23),
.B(n_148),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g438 ( 
.A(n_23),
.Y(n_438)
);

FAx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_91),
.CI(n_125),
.CON(n_23),
.SN(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_63),
.C(n_76),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_25),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_40),
.C(n_49),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_26),
.B(n_201),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_35),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_28),
.B(n_32),
.C(n_35),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_28),
.A2(n_29),
.B1(n_45),
.B2(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_41),
.C(n_45),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_31),
.A2(n_32),
.B1(n_97),
.B2(n_101),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_32),
.B(n_97),
.C(n_106),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_37),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_39),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_40),
.B(n_49),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_41),
.B(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_46),
.Y(n_181)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_48),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_48),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_55),
.C(n_58),
.Y(n_145)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_52),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_56),
.Y(n_137)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_57),
.Y(n_167)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g305 ( 
.A(n_60),
.Y(n_305)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_61),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_61),
.Y(n_361)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_63),
.B(n_76),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_64),
.B(n_70),
.C(n_75),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_70),
.A2(n_71),
.B1(n_88),
.B2(n_89),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_77),
.C(n_88),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_73),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_73),
.Y(n_340)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_74),
.Y(n_214)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_74),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_78),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.C(n_85),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_79),
.B(n_85),
.Y(n_156)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_83),
.B(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_84),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_84),
.Y(n_292)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_104),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_102),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_101),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_100),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_106),
.B(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_119),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_113),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_119),
.Y(n_147)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_124),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_142),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

INVx8_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_141),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_146),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_151),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_153),
.B(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_171),
.C(n_173),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_168),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_155),
.B(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_157),
.A2(n_158),
.B1(n_168),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_165),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_159),
.B(n_165),
.Y(n_410)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_162),
.B(n_410),
.Y(n_409)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_168),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_173),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_184),
.C(n_186),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_174),
.B(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.C(n_182),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_207),
.Y(n_206)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_179),
.B(n_182),
.Y(n_207)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_186),
.Y(n_229)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_247),
.B(n_435),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_193),
.B(n_195),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.C(n_202),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_197),
.B(n_200),
.Y(n_430)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_202),
.B(n_430),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_227),
.C(n_230),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_204),
.B(n_423),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.C(n_215),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_205),
.A2(n_206),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_208),
.A2(n_209),
.B(n_212),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_208),
.B(n_215),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.C(n_224),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_378)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_223),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_224),
.B(n_378),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_225),
.B(n_321),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_230),
.Y(n_424)
);

MAJx2_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_240),
.C(n_243),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_232),
.B(n_412),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_233),
.B(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_236),
.Y(n_391)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_240),
.B(n_243),
.Y(n_412)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI21x1_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_428),
.B(n_434),
.Y(n_247)
);

OAI21x1_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_415),
.B(n_427),
.Y(n_248)
);

AOI21x1_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_397),
.B(n_414),
.Y(n_249)
);

OAI21x1_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_371),
.B(n_396),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_345),
.B(n_370),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_313),
.B(n_344),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_294),
.B(n_312),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_275),
.B(n_293),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_269),
.B(n_274),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_265),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_261),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_261),
.Y(n_276)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx8_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_264),
.Y(n_273)
);

INVx4_ASAP7_75t_L g325 ( 
.A(n_264),
.Y(n_325)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_277),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_285),
.B2(n_286),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_278),
.B(n_288),
.C(n_290),
.Y(n_311)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_280),
.B(n_283),
.Y(n_302)
);

INVx8_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_311),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_311),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_303),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_302),
.C(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_300),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_303),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_304),
.B(n_333),
.C(n_334),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_310),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_310),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_316),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_316),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_331),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_317),
.B(n_332),
.C(n_335),
.Y(n_369)
);

XOR2x2_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_320),
.C(n_323),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

INVx4_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_326),
.B1(n_327),
.B2(n_330),
.Y(n_323)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_324),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_336),
.B(n_341),
.C(n_342),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_341),
.B1(n_342),
.B2(n_343),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_339),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_341),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_346),
.B(n_369),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_369),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_356),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_355),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_348),
.B(n_355),
.C(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_354),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_354),
.B(n_385),
.C(n_386),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_362),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_364),
.C(n_367),
.Y(n_374)
);

BUFx24_ASAP7_75t_SL g436 ( 
.A(n_357),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_359),
.CI(n_360),
.CON(n_357),
.SN(n_357)
);

MAJx2_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_359),
.C(n_360),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_364),
.B1(n_367),
.B2(n_368),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_365),
.B(n_366),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_368),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_394),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_394),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_383),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_374),
.B(n_375),
.C(n_383),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_379),
.B2(n_380),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_406),
.C(n_407),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_382),
.Y(n_380)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_381),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_382),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_384),
.B(n_388),
.C(n_393),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_392),
.B2(n_393),
.Y(n_387)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_388),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_413),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_413),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_403),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_403),
.C(n_426),
.Y(n_425)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_404),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_408),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_409),
.C(n_411),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_425),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_425),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.Y(n_416)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_417),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_432),
.C(n_433),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_422),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_431),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_431),
.Y(n_434)
);


endmodule