module fake_netlist_6_360_n_9051 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_98, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_54, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_100, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_108, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_103, n_111, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_9051);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_54;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_100;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_108;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_9051;

wire n_5643;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_6566;
wire n_2576;
wire n_5172;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_6872;
wire n_1351;
wire n_5254;
wire n_6441;
wire n_8668;
wire n_1212;
wire n_208;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_5019;
wire n_2332;
wire n_8713;
wire n_7111;
wire n_6141;
wire n_3849;
wire n_7933;
wire n_7967;
wire n_578;
wire n_5138;
wire n_4388;
wire n_4395;
wire n_6960;
wire n_1061;
wire n_3089;
wire n_8169;
wire n_9002;
wire n_783;
wire n_7180;
wire n_5653;
wire n_4978;
wire n_8604;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_188;
wire n_1854;
wire n_3088;
wire n_8168;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_7190;
wire n_1387;
wire n_3222;
wire n_7504;
wire n_8186;
wire n_677;
wire n_6126;
wire n_6725;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_8899;
wire n_2317;
wire n_5524;
wire n_442;
wire n_5345;
wire n_8023;
wire n_1975;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_8130;
wire n_2179;
wire n_8534;
wire n_5963;
wire n_5055;
wire n_1547;
wire n_3376;
wire n_4868;
wire n_893;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_4249;
wire n_5950;
wire n_1192;
wire n_3564;
wire n_1844;
wire n_6999;
wire n_1555;
wire n_5548;
wire n_5057;
wire n_8339;
wire n_8272;
wire n_7161;
wire n_3030;
wire n_830;
wire n_7868;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_447;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_3427;
wire n_852;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_7000;
wire n_8561;
wire n_7398;
wire n_2926;
wire n_1078;
wire n_544;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_8411;
wire n_2321;
wire n_8499;
wire n_2019;
wire n_8236;
wire n_5102;
wire n_3345;
wire n_2074;
wire n_6882;
wire n_2919;
wire n_4501;
wire n_2129;
wire n_6325;
wire n_4724;
wire n_945;
wire n_5598;
wire n_7983;
wire n_7389;
wire n_4997;
wire n_2399;
wire n_9018;
wire n_4843;
wire n_1232;
wire n_8070;
wire n_4696;
wire n_6660;
wire n_4347;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_3877;
wire n_3929;
wire n_8366;
wire n_3048;
wire n_1455;
wire n_8102;
wire n_7401;
wire n_7516;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_8175;
wire n_8977;
wire n_5239;
wire n_567;
wire n_1781;
wire n_1971;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_5332;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_5908;
wire n_3077;
wire n_2873;
wire n_3452;
wire n_8913;
wire n_3107;
wire n_155;
wire n_4956;
wire n_454;
wire n_7686;
wire n_1421;
wire n_3664;
wire n_6914;
wire n_1936;
wire n_5337;
wire n_5129;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_6585;
wire n_713;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_6374;
wire n_2843;
wire n_7651;
wire n_6628;
wire n_8125;
wire n_3760;
wire n_6015;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_6526;
wire n_1894;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_8556;
wire n_7196;
wire n_3347;
wire n_5136;
wire n_907;
wire n_8040;
wire n_5638;
wire n_4110;
wire n_6784;
wire n_1658;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_6323;
wire n_6110;
wire n_1967;
wire n_3999;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_7846;
wire n_8595;
wire n_2708;
wire n_1648;
wire n_5151;
wire n_1911;
wire n_8142;
wire n_2011;
wire n_5684;
wire n_8598;
wire n_5729;
wire n_7256;
wire n_281;
wire n_6404;
wire n_7331;
wire n_7774;
wire n_7856;
wire n_564;
wire n_5680;
wire n_6674;
wire n_6951;
wire n_6148;
wire n_7625;
wire n_279;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_2735;
wire n_4662;
wire n_8869;
wire n_6989;
wire n_4671;
wire n_7863;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_4314;
wire n_2080;
wire n_8958;
wire n_323;
wire n_5099;
wire n_6896;
wire n_7770;
wire n_8421;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_1381;
wire n_331;
wire n_1699;
wire n_2093;
wire n_4296;
wire n_7147;
wire n_2770;
wire n_8115;
wire n_608;
wire n_2101;
wire n_4507;
wire n_8389;
wire n_5902;
wire n_512;
wire n_3484;
wire n_4677;
wire n_792;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_1328;
wire n_2917;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_3923;
wire n_9042;
wire n_3900;
wire n_8412;
wire n_3488;
wire n_939;
wire n_3732;
wire n_2811;
wire n_6485;
wire n_8987;
wire n_6107;
wire n_2832;
wire n_4226;
wire n_8849;
wire n_1762;
wire n_5493;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_237;
wire n_6863;
wire n_6282;
wire n_6994;
wire n_1895;
wire n_4294;
wire n_4698;
wire n_4445;
wire n_4810;
wire n_7564;
wire n_3859;
wire n_2692;
wire n_175;
wire n_6768;
wire n_6383;
wire n_7234;
wire n_3914;
wire n_4456;
wire n_8119;
wire n_3397;
wire n_8641;
wire n_3575;
wire n_8151;
wire n_8118;
wire n_2469;
wire n_9038;
wire n_8748;
wire n_3927;
wire n_8436;
wire n_5452;
wire n_6794;
wire n_3888;
wire n_6151;
wire n_8718;
wire n_7110;
wire n_764;
wire n_5476;
wire n_2764;
wire n_2895;
wire n_6431;
wire n_6990;
wire n_8659;
wire n_733;
wire n_2922;
wire n_8223;
wire n_3882;
wire n_4856;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_7849;
wire n_8915;
wire n_4331;
wire n_7297;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_7298;
wire n_5536;
wire n_2072;
wire n_1354;
wire n_7533;
wire n_586;
wire n_423;
wire n_7221;
wire n_4375;
wire n_1701;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_2678;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_8246;
wire n_5897;
wire n_1726;
wire n_5532;
wire n_4613;
wire n_8952;
wire n_2434;
wire n_2878;
wire n_3012;
wire n_3875;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_4877;
wire n_3247;
wire n_871;
wire n_5922;
wire n_210;
wire n_7569;
wire n_2641;
wire n_7734;
wire n_7823;
wire n_7861;
wire n_7062;
wire n_8955;
wire n_5658;
wire n_4731;
wire n_3052;
wire n_178;
wire n_7039;
wire n_355;
wire n_8577;
wire n_8594;
wire n_5046;
wire n_8428;
wire n_2749;
wire n_3298;
wire n_8848;
wire n_2254;
wire n_5058;
wire n_1926;
wire n_3273;
wire n_4467;
wire n_7077;
wire n_1747;
wire n_195;
wire n_5667;
wire n_780;
wire n_8259;
wire n_2624;
wire n_5865;
wire n_8349;
wire n_6836;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_4681;
wire n_8164;
wire n_4072;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_7905;
wire n_8776;
wire n_8287;
wire n_2092;
wire n_7753;
wire n_1654;
wire n_6771;
wire n_7950;
wire n_1750;
wire n_1462;
wire n_8607;
wire n_2514;
wire n_604;
wire n_6248;
wire n_6952;
wire n_6795;
wire n_5314;
wire n_1588;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_2468;
wire n_4381;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_515;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_8066;
wire n_6831;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_5795;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_5226;
wire n_6715;
wire n_514;
wire n_6714;
wire n_687;
wire n_890;
wire n_7677;
wire n_5457;
wire n_8416;
wire n_2812;
wire n_190;
wire n_4518;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_1709;
wire n_7009;
wire n_8453;
wire n_2393;
wire n_2657;
wire n_7149;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_8949;
wire n_3500;
wire n_3834;
wire n_4589;
wire n_2075;
wire n_2972;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_2763;
wire n_2762;
wire n_3192;
wire n_8995;
wire n_760;
wire n_1546;
wire n_4394;
wire n_6581;
wire n_2279;
wire n_161;
wire n_6010;
wire n_1296;
wire n_3352;
wire n_8711;
wire n_3073;
wire n_7013;
wire n_5343;
wire n_2150;
wire n_1294;
wire n_4082;
wire n_1420;
wire n_3696;
wire n_7290;
wire n_595;
wire n_1779;
wire n_524;
wire n_4921;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_8306;
wire n_7488;
wire n_2558;
wire n_7315;
wire n_8887;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_3763;
wire n_6185;
wire n_2712;
wire n_5529;
wire n_3733;
wire n_7889;
wire n_6042;
wire n_1487;
wire n_3614;
wire n_874;
wire n_382;
wire n_5183;
wire n_8500;
wire n_7438;
wire n_2145;
wire n_7268;
wire n_7337;
wire n_898;
wire n_4964;
wire n_5957;
wire n_6965;
wire n_4228;
wire n_3423;
wire n_6357;
wire n_925;
wire n_1932;
wire n_1101;
wire n_6800;
wire n_4636;
wire n_7461;
wire n_8285;
wire n_4322;
wire n_3644;
wire n_6955;
wire n_8483;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_8332;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_2767;
wire n_7278;
wire n_6509;
wire n_4576;
wire n_7454;
wire n_5929;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_1521;
wire n_8741;
wire n_1366;
wire n_4000;
wire n_5445;
wire n_2897;
wire n_4389;
wire n_3970;
wire n_5501;
wire n_6839;
wire n_7232;
wire n_7377;
wire n_4345;
wire n_5342;
wire n_996;
wire n_532;
wire n_173;
wire n_6646;
wire n_8648;
wire n_1376;
wire n_413;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_7098;
wire n_7069;
wire n_7904;
wire n_6033;
wire n_977;
wire n_536;
wire n_3158;
wire n_1788;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_1835;
wire n_8394;
wire n_3470;
wire n_5076;
wire n_581;
wire n_5870;
wire n_4713;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_432;
wire n_3700;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_3104;
wire n_6809;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_7840;
wire n_4310;
wire n_6359;
wire n_7782;
wire n_1432;
wire n_5212;
wire n_989;
wire n_8800;
wire n_7080;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_2191;
wire n_8229;
wire n_1246;
wire n_4528;
wire n_8410;
wire n_5811;
wire n_899;
wire n_7739;
wire n_7624;
wire n_1035;
wire n_4914;
wire n_6766;
wire n_4939;
wire n_7629;
wire n_499;
wire n_1426;
wire n_3418;
wire n_705;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_4634;
wire n_2069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_7003;
wire n_3119;
wire n_5427;
wire n_3735;
wire n_2297;
wire n_4379;
wire n_486;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_1448;
wire n_5901;
wire n_6538;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_7010;
wire n_648;
wire n_8107;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_6519;
wire n_2103;
wire n_8983;
wire n_3770;
wire n_2772;
wire n_6530;
wire n_7219;
wire n_4440;
wire n_8774;
wire n_4402;
wire n_927;
wire n_5052;
wire n_7299;
wire n_4541;
wire n_5009;
wire n_4872;
wire n_929;
wire n_6402;
wire n_4551;
wire n_2857;
wire n_6195;
wire n_7243;
wire n_6609;
wire n_7326;
wire n_7471;
wire n_5326;
wire n_7067;
wire n_1183;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_8620;
wire n_8691;
wire n_3342;
wire n_6748;
wire n_7741;
wire n_998;
wire n_5035;
wire n_717;
wire n_7790;
wire n_6149;
wire n_1383;
wire n_7484;
wire n_3390;
wire n_3656;
wire n_7002;
wire n_1424;
wire n_6414;
wire n_1000;
wire n_8424;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_7528;
wire n_8026;
wire n_3810;
wire n_552;
wire n_4798;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_216;
wire n_8174;
wire n_7941;
wire n_912;
wire n_5010;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_5089;
wire n_2849;
wire n_1398;
wire n_1201;
wire n_884;
wire n_5394;
wire n_4592;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_2661;
wire n_8861;
wire n_731;
wire n_5359;
wire n_8644;
wire n_1955;
wire n_8907;
wire n_931;
wire n_474;
wire n_312;
wire n_1791;
wire n_958;
wire n_5137;
wire n_6902;
wire n_3331;
wire n_5104;
wire n_1897;
wire n_2064;
wire n_7117;
wire n_5741;
wire n_8324;
wire n_2773;
wire n_6205;
wire n_6380;
wire n_7478;
wire n_7913;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_589;
wire n_3606;
wire n_1310;
wire n_819;
wire n_1334;
wire n_3591;
wire n_7939;
wire n_2788;
wire n_964;
wire n_8503;
wire n_4756;
wire n_8196;
wire n_6449;
wire n_2797;
wire n_7458;
wire n_6723;
wire n_6440;
wire n_7436;
wire n_4746;
wire n_124;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_211;
wire n_2748;
wire n_8446;
wire n_5194;
wire n_1834;
wire n_9033;
wire n_2331;
wire n_2292;
wire n_7435;
wire n_3441;
wire n_3534;
wire n_6997;
wire n_5952;
wire n_3964;
wire n_2416;
wire n_311;
wire n_5947;
wire n_8923;
wire n_1877;
wire n_3944;
wire n_6124;
wire n_7685;
wire n_6736;
wire n_7363;
wire n_8192;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_5985;
wire n_8197;
wire n_556;
wire n_2209;
wire n_3605;
wire n_6622;
wire n_1602;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_3306;
wire n_276;
wire n_3026;
wire n_221;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_8082;
wire n_4428;
wire n_8730;
wire n_1533;
wire n_3323;
wire n_7917;
wire n_7261;
wire n_266;
wire n_9023;
wire n_6528;
wire n_2274;
wire n_7532;
wire n_8051;
wire n_5761;
wire n_518;
wire n_6773;
wire n_4618;
wire n_7375;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_317;
wire n_4805;
wire n_1679;
wire n_8651;
wire n_3454;
wire n_2160;
wire n_5760;
wire n_6885;
wire n_2146;
wire n_6531;
wire n_2131;
wire n_488;
wire n_7430;
wire n_5472;
wire n_3547;
wire n_8377;
wire n_5679;
wire n_7912;
wire n_2575;
wire n_5100;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_7728;
wire n_4410;
wire n_1933;
wire n_8281;
wire n_1179;
wire n_324;
wire n_3816;
wire n_4807;
wire n_8842;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_301;
wire n_2928;
wire n_5166;
wire n_9046;
wire n_6339;
wire n_1917;
wire n_8024;
wire n_1580;
wire n_7730;
wire n_8814;
wire n_8530;
wire n_2822;
wire n_4180;
wire n_1281;
wire n_8467;
wire n_7281;
wire n_3109;
wire n_3354;
wire n_2572;
wire n_7711;
wire n_1520;
wire n_3126;
wire n_8984;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_6417;
wire n_351;
wire n_5740;
wire n_259;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1832;
wire n_1645;
wire n_4676;
wire n_5180;
wire n_6763;
wire n_8956;
wire n_858;
wire n_2049;
wire n_5182;
wire n_7858;
wire n_8676;
wire n_956;
wire n_5534;
wire n_8003;
wire n_663;
wire n_4880;
wire n_8785;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_2781;
wire n_4126;
wire n_410;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_6556;
wire n_1594;
wire n_8692;
wire n_664;
wire n_1869;
wire n_6889;
wire n_7230;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_5196;
wire n_6199;
wire n_2016;
wire n_5171;
wire n_4470;
wire n_6726;
wire n_580;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_7011;
wire n_465;
wire n_8998;
wire n_1790;
wire n_5261;
wire n_4014;
wire n_4704;
wire n_341;
wire n_1744;
wire n_828;
wire n_2142;
wire n_4252;
wire n_607;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_2448;
wire n_8906;
wire n_5949;
wire n_4048;
wire n_4596;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_3406;
wire n_820;
wire n_951;
wire n_6100;
wire n_6516;
wire n_952;
wire n_3919;
wire n_8462;
wire n_6977;
wire n_7660;
wire n_6915;
wire n_2263;
wire n_7834;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_974;
wire n_6522;
wire n_8979;
wire n_5023;
wire n_2656;
wire n_4952;
wire n_2375;
wire n_5906;
wire n_1934;
wire n_8429;
wire n_8930;
wire n_628;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_7890;
wire n_3973;
wire n_2756;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_807;
wire n_4761;
wire n_6675;
wire n_6270;
wire n_1275;
wire n_2884;
wire n_6808;
wire n_485;
wire n_1510;
wire n_7620;
wire n_7265;
wire n_7986;
wire n_7006;
wire n_6931;
wire n_6207;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_6245;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_238;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_202;
wire n_1749;
wire n_3474;
wire n_6963;
wire n_8685;
wire n_2549;
wire n_4690;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_8264;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_5456;
wire n_248;
wire n_2302;
wire n_8135;
wire n_1667;
wire n_7837;
wire n_7717;
wire n_8445;
wire n_1037;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_3592;
wire n_468;
wire n_5500;
wire n_6412;
wire n_4230;
wire n_2637;
wire n_1639;
wire n_7627;
wire n_183;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_3195;
wire n_466;
wire n_2526;
wire n_6346;
wire n_4274;
wire n_7860;
wire n_5215;
wire n_8408;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_7335;
wire n_4189;
wire n_8895;
wire n_3817;
wire n_7811;
wire n_340;
wire n_1108;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_5003;
wire n_4827;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_8450;
wire n_3648;
wire n_8273;
wire n_1686;
wire n_6059;
wire n_7499;
wire n_3042;
wire n_6065;
wire n_7292;
wire n_5094;
wire n_4610;
wire n_4472;
wire n_7870;
wire n_5433;
wire n_9043;
wire n_6075;
wire n_3228;
wire n_3657;
wire n_7397;
wire n_3081;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_7211;
wire n_5618;
wire n_6861;
wire n_8312;
wire n_6781;
wire n_1586;
wire n_7847;
wire n_8506;
wire n_2264;
wire n_3464;
wire n_6494;
wire n_380;
wire n_6133;
wire n_3723;
wire n_1190;
wire n_8963;
wire n_7822;
wire n_397;
wire n_4380;
wire n_6453;
wire n_5978;
wire n_4990;
wire n_4996;
wire n_6127;
wire n_5247;
wire n_4398;
wire n_2498;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_6006;
wire n_2235;
wire n_7289;
wire n_4193;
wire n_3570;
wire n_7926;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_172;
wire n_7354;
wire n_8352;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_239;
wire n_7960;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_5689;
wire n_7482;
wire n_1043;
wire n_4090;
wire n_6115;
wire n_4165;
wire n_8143;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_352;
wire n_6838;
wire n_6867;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_6139;
wire n_1361;
wire n_662;
wire n_6256;
wire n_7965;
wire n_3262;
wire n_6613;
wire n_4008;
wire n_3356;
wire n_5221;
wire n_5641;
wire n_1642;
wire n_3210;
wire n_6361;
wire n_937;
wire n_4689;
wire n_8183;
wire n_1682;
wire n_4547;
wire n_6085;
wire n_7474;
wire n_5731;
wire n_6329;
wire n_8650;
wire n_6678;
wire n_3329;
wire n_8662;
wire n_330;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_1406;
wire n_4601;
wire n_962;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_8526;
wire n_1186;
wire n_4623;
wire n_7325;
wire n_5007;
wire n_7044;
wire n_3320;
wire n_6370;
wire n_8623;
wire n_2518;
wire n_5883;
wire n_7166;
wire n_6554;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_3988;
wire n_6560;
wire n_1720;
wire n_3476;
wire n_7838;
wire n_4842;
wire n_204;
wire n_482;
wire n_7028;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_7873;
wire n_2688;
wire n_394;
wire n_1845;
wire n_1489;
wire n_6535;
wire n_942;
wire n_7518;
wire n_2798;
wire n_7414;
wire n_6147;
wire n_2852;
wire n_1524;
wire n_8973;
wire n_6448;
wire n_7791;
wire n_1964;
wire n_8419;
wire n_1920;
wire n_2753;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_5934;
wire n_7431;
wire n_5434;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_1846;
wire n_3437;
wire n_4111;
wire n_6643;
wire n_533;
wire n_7146;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_2506;
wire n_6157;
wire n_4859;
wire n_2626;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_8351;
wire n_8430;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_8603;
wire n_5218;
wire n_8249;
wire n_7052;
wire n_3665;
wire n_273;
wire n_3007;
wire n_3528;
wire n_5960;
wire n_4571;
wire n_3698;
wire n_7888;
wire n_6397;
wire n_5358;
wire n_3355;
wire n_2454;
wire n_8234;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_1066;
wire n_1948;
wire n_157;
wire n_4215;
wire n_9010;
wire n_9003;
wire n_2154;
wire n_6073;
wire n_7502;
wire n_1484;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_7312;
wire n_7919;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_7085;
wire n_1373;
wire n_3958;
wire n_6939;
wire n_7848;
wire n_3985;
wire n_2427;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_6689;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_7580;
wire n_5149;
wire n_8980;
wire n_5571;
wire n_2680;
wire n_1047;
wire n_3375;
wire n_3899;
wire n_6698;
wire n_1385;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_502;
wire n_2668;
wire n_7288;
wire n_8558;
wire n_1257;
wire n_7707;
wire n_3197;
wire n_7223;
wire n_7833;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_7274;
wire n_9004;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_6206;
wire n_8136;
wire n_834;
wire n_5033;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_3124;
wire n_1741;
wire n_7466;
wire n_1002;
wire n_6529;
wire n_1949;
wire n_3759;
wire n_545;
wire n_2671;
wire n_4516;
wire n_6363;
wire n_6750;
wire n_2715;
wire n_1804;
wire n_8619;
wire n_251;
wire n_2508;
wire n_3511;
wire n_2054;
wire n_6290;
wire n_7429;
wire n_6025;
wire n_1337;
wire n_1477;
wire n_7277;
wire n_6455;
wire n_2614;
wire n_8146;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_5393;
wire n_8813;
wire n_5607;
wire n_3694;
wire n_7695;
wire n_2937;
wire n_7179;
wire n_7122;
wire n_7165;
wire n_7869;
wire n_4789;
wire n_5999;
wire n_8910;
wire n_4376;
wire n_6203;
wire n_1001;
wire n_6408;
wire n_2241;
wire n_6555;
wire n_7683;
wire n_6150;
wire n_7630;
wire n_4708;
wire n_8470;
wire n_4657;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_8643;
wire n_1076;
wire n_4512;
wire n_1378;
wire n_855;
wire n_1377;
wire n_8565;
wire n_695;
wire n_8550;
wire n_4081;
wire n_1542;
wire n_4542;
wire n_6892;
wire n_4462;
wire n_7061;
wire n_6401;
wire n_7322;
wire n_1716;
wire n_278;
wire n_6685;
wire n_4931;
wire n_4536;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_7051;
wire n_384;
wire n_8477;
wire n_1976;
wire n_7880;
wire n_4382;
wire n_2905;
wire n_1291;
wire n_8230;
wire n_6679;
wire n_8092;
wire n_749;
wire n_1824;
wire n_3954;
wire n_5911;
wire n_2122;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_6574;
wire n_6571;
wire n_5577;
wire n_1255;
wire n_568;
wire n_8876;
wire n_5124;
wire n_143;
wire n_3951;
wire n_8829;
wire n_823;
wire n_7824;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_7094;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_8140;
wire n_5413;
wire n_8971;
wire n_8060;
wire n_1338;
wire n_1097;
wire n_3027;
wire n_781;
wire n_4083;
wire n_7036;
wire n_6392;
wire n_1810;
wire n_182;
wire n_5915;
wire n_8527;
wire n_573;
wire n_9049;
wire n_7351;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_2295;
wire n_2746;
wire n_389;
wire n_814;
wire n_7608;
wire n_5779;
wire n_1643;
wire n_2020;
wire n_6260;
wire n_6832;
wire n_7394;
wire n_7909;
wire n_7413;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_222;
wire n_6286;
wire n_7675;
wire n_8267;
wire n_4023;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_6912;
wire n_721;
wire n_1461;
wire n_742;
wire n_7175;
wire n_691;
wire n_3617;
wire n_8276;
wire n_2076;
wire n_6019;
wire n_3567;
wire n_377;
wire n_1598;
wire n_7524;
wire n_4344;
wire n_2935;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_3807;
wire n_8925;
wire n_6214;
wire n_918;
wire n_1114;
wire n_763;
wire n_4027;
wire n_3154;
wire n_7783;
wire n_6692;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_3520;
wire n_191;
wire n_8978;
wire n_8093;
wire n_8245;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_946;
wire n_1303;
wire n_8454;
wire n_6552;
wire n_4095;
wire n_8327;
wire n_2881;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_8891;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_1780;
wire n_3897;
wire n_1689;
wire n_5591;
wire n_3372;
wire n_7697;
wire n_1944;
wire n_6403;
wire n_7306;
wire n_1347;
wire n_7947;
wire n_795;
wire n_1221;
wire n_7470;
wire n_7547;
wire n_7733;
wire n_6013;
wire n_1245;
wire n_7693;
wire n_3215;
wire n_6491;
wire n_448;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_6348;
wire n_6744;
wire n_1561;
wire n_8582;
wire n_1112;
wire n_6982;
wire n_5518;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_6661;
wire n_6293;
wire n_234;
wire n_5847;
wire n_7345;
wire n_6049;
wire n_1460;
wire n_911;
wire n_8847;
wire n_8957;
wire n_7385;
wire n_5159;
wire n_2862;
wire n_472;
wire n_2615;
wire n_4068;
wire n_6558;
wire n_4625;
wire n_2474;
wire n_3703;
wire n_2444;
wire n_2437;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_8488;
wire n_4863;
wire n_2267;
wire n_3035;
wire n_668;
wire n_4166;
wire n_8356;
wire n_1821;
wire n_6136;
wire n_1058;
wire n_3378;
wire n_6855;
wire n_3745;
wire n_3362;
wire n_4744;
wire n_8888;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_2222;
wire n_712;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_6551;
wire n_7691;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_6312;
wire n_8747;
wire n_2505;
wire n_334;
wire n_4817;
wire n_6668;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_470;
wire n_7653;
wire n_3680;
wire n_5381;
wire n_8354;
wire n_2408;
wire n_5723;
wire n_6859;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_8353;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_9027;
wire n_1972;
wire n_4383;
wire n_6995;
wire n_4491;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_455;
wire n_8211;
wire n_363;
wire n_4486;
wire n_6971;
wire n_1816;
wire n_393;
wire n_503;
wire n_6131;
wire n_5848;
wire n_3024;
wire n_7475;
wire n_4612;
wire n_6435;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_6351;
wire n_5163;
wire n_7668;
wire n_6212;
wire n_307;
wire n_4529;
wire n_500;
wire n_3361;
wire n_714;
wire n_3478;
wire n_8018;
wire n_8653;
wire n_3936;
wire n_1349;
wire n_291;
wire n_8920;
wire n_7937;
wire n_6829;
wire n_2723;
wire n_5485;
wire n_7819;
wire n_5823;
wire n_7305;
wire n_2800;
wire n_3496;
wire n_5473;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_4390;
wire n_3096;
wire n_8678;
wire n_2651;
wire n_8884;
wire n_8803;
wire n_2095;
wire n_3239;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_8222;
wire n_6822;
wire n_4062;
wire n_3902;
wire n_3295;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_1998;
wire n_1574;
wire n_3101;
wire n_240;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_3374;
wire n_2640;
wire n_253;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_8751;
wire n_4307;
wire n_3992;
wire n_3876;
wire n_249;
wire n_3125;
wire n_7391;
wire n_8790;
wire n_6617;
wire n_4293;
wire n_941;
wire n_3552;
wire n_1031;
wire n_115;
wire n_7511;
wire n_6533;
wire n_849;
wire n_4684;
wire n_3116;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_1753;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_2471;
wire n_8338;
wire n_6983;
wire n_8398;
wire n_4412;
wire n_2807;
wire n_8178;
wire n_6801;
wire n_1921;
wire n_8491;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_5630;
wire n_4758;
wire n_4781;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_271;
wire n_206;
wire n_4057;
wire n_633;
wire n_1170;
wire n_5379;
wire n_5335;
wire n_308;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_6113;
wire n_2634;
wire n_1761;
wire n_5424;
wire n_8750;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_8560;
wire n_2308;
wire n_2333;
wire n_8439;
wire n_3001;
wire n_1089;
wire n_3795;
wire n_7321;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_8200;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_8304;
wire n_3896;
wire n_3815;
wire n_6655;
wire n_8674;
wire n_5274;
wire n_3274;
wire n_5401;
wire n_7584;
wire n_4457;
wire n_7537;
wire n_4093;
wire n_1616;
wire n_8675;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_339;
wire n_434;
wire n_288;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_4794;
wire n_722;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_629;
wire n_1621;
wire n_9016;
wire n_2547;
wire n_2415;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_5073;
wire n_827;
wire n_8846;
wire n_8315;
wire n_4834;
wire n_8760;
wire n_4762;
wire n_192;
wire n_5581;
wire n_9029;
wire n_3113;
wire n_6837;
wire n_992;
wire n_3813;
wire n_3660;
wire n_3766;
wire n_1613;
wire n_1458;
wire n_5303;
wire n_7486;
wire n_6756;
wire n_1027;
wire n_3266;
wire n_7023;
wire n_3574;
wire n_7496;
wire n_1189;
wire n_223;
wire n_4154;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_7410;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_365;
wire n_3844;
wire n_8777;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_8535;
wire n_6373;
wire n_5375;
wire n_2451;
wire n_5370;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_5784;
wire n_5601;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_509;
wire n_4819;
wire n_1209;
wire n_7906;
wire n_5248;
wire n_1708;
wire n_7131;
wire n_805;
wire n_396;
wire n_6411;
wire n_350;
wire n_2051;
wire n_4370;
wire n_8909;
wire n_2359;
wire n_5112;
wire n_480;
wire n_142;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_7302;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_4645;
wire n_7797;
wire n_3668;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_7687;
wire n_2491;
wire n_1264;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_7582;
wire n_4933;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_287;
wire n_4302;
wire n_5111;
wire n_8959;
wire n_6534;
wire n_3340;
wire n_230;
wire n_5227;
wire n_7809;
wire n_461;
wire n_873;
wire n_3946;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_8425;
wire n_8087;
wire n_3395;
wire n_7060;
wire n_7607;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_2513;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_250;
wire n_1711;
wire n_4884;
wire n_1579;
wire n_7867;
wire n_3275;
wire n_8361;
wire n_836;
wire n_6135;
wire n_7761;
wire n_8007;
wire n_522;
wire n_3678;
wire n_6814;
wire n_3440;
wire n_8669;
wire n_8001;
wire n_2094;
wire n_7525;
wire n_1511;
wire n_2356;
wire n_7257;
wire n_7553;
wire n_1422;
wire n_7529;
wire n_1772;
wire n_4692;
wire n_6791;
wire n_616;
wire n_8496;
wire n_3165;
wire n_1119;
wire n_6824;
wire n_5788;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2739;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_641;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_7650;
wire n_3316;
wire n_8568;
wire n_516;
wire n_6903;
wire n_2418;
wire n_2864;
wire n_8852;
wire n_4311;
wire n_1180;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_6881;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_6450;
wire n_3261;
wire n_666;
wire n_7520;
wire n_4187;
wire n_6309;
wire n_940;
wire n_7903;
wire n_2058;
wire n_405;
wire n_213;
wire n_2660;
wire n_6733;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_1094;
wire n_8610;
wire n_5942;
wire n_5430;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_494;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_6300;
wire n_8256;
wire n_3532;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_3948;
wire n_9039;
wire n_8573;
wire n_2124;
wire n_8265;
wire n_4619;
wire n_381;
wire n_7639;
wire n_8704;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_5036;
wire n_4221;
wire n_3297;
wire n_6179;
wire n_6395;
wire n_976;
wire n_7605;
wire n_7054;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_5327;
wire n_2364;
wire n_4392;
wire n_2996;
wire n_7433;
wire n_8131;
wire n_3803;
wire n_2085;
wire n_8941;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_6171;
wire n_8775;
wire n_808;
wire n_5519;
wire n_4047;
wire n_6269;
wire n_5753;
wire n_3413;
wire n_7092;
wire n_6980;
wire n_1193;
wire n_5233;
wire n_3412;
wire n_8279;
wire n_6654;
wire n_8019;
wire n_3791;
wire n_6083;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_551;
wire n_699;
wire n_4320;
wire n_8257;
wire n_7832;
wire n_3884;
wire n_5808;
wire n_451;
wire n_8390;
wire n_8898;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_757;
wire n_594;
wire n_5231;
wire n_2190;
wire n_6120;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_3438;
wire n_166;
wire n_4141;
wire n_8464;
wire n_6547;
wire n_8799;
wire n_5193;
wire n_6423;
wire n_2850;
wire n_572;
wire n_6342;
wire n_6641;
wire n_1481;
wire n_6984;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_2104;
wire n_7441;
wire n_513;
wire n_7106;
wire n_7213;
wire n_3883;
wire n_5961;
wire n_261;
wire n_5866;
wire n_9050;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_6687;
wire n_121;
wire n_5822;
wire n_433;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_3949;
wire n_5726;
wire n_2792;
wire n_219;
wire n_5364;
wire n_3315;
wire n_7031;
wire n_263;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_788;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_329;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_7133;
wire n_4720;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_243;
wire n_1873;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_1866;
wire n_117;
wire n_8661;
wire n_2130;
wire n_7424;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_7523;
wire n_2228;
wire n_8654;
wire n_5039;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_6790;
wire n_8746;
wire n_5953;
wire n_3099;
wire n_8531;
wire n_7141;
wire n_5198;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_6459;
wire n_1663;
wire n_6505;
wire n_8379;
wire n_8609;
wire n_4172;
wire n_3403;
wire n_7626;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_1107;
wire n_2457;
wire n_3294;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_7311;
wire n_3686;
wire n_7669;
wire n_4502;
wire n_5958;
wire n_8793;
wire n_8103;
wire n_318;
wire n_2971;
wire n_1713;
wire n_715;
wire n_4526;
wire n_4277;
wire n_1265;
wire n_3490;
wire n_4849;
wire n_530;
wire n_277;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_8873;
wire n_8367;
wire n_618;
wire n_7367;
wire n_199;
wire n_5792;
wire n_3581;
wire n_8543;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_7323;
wire n_7189;
wire n_7301;
wire n_6258;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_6905;
wire n_612;
wire n_8682;
wire n_3725;
wire n_8089;
wire n_6704;
wire n_3933;
wire n_8533;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_1175;
wire n_7244;
wire n_7368;
wire n_2311;
wire n_429;
wire n_1012;
wire n_3691;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_903;
wire n_7633;
wire n_4146;
wire n_5711;
wire n_1802;
wire n_1504;
wire n_4340;
wire n_5790;
wire n_286;
wire n_8640;
wire n_254;
wire n_8063;
wire n_3961;
wire n_4855;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_7878;
wire n_6186;
wire n_6803;
wire n_816;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_1188;
wire n_7427;
wire n_2206;
wire n_4004;
wire n_2967;
wire n_5404;
wire n_2916;
wire n_5739;
wire n_4292;
wire n_8570;
wire n_6163;
wire n_7628;
wire n_5972;
wire n_2467;
wire n_5549;
wire n_267;
wire n_3145;
wire n_6785;
wire n_6553;
wire n_1124;
wire n_1624;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_3280;
wire n_8039;
wire n_5757;
wire n_1515;
wire n_8902;
wire n_8916;
wire n_961;
wire n_7557;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_593;
wire n_8843;
wire n_7128;
wire n_637;
wire n_2377;
wire n_701;
wire n_6849;
wire n_7594;
wire n_950;
wire n_8129;
wire n_8162;
wire n_7457;
wire n_8744;
wire n_3009;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_7788;
wire n_4361;
wire n_5488;
wire n_6760;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_7752;
wire n_3889;
wire n_2687;
wire n_1630;
wire n_2887;
wire n_4245;
wire n_4136;
wire n_8286;
wire n_3526;
wire n_2194;
wire n_2619;
wire n_5329;
wire n_9015;
wire n_4367;
wire n_5637;
wire n_6825;
wire n_1987;
wire n_7586;
wire n_6452;
wire n_507;
wire n_968;
wire n_7767;
wire n_8294;
wire n_2271;
wire n_1008;
wire n_6611;
wire n_8562;
wire n_2583;
wire n_4560;
wire n_2606;
wire n_4899;
wire n_5728;
wire n_5471;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_5164;
wire n_2391;
wire n_304;
wire n_2431;
wire n_7207;
wire n_8218;
wire n_5843;
wire n_8170;
wire n_7744;
wire n_125;
wire n_2078;
wire n_7021;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_7748;
wire n_8537;
wire n_3450;
wire n_6827;
wire n_449;
wire n_4663;
wire n_2893;
wire n_1208;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_2728;
wire n_1072;
wire n_815;
wire n_6227;
wire n_7215;
wire n_7485;
wire n_3421;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_1067;
wire n_3405;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_255;
wire n_284;
wire n_1952;
wire n_5074;
wire n_4044;
wire n_6564;
wire n_3436;
wire n_8709;
wire n_8782;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_289;
wire n_6468;
wire n_3937;
wire n_1293;
wire n_3159;
wire n_4701;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_6857;
wire n_3240;
wire n_8144;
wire n_3576;
wire n_1863;
wire n_3385;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_3293;
wire n_872;
wire n_3922;
wire n_8049;
wire n_7762;
wire n_5204;
wire n_5333;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_5422;
wire n_6871;
wire n_1513;
wire n_1913;
wire n_4934;
wire n_837;
wire n_8357;
wire n_6904;
wire n_5087;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_7017;
wire n_7777;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_7652;
wire n_5551;
wire n_3150;
wire n_8701;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_6499;
wire n_7830;
wire n_4011;
wire n_5131;
wire n_1959;
wire n_3133;
wire n_7138;
wire n_5257;
wire n_8097;
wire n_765;
wire n_1492;
wire n_8084;
wire n_8645;
wire n_1340;
wire n_4688;
wire n_4753;
wire n_8712;
wire n_4058;
wire n_631;
wire n_8289;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_7966;
wire n_8591;
wire n_5059;
wire n_156;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_843;
wire n_8824;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_7191;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_5242;
wire n_5219;
wire n_8417;
wire n_2675;
wire n_6276;
wire n_5631;
wire n_3537;
wire n_8340;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_1022;
wire n_614;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_8455;
wire n_7208;
wire n_2119;
wire n_947;
wire n_1117;
wire n_7961;
wire n_1992;
wire n_5686;
wire n_5899;
wire n_6893;
wire n_7406;
wire n_8681;
wire n_8905;
wire n_3223;
wire n_3140;
wire n_7807;
wire n_3185;
wire n_4749;
wire n_2605;
wire n_5155;
wire n_7680;
wire n_118;
wire n_926;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_8172;
wire n_1698;
wire n_8106;
wire n_4100;
wire n_6447;
wire n_4264;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_5937;
wire n_777;
wire n_6422;
wire n_1299;
wire n_6751;
wire n_5339;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_3325;
wire n_2238;
wire n_6040;
wire n_8375;
wire n_4085;
wire n_4464;
wire n_8612;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_4659;
wire n_3600;
wire n_6741;
wire n_8459;
wire n_5217;
wire n_5465;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_8268;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_6160;
wire n_6650;
wire n_8221;
wire n_7066;
wire n_8255;
wire n_7183;
wire n_796;
wire n_1195;
wire n_7789;
wire n_184;
wire n_7606;
wire n_8461;
wire n_6192;
wire n_1811;
wire n_6368;
wire n_7140;
wire n_7193;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_6039;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_1142;
wire n_623;
wire n_1048;
wire n_5721;
wire n_3638;
wire n_4816;
wire n_8515;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_8812;
wire n_6012;
wire n_3451;
wire n_1418;
wire n_1250;
wire n_292;
wire n_4937;
wire n_5277;
wire n_8792;
wire n_3615;
wire n_7344;
wire n_3072;
wire n_3087;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_4222;
wire n_6707;
wire n_4874;
wire n_4401;
wire n_889;
wire n_2710;
wire n_6064;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_477;
wire n_6787;
wire n_8523;
wire n_1110;
wire n_4709;
wire n_2213;
wire n_7710;
wire n_4976;
wire n_2389;
wire n_7892;
wire n_2132;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_1564;
wire n_5578;
wire n_4658;
wire n_231;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_1457;
wire n_505;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_1787;
wire n_6769;
wire n_537;
wire n_1993;
wire n_2281;
wire n_8406;
wire n_6277;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_3705;
wire n_3211;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_8554;
wire n_546;
wire n_386;
wire n_1220;
wire n_6051;
wire n_1893;
wire n_8896;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_7206;
wire n_4223;
wire n_7538;
wire n_2387;
wire n_5674;
wire n_3270;
wire n_5539;
wire n_6895;
wire n_2846;
wire n_5282;
wire n_970;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_6799;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_444;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_7716;
wire n_6487;
wire n_511;
wire n_5121;
wire n_8758;
wire n_6026;
wire n_6070;
wire n_1286;
wire n_8818;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_4348;
wire n_5013;
wire n_1597;
wire n_6807;
wire n_8954;
wire n_7251;
wire n_4489;
wire n_4839;
wire n_7254;
wire n_2596;
wire n_3163;
wire n_7540;
wire n_775;
wire n_4404;
wire n_1153;
wire n_5589;
wire n_439;
wire n_6563;
wire n_1531;
wire n_7882;
wire n_2828;
wire n_453;
wire n_8552;
wire n_7554;
wire n_2384;
wire n_8069;
wire n_7558;
wire n_4261;
wire n_4204;
wire n_8373;
wire n_759;
wire n_2724;
wire n_426;
wire n_6481;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_4006;
wire n_2226;
wire n_2801;
wire n_6341;
wire n_6384;
wire n_1901;
wire n_3869;
wire n_7421;
wire n_2556;
wire n_7489;
wire n_4747;
wire n_6906;
wire n_7541;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_3742;
wire n_3683;
wire n_8318;
wire n_4801;
wire n_401;
wire n_3260;
wire n_2550;
wire n_8341;
wire n_3175;
wire n_7188;
wire n_3736;
wire n_5475;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_7991;
wire n_6233;
wire n_2227;
wire n_6377;
wire n_5216;
wire n_3284;
wire n_4869;
wire n_8239;
wire n_427;
wire n_8926;
wire n_6257;
wire n_2159;
wire n_688;
wire n_2315;
wire n_1077;
wire n_4386;
wire n_4132;
wire n_2995;
wire n_5273;
wire n_7898;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_4955;
wire n_8965;
wire n_4149;
wire n_5936;
wire n_4355;
wire n_7646;
wire n_501;
wire n_2276;
wire n_3234;
wire n_856;
wire n_2803;
wire n_8817;
wire n_379;
wire n_8190;
wire n_1668;
wire n_2777;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_6587;
wire n_1129;
wire n_7781;
wire n_6987;
wire n_602;
wire n_7360;
wire n_2181;
wire n_6069;
wire n_171;
wire n_2911;
wire n_7497;
wire n_169;
wire n_4655;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_7665;
wire n_3429;
wire n_2379;
wire n_326;
wire n_7793;
wire n_587;
wire n_8355;
wire n_3554;
wire n_1593;
wire n_6991;
wire n_1202;
wire n_7101;
wire n_7671;
wire n_1635;
wire n_7530;
wire n_8489;
wire n_5431;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_7204;
wire n_8649;
wire n_6887;
wire n_7578;
wire n_3462;
wire n_7654;
wire n_2851;
wire n_8303;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_8369;
wire n_9022;
wire n_358;
wire n_160;
wire n_8059;
wire n_6633;
wire n_2420;
wire n_5627;
wire n_5774;
wire n_6579;
wire n_3722;
wire n_186;
wire n_4846;
wire n_4400;
wire n_5798;
wire n_2984;
wire n_575;
wire n_5187;
wire n_5875;
wire n_4024;
wire n_8831;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_732;
wire n_6569;
wire n_2983;
wire n_6335;
wire n_7120;
wire n_8728;
wire n_2240;
wire n_392;
wire n_2538;
wire n_724;
wire n_3250;
wire n_6789;
wire n_8386;
wire n_8853;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_6252;
wire n_557;
wire n_1871;
wire n_4860;
wire n_6211;
wire n_845;
wire n_140;
wire n_5844;
wire n_8862;
wire n_3414;
wire n_1549;
wire n_4870;
wire n_6164;
wire n_768;
wire n_7576;
wire n_6173;
wire n_8081;
wire n_7786;
wire n_3651;
wire n_7313;
wire n_2102;
wire n_2563;
wire n_4989;
wire n_7676;
wire n_7609;
wire n_7757;
wire n_3449;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_8900;
wire n_597;
wire n_280;
wire n_6630;
wire n_6934;
wire n_9017;
wire n_1187;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_6737;
wire n_4488;
wire n_3767;
wire n_8396;
wire n_6612;
wire n_8478;
wire n_6606;
wire n_2544;
wire n_6695;
wire n_3550;
wire n_8865;
wire n_4211;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_1206;
wire n_4016;
wire n_5867;
wire n_621;
wire n_750;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_3839;
wire n_8497;
wire n_2823;
wire n_8820;
wire n_6410;
wire n_6158;
wire n_5597;
wire n_9028;
wire n_4915;
wire n_4328;
wire n_6413;
wire n_8020;
wire n_6090;
wire n_1057;
wire n_7419;
wire n_6506;
wire n_2785;
wire n_235;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1818;
wire n_3730;
wire n_6935;
wire n_1298;
wire n_5862;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_1611;
wire n_5050;
wire n_2740;
wire n_746;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_3416;
wire n_3498;
wire n_5767;
wire n_2401;
wire n_8992;
wire n_1589;
wire n_4712;
wire n_8880;
wire n_8690;
wire n_2309;
wire n_2900;
wire n_6234;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_1497;
wire n_6688;
wire n_133;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_8770;
wire n_3672;
wire n_7182;
wire n_5318;
wire n_7365;
wire n_6608;
wire n_3533;
wire n_1622;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_8075;
wire n_6798;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_7885;
wire n_6860;
wire n_6557;
wire n_8466;
wire n_6753;
wire n_2171;
wire n_6527;
wire n_7341;
wire n_2988;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_8094;
wire n_4109;
wire n_4192;
wire n_6639;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_6430;
wire n_5150;
wire n_782;
wire n_809;
wire n_8832;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_1797;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_402;
wire n_1870;
wire n_1171;
wire n_460;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_1827;
wire n_4904;
wire n_2187;
wire n_7517;
wire n_1152;
wire n_6627;
wire n_8080;
wire n_450;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_6058;
wire n_711;
wire n_7745;
wire n_3105;
wire n_2872;
wire n_6666;
wire n_3692;
wire n_4616;
wire n_8321;
wire n_8772;
wire n_8735;
wire n_4982;
wire n_370;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_8592;
wire n_8786;
wire n_8684;
wire n_6190;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_6249;
wire n_2738;
wire n_972;
wire n_8083;
wire n_5348;
wire n_6594;
wire n_1332;
wire n_5480;
wire n_4323;
wire n_624;
wire n_8157;
wire n_2346;
wire n_4831;
wire n_7095;
wire n_936;
wire n_3045;
wire n_3821;
wire n_6969;
wire n_885;
wire n_7459;
wire n_6161;
wire n_6615;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_7294;
wire n_3676;
wire n_4896;
wire n_8206;
wire n_2882;
wire n_3675;
wire n_3666;
wire n_4017;
wire n_4260;
wire n_4916;
wire n_2541;
wire n_8622;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_7184;
wire n_6607;
wire n_599;
wire n_6062;
wire n_7908;
wire n_1974;
wire n_4122;
wire n_7974;
wire n_7551;
wire n_934;
wire n_4209;
wire n_8104;
wire n_8344;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_4298;
wire n_2314;
wire n_8120;
wire n_3502;
wire n_8513;
wire n_5461;
wire n_3003;
wire n_6482;
wire n_4128;
wire n_6294;
wire n_543;
wire n_5147;
wire n_4271;
wire n_4644;
wire n_9021;
wire n_1355;
wire n_8779;
wire n_2258;
wire n_8621;
wire n_5503;
wire n_325;
wire n_5845;
wire n_5945;
wire n_804;
wire n_2390;
wire n_6246;
wire n_8868;
wire n_959;
wire n_2562;
wire n_8134;
wire n_4716;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_7250;
wire n_1782;
wire n_5755;
wire n_5600;
wire n_8762;
wire n_8043;
wire n_8694;
wire n_707;
wire n_1900;
wire n_5048;
wire n_6053;
wire n_7252;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_3208;
wire n_2195;
wire n_4944;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_6901;
wire n_4935;
wire n_4694;
wire n_8191;
wire n_6841;
wire n_4672;
wire n_8101;
wire n_5054;
wire n_2962;
wire n_8376;
wire n_8171;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_2939;
wire n_7698;
wire n_5749;
wire n_1672;
wire n_6774;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_1925;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_8710;
wire n_737;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_4598;
wire n_3061;
wire n_3893;
wire n_3932;
wire n_3469;
wire n_8599;
wire n_2960;
wire n_8549;
wire n_5993;
wire n_8054;
wire n_6716;
wire n_138;
wire n_3258;
wire n_8616;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_333;
wire n_4084;
wire n_3149;
wire n_6844;
wire n_7914;
wire n_8628;
wire n_3365;
wire n_6521;
wire n_7891;
wire n_3379;
wire n_8857;
wire n_8517;
wire n_459;
wire n_4850;
wire n_8547;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_3008;
wire n_1751;
wire n_6162;
wire n_2840;
wire n_6779;
wire n_8010;
wire n_285;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_1375;
wire n_3972;
wire n_4153;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_7216;
wire n_1928;
wire n_3091;
wire n_4317;
wire n_8275;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_6762;
wire n_6178;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_9035;
wire n_1019;
wire n_8291;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_3642;
wire n_2845;
wire n_4650;
wire n_7706;
wire n_438;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_479;
wire n_6458;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_7642;
wire n_8247;
wire n_6577;
wire n_6740;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_6315;
wire n_2366;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_2210;
wire n_7156;
wire n_4735;
wire n_3602;
wire n_187;
wire n_3300;
wire n_2978;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_6910;
wire n_6262;
wire n_7604;
wire n_2827;
wire n_1177;
wire n_7703;
wire n_3515;
wire n_1150;
wire n_6319;
wire n_566;
wire n_1023;
wire n_2951;
wire n_1118;
wire n_194;
wire n_2949;
wire n_1807;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_6536;
wire n_256;
wire n_440;
wire n_6175;
wire n_3806;
wire n_7040;
wire n_8827;
wire n_8280;
wire n_5514;
wire n_2931;
wire n_209;
wire n_367;
wire n_8388;
wire n_2569;
wire n_3866;
wire n_6978;
wire n_5351;
wire n_5909;
wire n_671;
wire n_6093;
wire n_4543;
wire n_740;
wire n_7378;
wire n_703;
wire n_4157;
wire n_8988;
wire n_6845;
wire n_6947;
wire n_4229;
wire n_5293;
wire n_8203;
wire n_6099;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_8569;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_8877;
wire n_1401;
wire n_7498;
wire n_1516;
wire n_3846;
wire n_6321;
wire n_180;
wire n_3512;
wire n_6819;
wire n_5201;
wire n_2029;
wire n_7501;
wire n_5890;
wire n_6415;
wire n_6465;
wire n_4439;
wire n_1394;
wire n_1326;
wire n_4783;
wire n_1379;
wire n_214;
wire n_7931;
wire n_8688;
wire n_935;
wire n_4910;
wire n_1130;
wire n_3083;
wire n_6899;
wire n_7549;
wire n_7373;
wire n_7895;
wire n_676;
wire n_832;
wire n_6592;
wire n_3049;
wire n_8686;
wire n_8871;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_9011;
wire n_8418;
wire n_3830;
wire n_7740;
wire n_8403;
wire n_3679;
wire n_5891;
wire n_7613;
wire n_3541;
wire n_6101;
wire n_3117;
wire n_5935;
wire n_7556;
wire n_4930;
wire n_372;
wire n_8588;
wire n_314;
wire n_378;
wire n_5623;
wire n_8564;
wire n_6944;
wire n_338;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_506;
wire n_360;
wire n_2149;
wire n_9012;
wire n_2396;
wire n_4557;
wire n_4917;
wire n_8698;
wire n_895;
wire n_8924;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_4593;
wire n_7238;
wire n_344;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_8780;
wire n_7309;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_1392;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_525;
wire n_2463;
wire n_3363;
wire n_7572;
wire n_8214;
wire n_1677;
wire n_5990;
wire n_611;
wire n_7043;
wire n_3721;
wire n_3062;
wire n_2679;
wire n_5024;
wire n_7760;
wire n_4559;
wire n_8514;
wire n_8722;
wire n_8241;
wire n_8589;
wire n_838;
wire n_3969;
wire n_129;
wire n_3336;
wire n_7573;
wire n_4160;
wire n_8442;
wire n_4231;
wire n_6281;
wire n_7364;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_8608;
wire n_5203;
wire n_6846;
wire n_6311;
wire n_445;
wire n_930;
wire n_7590;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_1945;
wire n_5426;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_1414;
wire n_5285;
wire n_7048;
wire n_6886;
wire n_2721;
wire n_944;
wire n_4335;
wire n_2034;
wire n_576;
wire n_6593;
wire n_8630;
wire n_270;
wire n_2683;
wire n_563;
wire n_5365;
wire n_8583;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_8145;
wire n_8405;
wire n_7176;
wire n_8928;
wire n_7682;
wire n_626;
wire n_990;
wire n_6231;
wire n_8948;
wire n_8672;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_6746;
wire n_498;
wire n_8447;
wire n_7901;
wire n_870;
wire n_5395;
wire n_1253;
wire n_366;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_1693;
wire n_6446;
wire n_7980;
wire n_3256;
wire n_348;
wire n_3802;
wire n_7218;
wire n_6996;
wire n_8828;
wire n_376;
wire n_2118;
wire n_2111;
wire n_390;
wire n_2915;
wire n_1148;
wire n_6749;
wire n_2188;
wire n_8440;
wire n_1989;
wire n_7005;
wire n_2802;
wire n_8572;
wire n_7732;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_7447;
wire n_2425;
wire n_6777;
wire n_4265;
wire n_8227;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_8475;
wire n_3060;
wire n_3098;
wire n_6924;
wire n_8029;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_4064;
wire n_7405;
wire n_4926;
wire n_1518;
wire n_1362;
wire n_3123;
wire n_8314;
wire n_3380;
wire n_5617;
wire n_1829;
wire n_7922;
wire n_5580;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_3038;
wire n_570;
wire n_1789;
wire n_6310;
wire n_620;
wire n_519;
wire n_8311;
wire n_2523;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_5310;
wire n_8764;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_5390;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_6683;
wire n_4769;
wire n_5764;
wire n_8934;
wire n_2282;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_2047;
wire n_8407;
wire n_6229;
wire n_8567;
wire n_5385;
wire n_1609;
wire n_8729;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_409;
wire n_1763;
wire n_5322;
wire n_6907;
wire n_3989;
wire n_7144;
wire n_2490;
wire n_7089;
wire n_7286;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_635;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_4254;
wire n_8253;
wire n_6177;
wire n_1996;
wire n_6332;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_8283;
wire n_5982;
wire n_1158;
wire n_2248;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_5011;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_2662;
wire n_3147;
wire n_4909;
wire n_6696;
wire n_753;
wire n_3925;
wire n_3180;
wire n_8566;
wire n_7343;
wire n_2795;
wire n_3472;
wire n_8516;
wire n_8302;
wire n_8317;
wire n_5376;
wire n_5106;
wire n_269;
wire n_6116;
wire n_359;
wire n_8167;
wire n_7859;
wire n_6730;
wire n_7492;
wire n_7872;
wire n_7972;
wire n_1479;
wire n_4768;
wire n_1675;
wire n_7916;
wire n_3717;
wire n_7480;
wire n_7694;
wire n_5561;
wire n_5410;
wire n_571;
wire n_2215;
wire n_404;
wire n_8944;
wire n_6167;
wire n_158;
wire n_1884;
wire n_8008;
wire n_6170;
wire n_665;
wire n_8109;
wire n_2055;
wire n_5156;
wire n_2553;
wire n_6307;
wire n_149;
wire n_632;
wire n_6094;
wire n_2038;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_7434;
wire n_4826;
wire n_3445;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_373;
wire n_8975;
wire n_6267;
wire n_7787;
wire n_1833;
wire n_3903;
wire n_5998;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_6568;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_5378;
wire n_6028;
wire n_1417;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_5916;
wire n_681;
wire n_4648;
wire n_3094;
wire n_412;
wire n_8697;
wire n_6299;
wire n_6813;
wire n_965;
wire n_8825;
wire n_1428;
wire n_1576;
wire n_1856;
wire n_2077;
wire n_7425;
wire n_6669;
wire n_8581;
wire n_8266;
wire n_5691;
wire n_1059;
wire n_4951;
wire n_8981;
wire n_422;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_3079;
wire n_165;
wire n_4360;
wire n_8771;
wire n_540;
wire n_4039;
wire n_457;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_1748;
wire n_8639;
wire n_8058;
wire n_8138;
wire n_3504;
wire n_6638;
wire n_531;
wire n_7719;
wire n_4272;
wire n_8333;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_6220;
wire n_7562;
wire n_3111;
wire n_336;
wire n_6985;
wire n_7619;
wire n_7170;
wire n_1885;
wire n_8176;
wire n_8124;
wire n_8823;
wire n_7366;
wire n_5269;
wire n_9026;
wire n_3054;
wire n_1538;
wire n_8147;
wire n_1240;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_1234;
wire n_5262;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_4882;
wire n_4620;
wire n_3152;
wire n_7935;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_8458;
wire n_6772;
wire n_8113;
wire n_3335;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_1003;
wire n_5713;
wire n_5256;
wire n_168;
wire n_6318;
wire n_2353;
wire n_4099;
wire n_7918;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_6916;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_6651;
wire n_1923;
wire n_2260;
wire n_3952;
wire n_7845;
wire n_5550;
wire n_3911;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_1743;
wire n_6366;
wire n_6230;
wire n_2997;
wire n_6604;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_3708;
wire n_4078;
wire n_3046;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5939;
wire n_5509;
wire n_8160;
wire n_6391;
wire n_5382;
wire n_5659;
wire n_8099;
wire n_8840;
wire n_3619;
wire n_1415;
wire n_5881;
wire n_8522;
wire n_1370;
wire n_7222;
wire n_1786;
wire n_7942;
wire n_6473;
wire n_8578;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2291;
wire n_415;
wire n_1371;
wire n_7725;
wire n_383;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_200;
wire n_2184;
wire n_2982;
wire n_6483;
wire n_1803;
wire n_4065;
wire n_5863;
wire n_229;
wire n_7647;
wire n_8626;
wire n_2645;
wire n_3904;
wire n_8611;
wire n_8036;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_8819;
wire n_2630;
wire n_1444;
wire n_1603;
wire n_7300;
wire n_6697;
wire n_7875;
wire n_6975;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_4417;
wire n_5466;
wire n_7643;
wire n_4733;
wire n_6728;
wire n_6729;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_2286;
wire n_4743;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_5955;
wire n_7242;
wire n_658;
wire n_1874;
wire n_2865;
wire n_2825;
wire n_8441;
wire n_2013;
wire n_6076;
wire n_8933;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_7778;
wire n_758;
wire n_5851;
wire n_7073;
wire n_2256;
wire n_943;
wire n_4060;
wire n_5110;
wire n_8397;
wire n_4879;
wire n_6390;
wire n_5796;
wire n_772;
wire n_8726;
wire n_2806;
wire n_6665;
wire n_8797;
wire n_7224;
wire n_770;
wire n_3028;
wire n_7746;
wire n_3662;
wire n_2981;
wire n_6958;
wire n_3076;
wire n_886;
wire n_7563;
wire n_343;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_6549;
wire n_539;
wire n_8414;
wire n_6297;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_6096;
wire n_4117;
wire n_7853;
wire n_4687;
wire n_2836;
wire n_7531;
wire n_638;
wire n_1404;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_8615;
wire n_2378;
wire n_7721;
wire n_887;
wire n_7192;
wire n_5905;
wire n_2655;
wire n_4600;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_126;
wire n_1467;
wire n_8316;
wire n_4250;
wire n_5829;
wire n_3906;
wire n_224;
wire n_8057;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_8505;
wire n_3963;
wire n_3368;
wire n_7884;
wire n_2370;
wire n_2612;
wire n_8970;
wire n_7527;
wire n_7417;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_2214;
wire n_4253;
wire n_407;
wire n_913;
wire n_6582;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_7388;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_8717;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_3189;
wire n_7635;
wire n_5525;
wire n_163;
wire n_1644;
wire n_2725;
wire n_2277;
wire n_7090;
wire n_4691;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_8571;
wire n_4305;
wire n_7227;
wire n_7415;
wire n_824;
wire n_6745;
wire n_6972;
wire n_4297;
wire n_8030;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_2907;
wire n_577;
wire n_5374;
wire n_5575;
wire n_8725;
wire n_1843;
wire n_619;
wire n_5675;
wire n_4227;
wire n_521;
wire n_2778;
wire n_395;
wire n_1909;
wire n_6240;
wire n_8243;
wire n_6347;
wire n_8633;
wire n_5020;
wire n_7689;
wire n_6511;
wire n_606;
wire n_5297;
wire n_7121;
wire n_1309;
wire n_1123;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_483;
wire n_6804;
wire n_1970;
wire n_8449;
wire n_6358;
wire n_630;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_6603;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_476;
wire n_4364;
wire n_7534;
wire n_1957;
wire n_8201;
wire n_8967;
wire n_4354;
wire n_6986;
wire n_8801;
wire n_3912;
wire n_4732;
wire n_3118;
wire n_5959;
wire n_3720;
wire n_1907;
wire n_2529;
wire n_8031;
wire n_8918;
wire n_264;
wire n_860;
wire n_8219;
wire n_1530;
wire n_8696;
wire n_4745;
wire n_938;
wire n_1302;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_4581;
wire n_6890;
wire n_549;
wire n_4377;
wire n_7827;
wire n_2143;
wire n_8180;
wire n_905;
wire n_6109;
wire n_4792;
wire n_7731;
wire n_1680;
wire n_3842;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_4979;
wire n_1988;
wire n_558;
wire n_6770;
wire n_2654;
wire n_3036;
wire n_7943;
wire n_8892;
wire n_5302;
wire n_966;
wire n_4511;
wire n_2908;
wire n_3357;
wire n_692;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_487;
wire n_8943;
wire n_8486;
wire n_241;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_2459;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_7132;
wire n_2711;
wire n_7081;
wire n_4199;
wire n_5885;
wire n_6663;
wire n_1912;
wire n_5356;
wire n_4441;
wire n_7319;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_1312;
wire n_8155;
wire n_5668;
wire n_5038;
wire n_268;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_2664;
wire n_1722;
wire n_1664;
wire n_5463;
wire n_3022;
wire n_8098;
wire n_247;
wire n_8833;
wire n_5489;
wire n_1165;
wire n_5892;
wire n_7828;
wire n_4773;
wire n_7940;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_2008;
wire n_6009;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_9034;
wire n_328;
wire n_1386;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_5113;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_8074;
wire n_8485;
wire n_8860;
wire n_5510;
wire n_2676;
wire n_3940;
wire n_6621;
wire n_7001;
wire n_4822;
wire n_1214;
wire n_690;
wire n_850;
wire n_8271;
wire n_5692;
wire n_8473;
wire n_4800;
wire n_1157;
wire n_3453;
wire n_5555;
wire n_3410;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_6783;
wire n_825;
wire n_6066;
wire n_8699;
wire n_3785;
wire n_6897;
wire n_2963;
wire n_8587;
wire n_5366;
wire n_2602;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_8225;
wire n_2980;
wire n_696;
wire n_4886;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_6296;
wire n_7708;
wire n_4055;
wire n_2178;
wire n_5968;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_6497;
wire n_8319;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_7108;
wire n_6470;
wire n_1796;
wire n_8368;
wire n_8322;
wire n_7333;
wire n_2082;
wire n_3519;
wire n_6187;
wire n_7876;
wire n_8546;
wire n_8300;
wire n_7371;
wire n_8152;
wire n_678;
wire n_7463;
wire n_8525;
wire n_6573;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_283;
wire n_8148;
wire n_8150;
wire n_3578;
wire n_909;
wire n_6693;
wire n_4737;
wire n_590;
wire n_4925;
wire n_4116;
wire n_5415;
wire n_8986;
wire n_362;
wire n_7285;
wire n_5419;
wire n_1990;
wire n_3805;
wire n_8929;
wire n_7260;
wire n_2943;
wire n_5205;
wire n_6409;
wire n_1634;
wire n_3252;
wire n_627;
wire n_3253;
wire n_7954;
wire n_1465;
wire n_342;
wire n_2622;
wire n_7951;
wire n_2658;
wire n_7552;
wire n_8096;
wire n_2665;
wire n_2133;
wire n_1712;
wire n_6130;
wire n_4603;
wire n_8233;
wire n_7273;
wire n_1523;
wire n_7231;
wire n_1627;
wire n_5080;
wire n_5976;
wire n_3128;
wire n_1527;
wire n_495;
wire n_5732;
wire n_5372;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_7449;
wire n_7772;
wire n_2230;
wire n_8763;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_8679;
wire n_1565;
wire n_7239;
wire n_1493;
wire n_5690;
wire n_8187;
wire n_7050;
wire n_8996;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_6623;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_615;
wire n_3838;
wire n_5371;
wire n_4651;
wire n_3941;
wire n_3793;
wire n_8139;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_605;
wire n_1514;
wire n_7597;
wire n_5801;
wire n_6047;
wire n_8292;
wire n_3037;
wire n_1646;
wire n_3729;
wire n_8601;
wire n_4994;
wire n_6652;
wire n_2537;
wire n_8830;
wire n_4483;
wire n_6921;
wire n_6970;
wire n_5347;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_4988;
wire n_7674;
wire n_3171;
wire n_7568;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_4540;
wire n_6344;
wire n_2097;
wire n_3459;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_3499;
wire n_6624;
wire n_6956;
wire n_4284;
wire n_6305;
wire n_1005;
wire n_1947;
wire n_6209;
wire n_8310;
wire n_3426;
wire n_4971;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_7329;
wire n_8646;
wire n_7408;
wire n_2650;
wire n_7107;
wire n_5652;
wire n_6457;
wire n_8597;
wire n_987;
wire n_7690;
wire n_8969;
wire n_7123;
wire n_5499;
wire n_720;
wire n_8117;
wire n_153;
wire n_3348;
wire n_3229;
wire n_1707;
wire n_656;
wire n_6950;
wire n_8208;
wire n_9048;
wire n_5228;
wire n_797;
wire n_2933;
wire n_2717;
wire n_1723;
wire n_1878;
wire n_189;
wire n_738;
wire n_2012;
wire n_6694;
wire n_3497;
wire n_6880;
wire n_5066;
wire n_7418;
wire n_2842;
wire n_3580;
wire n_2335;
wire n_8536;
wire n_7229;
wire n_8350;
wire n_529;
wire n_2307;
wire n_3704;
wire n_684;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_8328;
wire n_8914;
wire n_1181;
wire n_7258;
wire n_5190;
wire n_8391;
wire n_3173;
wire n_3677;
wire n_8336;
wire n_6856;
wire n_3996;
wire n_1049;
wire n_6466;
wire n_7864;
wire n_6727;
wire n_4097;
wire n_1666;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_2449;
wire n_3880;
wire n_3685;
wire n_8216;
wire n_2868;
wire n_7709;
wire n_2231;
wire n_3609;
wire n_1228;
wire n_5455;
wire n_417;
wire n_5442;
wire n_6386;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_272;
wire n_6820;
wire n_2896;
wire n_8313;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_7656;
wire n_2898;
wire n_5511;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_2368;
wire n_8041;
wire n_8202;
wire n_8263;
wire n_458;
wire n_4175;
wire n_6438;
wire n_5490;
wire n_3200;
wire n_4771;
wire n_7332;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_3867;
wire n_3593;
wire n_4455;
wire n_8374;
wire n_1073;
wire n_252;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_5584;
wire n_7512;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_7766;
wire n_8738;
wire n_6469;
wire n_6700;
wire n_2682;
wire n_3032;
wire n_6223;
wire n_6758;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_8798;
wire n_2877;
wire n_8085;
wire n_5098;
wire n_1021;
wire n_8123;
wire n_7955;
wire n_811;
wire n_683;
wire n_1207;
wire n_5707;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_7287;
wire n_5497;
wire n_8721;
wire n_880;
wire n_6464;
wire n_6356;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_7637;
wire n_2432;
wire n_150;
wire n_1478;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3777;
wire n_4203;
wire n_3641;
wire n_7127;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_5481;
wire n_3590;
wire n_8666;
wire n_2435;
wire n_5344;
wire n_954;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_7638;
wire n_1382;
wire n_7801;
wire n_5408;
wire n_1736;
wire n_4053;
wire n_8460;
wire n_1483;
wire n_3848;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_8836;
wire n_7959;
wire n_319;
wire n_7019;
wire n_8181;
wire n_2701;
wire n_2511;
wire n_8254;
wire n_4167;
wire n_8071;
wire n_1427;
wire n_2745;
wire n_7735;
wire n_8004;
wire n_1080;
wire n_6667;
wire n_7409;
wire n_5271;
wire n_123;
wire n_562;
wire n_6004;
wire n_5964;
wire n_2323;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_162;
wire n_7546;
wire n_4431;
wire n_5234;
wire n_2421;
wire n_1136;
wire n_6272;
wire n_4387;
wire n_2618;
wire n_6588;
wire n_3265;
wire n_2464;
wire n_128;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_5128;
wire n_9001;
wire n_2224;
wire n_2329;
wire n_1092;
wire n_441;
wire n_5467;
wire n_7296;
wire n_8013;
wire n_4299;
wire n_4890;
wire n_146;
wire n_1784;
wire n_7575;
wire n_3571;
wire n_9045;
wire n_7083;
wire n_193;
wire n_1775;
wire n_2410;
wire n_7720;
wire n_6222;
wire n_1093;
wire n_1783;
wire n_6268;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_6456;
wire n_296;
wire n_7521;
wire n_651;
wire n_3407;
wire n_5992;
wire n_217;
wire n_5313;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_7187;
wire n_3425;
wire n_215;
wire n_3894;
wire n_3127;
wire n_1831;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_6467;
wire n_5079;
wire n_6540;
wire n_6625;
wire n_1453;
wire n_6336;
wire n_6796;
wire n_2502;
wire n_3646;
wire n_5513;
wire n_5614;
wire n_497;
wire n_6541;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_3243;
wire n_2462;
wire n_1135;
wire n_2889;
wire n_8487;
wire n_4034;
wire n_4056;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_8141;
wire n_7603;
wire n_4887;
wire n_8438;
wire n_2732;
wire n_4693;
wire n_4206;
wire n_8791;
wire n_2249;
wire n_8288;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_7979;
wire n_6732;
wire n_6876;
wire n_2270;
wire n_1425;
wire n_5049;
wire n_983;
wire n_6757;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_8323;
wire n_1733;
wire n_8006;
wire n_8296;
wire n_8657;
wire n_7636;
wire n_2955;
wire n_5592;
wire n_6954;
wire n_2158;
wire n_7866;
wire n_4609;
wire n_6938;
wire n_1855;
wire n_3051;
wire n_3367;
wire n_7205;
wire n_385;
wire n_1687;
wire n_8757;
wire n_1439;
wire n_2328;
wire n_7020;
wire n_7990;
wire n_2859;
wire n_2202;
wire n_1331;
wire n_613;
wire n_736;
wire n_5278;
wire n_8596;
wire n_5157;
wire n_3314;
wire n_2100;
wire n_3525;
wire n_2993;
wire n_3016;
wire n_4754;
wire n_4647;
wire n_1134;
wire n_3688;
wire n_8590;
wire n_8720;
wire n_4003;
wire n_5708;
wire n_554;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_6298;
wire n_4894;
wire n_5474;
wire n_4113;
wire n_1889;
wire n_4760;
wire n_5649;
wire n_6421;
wire n_435;
wire n_1905;
wire n_7407;
wire n_3466;
wire n_762;
wire n_5704;
wire n_4983;
wire n_1778;
wire n_7148;
wire n_6328;
wire n_5956;
wire n_5287;
wire n_6236;
wire n_1079;
wire n_2139;
wire n_419;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_6007;
wire n_2875;
wire n_1103;
wire n_3907;
wire n_6144;
wire n_3338;
wire n_144;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_2219;
wire n_6835;
wire n_1203;
wire n_8834;
wire n_3636;
wire n_2327;
wire n_8826;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_7075;
wire n_6247;
wire n_4897;
wire n_7104;
wire n_7124;
wire n_3539;
wire n_3291;
wire n_7467;
wire n_4399;
wire n_2304;
wire n_7799;
wire n_8364;
wire n_2487;
wire n_5698;
wire n_3276;
wire n_2597;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_7513;
wire n_3572;
wire n_349;
wire n_6602;
wire n_3886;
wire n_6708;
wire n_8854;
wire n_8917;
wire n_6645;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_443;
wire n_892;
wire n_3637;
wire n_6242;
wire n_4574;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2156;
wire n_9019;
wire n_1718;
wire n_8985;
wire n_7692;
wire n_5174;
wire n_4234;
wire n_7469;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_1768;
wire n_3974;
wire n_198;
wire n_1847;
wire n_3634;
wire n_7560;
wire n_8548;
wire n_7645;
wire n_1397;
wire n_3236;
wire n_901;
wire n_2755;
wire n_3141;
wire n_923;
wire n_5096;
wire n_1841;
wire n_4660;
wire n_5241;
wire n_1623;
wire n_1015;
wire n_7082;
wire n_3112;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_4270;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_3417;
wire n_9000;
wire n_5677;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_5570;
wire n_6418;
wire n_8742;
wire n_785;
wire n_8307;
wire n_5153;
wire n_609;
wire n_4611;
wire n_8874;
wire n_5927;
wire n_7392;
wire n_7495;
wire n_5435;
wire n_2337;
wire n_1356;
wire n_3213;
wire n_4333;
wire n_127;
wire n_3820;
wire n_5200;
wire n_8706;
wire n_6400;
wire n_2607;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_6941;
wire n_1943;
wire n_5566;
wire n_7829;
wire n_3249;
wire n_1320;
wire n_7543;
wire n_8680;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_7877;
wire n_7963;
wire n_2499;
wire n_4152;
wire n_5487;
wire n_8855;
wire n_6398;
wire n_8885;
wire n_8329;
wire n_302;
wire n_5486;
wire n_137;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_8270;
wire n_4832;
wire n_2902;
wire n_5889;
wire n_3217;
wire n_7284;
wire n_1983;
wire n_7264;
wire n_5391;
wire n_1938;
wire n_7737;
wire n_6537;
wire n_8614;
wire n_2472;
wire n_7328;
wire n_3394;
wire n_1715;
wire n_3536;
wire n_8816;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_4195;
wire n_5849;
wire n_4554;
wire n_7135;
wire n_6578;
wire n_6224;
wire n_3040;
wire n_8802;
wire n_3279;
wire n_8555;
wire n_5240;
wire n_8636;
wire n_7024;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_6092;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_1692;
wire n_1084;
wire n_6614;
wire n_8508;
wire n_5912;
wire n_8667;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_3475;
wire n_3501;
wire n_374;
wire n_1705;
wire n_8121;
wire n_3905;
wire n_8207;
wire n_8035;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_3013;
wire n_921;
wire n_579;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_2257;
wire n_4927;
wire n_5574;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_7152;
wire n_2200;
wire n_650;
wire n_6165;
wire n_8320;
wire n_1940;
wire n_4548;
wire n_4862;
wire n_1405;
wire n_2376;
wire n_5469;
wire n_8766;
wire n_456;
wire n_3878;
wire n_6567;
wire n_2670;
wire n_313;
wire n_2700;
wire n_5910;
wire n_5895;
wire n_1041;
wire n_5804;
wire n_565;
wire n_3134;
wire n_5965;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_7240;
wire n_7570;
wire n_896;
wire n_4553;
wire n_3278;
wire n_7033;
wire n_2084;
wire n_4875;
wire n_7817;
wire n_5682;
wire n_5387;
wire n_654;
wire n_5557;
wire n_411;
wire n_2458;
wire n_8850;
wire n_1222;
wire n_3050;
wire n_2673;
wire n_2456;
wire n_8002;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_420;
wire n_4321;
wire n_4183;
wire n_8370;
wire n_7237;
wire n_164;
wire n_5681;
wire n_6877;
wire n_7423;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_1271;
wire n_4901;
wire n_1545;
wire n_4145;
wire n_3121;
wire n_4821;
wire n_1640;
wire n_4040;
wire n_8301;
wire n_2406;
wire n_7617;
wire n_806;
wire n_584;
wire n_2141;
wire n_7718;
wire n_5316;
wire n_244;
wire n_6940;
wire n_548;
wire n_7396;
wire n_282;
wire n_5703;
wire n_7835;
wire n_833;
wire n_523;
wire n_6320;
wire n_8126;
wire n_345;
wire n_7998;
wire n_3930;
wire n_4943;
wire n_799;
wire n_3044;
wire n_4757;
wire n_7561;
wire n_7842;
wire n_6810;
wire n_2196;
wire n_2629;
wire n_2809;
wire n_787;
wire n_2172;
wire n_6202;
wire n_4682;
wire n_5564;
wire n_5620;
wire n_7163;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_4942;
wire n_159;
wire n_1086;
wire n_5406;
wire n_2125;
wire n_8072;
wire n_2561;
wire n_8277;
wire n_7236;
wire n_652;
wire n_4604;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_5724;
wire n_7130;
wire n_1241;
wire n_7201;
wire n_3157;
wire n_4841;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_4338;
wire n_3457;
wire n_306;
wire n_3762;
wire n_8724;
wire n_5738;
wire n_3005;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_7491;
wire n_5353;
wire n_1706;
wire n_5186;
wire n_5710;
wire n_1498;
wire n_2417;
wire n_6792;
wire n_1210;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_5979;
wire n_3558;
wire n_7559;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_6044;
wire n_8867;
wire n_4326;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_5605;
wire n_2441;
wire n_3401;
wire n_3242;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_655;
wire n_4726;
wire n_7678;
wire n_1045;
wire n_5907;
wire n_786;
wire n_1559;
wire n_6045;
wire n_1872;
wire n_8132;
wire n_6731;
wire n_7526;
wire n_5040;
wire n_6063;
wire n_1325;
wire n_6504;
wire n_3761;
wire n_4315;
wire n_2888;
wire n_2923;
wire n_7004;
wire n_7821;
wire n_1727;
wire n_8308;
wire n_6154;
wire n_6943;
wire n_4301;
wire n_151;
wire n_3744;
wire n_8165;
wire n_4788;
wire n_8400;
wire n_2041;
wire n_8210;
wire n_1360;
wire n_5977;
wire n_7879;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_2484;
wire n_2126;
wire n_7696;
wire n_6003;
wire n_6684;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_6600;
wire n_2045;
wire n_817;
wire n_5451;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_6673;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_3621;
wire n_6031;
wire n_8331;
wire n_8217;
wire n_6962;
wire n_2903;
wire n_3216;
wire n_332;
wire n_3808;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_398;
wire n_4365;
wire n_6060;
wire n_1882;
wire n_7929;
wire n_3726;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_7270;
wire n_591;
wire n_3758;
wire n_8689;
wire n_5417;
wire n_6967;
wire n_2587;
wire n_7550;
wire n_3199;
wire n_680;
wire n_3339;
wire n_6853;
wire n_6742;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_6691;
wire n_8743;
wire n_7087;
wire n_8753;
wire n_1953;
wire n_6191;
wire n_4741;
wire n_6172;
wire n_3343;
wire n_2752;
wire n_8627;
wire n_4885;
wire n_751;
wire n_5432;
wire n_1399;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_7851;
wire n_6894;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_2186;
wire n_2163;
wire n_2815;
wire n_3034;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_643;
wire n_6817;
wire n_5842;
wire n_6927;
wire n_400;
wire n_337;
wire n_5814;
wire n_2814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_6215;
wire n_789;
wire n_3231;
wire n_4212;
wire n_2979;
wire n_5699;
wire n_181;
wire n_5531;
wire n_5765;
wire n_2953;
wire n_6517;
wire n_327;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_7862;
wire n_2946;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_4225;
wire n_6883;
wire n_8808;
wire n_300;
wire n_8528;
wire n_747;
wire n_8204;
wire n_2565;
wire n_5495;
wire n_1389;
wire n_535;
wire n_7100;
wire n_3583;
wire n_3860;
wire n_3851;
wire n_5655;
wire n_6393;
wire n_5064;
wire n_7825;
wire n_7119;
wire n_5610;
wire n_7212;
wire n_8154;
wire n_6966;
wire n_8889;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_6722;
wire n_1506;
wire n_119;
wire n_3473;
wire n_1652;
wire n_6035;
wire n_957;
wire n_1994;
wire n_7874;
wire n_8490;
wire n_7622;
wire n_9014;
wire n_8509;
wire n_8767;
wire n_8512;
wire n_8634;
wire n_2566;
wire n_6364;
wire n_387;
wire n_744;
wire n_971;
wire n_8635;
wire n_2702;
wire n_3241;
wire n_7102;
wire n_7420;
wire n_2906;
wire n_4342;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_1205;
wire n_6061;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_7831;
wire n_6253;
wire n_2914;
wire n_5786;
wire n_8532;
wire n_8624;
wire n_8991;
wire n_8065;
wire n_3100;
wire n_2180;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_1016;
wire n_8796;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_4373;
wire n_8518;
wire n_8919;
wire n_197;
wire n_4711;
wire n_3068;
wire n_2685;
wire n_6419;
wire n_1083;
wire n_7784;
wire n_8372;
wire n_5768;
wire n_3553;
wire n_2465;
wire n_2275;
wire n_7225;
wire n_8077;
wire n_2568;
wire n_2022;
wire n_3811;
wire n_910;
wire n_3494;
wire n_1721;
wire n_6244;
wire n_6900;
wire n_1737;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_6755;
wire n_7361;
wire n_6565;
wire n_1028;
wire n_6942;
wire n_7705;
wire n_2106;
wire n_2265;
wire n_7228;
wire n_5350;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_7932;
wire n_4409;
wire n_7509;
wire n_5872;
wire n_6862;
wire n_7058;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_708;
wire n_1973;
wire n_6840;
wire n_3181;
wire n_6338;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_1500;
wire n_6037;
wire n_7981;
wire n_3699;
wire n_854;
wire n_4913;
wire n_2312;
wire n_6266;
wire n_5874;
wire n_6488;
wire n_904;
wire n_8337;
wire n_709;
wire n_1266;
wire n_2242;
wire n_7164;
wire n_3328;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_185;
wire n_3868;
wire n_1276;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_2530;
wire n_7018;
wire n_5873;
wire n_7975;
wire n_8358;
wire n_1085;
wire n_2042;
wire n_771;
wire n_6317;
wire n_475;
wire n_924;
wire n_8199;
wire n_298;
wire n_1582;
wire n_492;
wire n_5588;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_8656;
wire n_7167;
wire n_265;
wire n_6480;
wire n_3645;
wire n_5075;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_7865;
wire n_2666;
wire n_1585;
wire n_1799;
wire n_2564;
wire n_5085;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_2035;
wire n_8881;
wire n_7844;
wire n_7134;
wire n_3422;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_406;
wire n_4104;
wire n_4845;
wire n_6875;
wire n_1770;
wire n_878;
wire n_8346;
wire n_5120;
wire n_130;
wire n_3285;
wire n_4208;
wire n_8761;
wire n_8226;
wire n_8402;
wire n_7079;
wire n_981;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_2071;
wire n_3219;
wire n_3702;
wire n_8754;
wire n_2233;
wire n_4779;
wire n_7267;
wire n_481;
wire n_3233;
wire n_4599;
wire n_997;
wire n_4437;
wire n_5222;
wire n_7316;
wire n_7850;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_7812;
wire n_1198;
wire n_7103;
wire n_4061;
wire n_8133;
wire n_7460;
wire n_6176;
wire n_2174;
wire n_436;
wire n_6367;
wire n_3881;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_2426;
wire n_2478;
wire n_7056;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_1133;
wire n_4429;
wire n_7962;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_7813;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_6080;
wire n_4865;
wire n_8182;
wire n_8387;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_7473;
wire n_7200;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_7688;
wire n_4562;
wire n_553;
wire n_3383;
wire n_8707;
wire n_4903;
wire n_3709;
wire n_3738;
wire n_7611;
wire n_6873;
wire n_4186;
wire n_8494;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_8544;
wire n_3610;
wire n_4998;
wire n_3330;
wire n_7795;
wire n_2065;
wire n_2879;
wire n_8788;
wire n_967;
wire n_4522;
wire n_7038;
wire n_2001;
wire n_7723;
wire n_4341;
wire n_679;
wire n_1629;
wire n_7404;
wire n_5368;
wire n_4263;
wire n_225;
wire n_1260;
wire n_1819;
wire n_309;
wire n_8177;
wire n_3555;
wire n_7059;
wire n_7450;
wire n_8962;
wire n_915;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_812;
wire n_6145;
wire n_1131;
wire n_3155;
wire n_6539;
wire n_6926;
wire n_1006;
wire n_3110;
wire n_7271;
wire n_1632;
wire n_7826;
wire n_5933;
wire n_257;
wire n_1888;
wire n_8993;
wire n_6204;
wire n_1311;
wire n_7076;
wire n_4780;
wire n_670;
wire n_2697;
wire n_3908;
wire n_4973;
wire n_6842;
wire n_3467;
wire n_6866;
wire n_1887;
wire n_9044;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_6451;
wire n_3039;
wire n_1226;
wire n_6514;
wire n_3740;
wire n_5996;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_640;
wire n_1322;
wire n_7105;
wire n_1958;
wire n_315;
wire n_7049;
wire n_5903;
wire n_5986;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_2579;
wire n_6345;
wire n_2105;
wire n_135;
wire n_1423;
wire n_8618;
wire n_3387;
wire n_364;
wire n_5782;
wire n_7535;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_4283;
wire n_4959;
wire n_900;
wire n_8248;
wire n_8911;
wire n_4426;
wire n_2912;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_4449;
wire n_2116;
wire n_2320;
wire n_7057;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_3002;
wire n_6957;
wire n_649;
wire n_1612;
wire n_4809;
wire n_8495;
wire n_8783;
wire n_1199;
wire n_3392;
wire n_8529;
wire n_8733;
wire n_8990;
wire n_6050;
wire n_625;
wire n_7976;
wire n_6444;
wire n_226;
wire n_7944;
wire n_7262;
wire n_212;
wire n_3773;
wire n_8647;
wire n_2003;
wire n_8574;
wire n_1038;
wire n_1581;
wire n_7016;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_6379;
wire n_798;
wire n_2324;
wire n_5563;
wire n_245;
wire n_1348;
wire n_8044;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_6719;
wire n_7178;
wire n_1380;
wire n_2847;
wire n_7506;
wire n_2557;
wire n_8551;
wire n_8330;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_6232;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_6017;
wire n_2521;
wire n_8879;
wire n_1099;
wire n_471;
wire n_424;
wire n_8052;
wire n_4578;
wire n_2211;
wire n_6362;
wire n_4777;
wire n_5720;
wire n_369;
wire n_8903;
wire n_2672;
wire n_4702;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_7142;
wire n_141;
wire n_1285;
wire n_1985;
wire n_6326;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_1172;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_4531;
wire n_3282;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_7241;
wire n_7247;
wire n_7172;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_2365;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_4029;
wire n_375;
wire n_7235;
wire n_8540;
wire n_2447;
wire n_6239;
wire n_4617;
wire n_2340;
wire n_4010;
wire n_5896;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_7588;
wire n_5650;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_7340;
wire n_6974;
wire n_5105;
wire n_1572;
wire n_4308;
wire n_5021;
wire n_3463;
wire n_8939;
wire n_428;
wire n_5263;
wire n_2510;
wire n_1954;
wire n_6713;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_822;
wire n_8468;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_5134;
wire n_7096;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_8778;
wire n_491;
wire n_3998;
wire n_7442;
wire n_1591;
wire n_3632;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_2495;
wire n_7999;
wire n_7593;
wire n_371;
wire n_6087;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_8068;
wire n_538;
wire n_3829;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_9007;
wire n_7764;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_5969;
wire n_3655;
wire n_8198;
wire n_493;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2108;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_1211;
wire n_6454;
wire n_5022;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_5670;
wire n_8557;
wire n_1280;
wire n_6041;
wire n_6918;
wire n_3296;
wire n_7350;
wire n_5276;
wire n_8012;
wire n_1445;
wire n_7672;
wire n_2551;
wire n_6664;
wire n_1526;
wire n_5047;
wire n_196;
wire n_7318;
wire n_2985;
wire n_1978;
wire n_6472;
wire n_574;
wire n_8114;
wire n_3792;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_3507;
wire n_5879;
wire n_8062;
wire n_4403;
wire n_5238;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_3531;
wire n_6375;
wire n_473;
wire n_6352;
wire n_1054;
wire n_559;
wire n_8542;
wire n_7063;
wire n_1956;
wire n_7047;
wire n_4139;
wire n_6632;
wire n_4549;
wire n_8576;
wire n_6238;
wire n_1986;
wire n_8038;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_6081;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_3603;
wire n_6724;
wire n_5429;
wire n_6545;
wire n_813;
wire n_8716;
wire n_6705;
wire n_3822;
wire n_8629;
wire n_4163;
wire n_818;
wire n_5535;
wire n_645;
wire n_7074;
wire n_3812;
wire n_3910;
wire n_8734;
wire n_2633;
wire n_6591;
wire n_2207;
wire n_7585;
wire n_4948;
wire n_5268;
wire n_6946;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_2198;
wire n_3319;
wire n_541;
wire n_2073;
wire n_2273;
wire n_6289;
wire n_7037;
wire n_3748;
wire n_3272;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_9025;
wire n_8524;
wire n_3396;
wire n_7599;
wire n_7928;
wire n_8768;
wire n_4393;
wire n_1162;
wire n_6532;
wire n_821;
wire n_4372;
wire n_1068;
wire n_7293;
wire n_982;
wire n_5640;
wire n_7600;
wire n_408;
wire n_932;
wire n_2831;
wire n_4318;
wire n_6778;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_6721;
wire n_5560;
wire n_6644;
wire n_2123;
wire n_1697;
wire n_6512;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_6108;
wire n_8258;
wire n_4918;
wire n_3824;
wire n_5067;
wire n_5744;
wire n_4013;
wire n_6703;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_354;
wire n_5841;
wire n_7614;
wire n_134;
wire n_2941;
wire n_1278;
wire n_547;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_7347;
wire n_4032;
wire n_1064;
wire n_6086;
wire n_1396;
wire n_634;
wire n_2355;
wire n_4147;
wire n_136;
wire n_4477;
wire n_3168;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_4130;
wire n_5941;
wire n_2009;
wire n_7759;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_6340;
wire n_3092;
wire n_1289;
wire n_6219;
wire n_3055;
wire n_7479;
wire n_6706;
wire n_3966;
wire n_2866;
wire n_7395;
wire n_8947;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_1703;
wire n_7078;
wire n_2580;
wire n_8188;
wire n_6761;
wire n_882;
wire n_8972;
wire n_3649;
wire n_2821;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_8510;
wire n_3384;
wire n_1950;
wire n_6811;
wire n_1563;
wire n_3419;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_7372;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_674;
wire n_3921;
wire n_6868;
wire n_8664;
wire n_922;
wire n_1335;
wire n_1927;
wire n_4838;
wire n_5970;
wire n_7174;
wire n_5202;
wire n_702;
wire n_4965;
wire n_347;
wire n_8021;
wire n_3346;
wire n_7803;
wire n_1896;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_3861;
wire n_675;
wire n_1540;
wire n_1977;
wire n_3891;
wire n_2193;
wire n_6659;
wire n_4523;
wire n_1655;
wire n_242;
wire n_6011;
wire n_1886;
wire n_4371;
wire n_6225;
wire n_2994;
wire n_5502;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_8982;
wire n_877;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_7086;
wire n_728;
wire n_3415;
wire n_1063;
wire n_6648;
wire n_4607;
wire n_7226;
wire n_6182;
wire n_7927;
wire n_9013;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_3918;
wire n_5876;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_6601;
wire n_598;
wire n_8584;
wire n_7920;
wire n_437;
wire n_7810;
wire n_8501;
wire n_4169;
wire n_8480;
wire n_697;
wire n_3271;
wire n_295;
wire n_5088;
wire n_4248;
wire n_8034;
wire n_388;
wire n_484;
wire n_7025;
wire n_8228;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_8076;
wire n_6826;
wire n_1825;
wire n_1757;
wire n_170;
wire n_1792;
wire n_5856;
wire n_8484;
wire n_1412;
wire n_2497;
wire n_3809;
wire n_3139;
wire n_8100;
wire n_4070;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_8014;
wire n_3993;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_4031;
wire n_5837;
wire n_148;
wire n_4675;
wire n_7768;
wire n_2663;
wire n_8638;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_7982;
wire n_8804;
wire n_297;
wire n_3337;
wire n_4002;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_2165;
wire n_5547;
wire n_1391;
wire n_8158;
wire n_131;
wire n_2750;
wire n_2775;
wire n_6879;
wire n_1295;
wire n_8469;
wire n_7567;
wire n_8765;
wire n_3477;
wire n_8433;
wire n_2349;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_5983;
wire n_8213;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_585;
wire n_4653;
wire n_4435;
wire n_7684;
wire n_5604;
wire n_1756;
wire n_8451;
wire n_1128;
wire n_5411;
wire n_673;
wire n_8334;
wire n_4019;
wire n_1071;
wire n_8731;
wire n_8385;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_4922;
wire n_865;
wire n_3616;
wire n_5815;
wire n_7370;
wire n_7771;
wire n_4191;
wire n_6595;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_8539;
wire n_2151;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_1839;
wire n_2341;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_2707;
wire n_6306;
wire n_6720;
wire n_6888;
wire n_826;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_1714;
wire n_8122;
wire n_718;
wire n_6095;
wire n_8432;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_542;
wire n_5311;
wire n_305;
wire n_6590;
wire n_2089;
wire n_7583;
wire n_3522;
wire n_6559;
wire n_2747;
wire n_3924;
wire n_791;
wire n_4621;
wire n_4216;
wire n_5797;
wire n_510;
wire n_4240;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_704;
wire n_2148;
wire n_7151;
wire n_4162;
wire n_5565;
wire n_8950;
wire n_2339;
wire n_2861;
wire n_1999;
wire n_2731;
wire n_622;
wire n_5520;
wire n_147;
wire n_3353;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_1838;
wire n_6287;
wire n_2638;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_1776;
wire n_1766;
wire n_7353;
wire n_2002;
wire n_2138;
wire n_7758;
wire n_4021;
wire n_2414;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_5060;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_9024;
wire n_5772;
wire n_7571;
wire n_145;
wire n_2208;
wire n_4775;
wire n_5884;
wire n_6671;
wire n_6812;
wire n_4864;
wire n_5758;
wire n_4674;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_1304;
wire n_294;
wire n_8242;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_2134;
wire n_1176;
wire n_8284;
wire n_7792;
wire n_8161;
wire n_7510;
wire n_6662;
wire n_8184;
wire n_425;
wire n_5603;
wire n_6525;
wire n_7422;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_5763;
wire n_2958;
wire n_8703;
wire n_7109;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_6128;
wire n_2489;
wire n_6029;
wire n_1087;
wire n_8822;
wire n_657;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_5924;
wire n_1505;
wire n_290;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_2610;
wire n_3129;
wire n_8476;
wire n_6702;
wire n_3620;
wire n_478;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_2520;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_3693;
wire n_446;
wire n_8545;
wire n_8736;
wire n_4497;
wire n_7749;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_8705;
wire n_526;
wire n_2251;
wire n_7508;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_4871;
wire n_8708;
wire n_293;
wire n_7574;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_1665;
wire n_4306;
wire n_154;
wire n_4224;
wire n_2127;
wire n_3341;
wire n_6005;
wire n_8872;
wire n_4453;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_6169;
wire n_8238;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_7713;
wire n_4564;
wire n_5146;
wire n_3056;
wire n_745;
wire n_2424;
wire n_3201;
wire n_3447;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_716;
wire n_1475;
wire n_1774;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_6936;
wire n_2589;
wire n_4535;
wire n_7704;
wire n_7487;
wire n_755;
wire n_8844;
wire n_6302;
wire n_527;
wire n_2442;
wire n_7641;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_7203;
wire n_1137;
wire n_7169;
wire n_7670;
wire n_3612;
wire n_4695;
wire n_6848;
wire n_2545;
wire n_8642;
wire n_3509;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_8912;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_7439;
wire n_1314;
wire n_600;
wire n_3196;
wire n_8110;
wire n_864;
wire n_5319;
wire n_2504;
wire n_2623;
wire n_9008;
wire n_399;
wire n_6343;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_8805;
wire n_1534;
wire n_6850;
wire n_5005;
wire n_8989;
wire n_6098;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_1339;
wire n_2475;
wire n_5181;
wire n_6979;
wire n_7815;
wire n_403;
wire n_7934;
wire n_723;
wire n_3144;
wire n_8111;
wire n_3244;
wire n_596;
wire n_6865;
wire n_1141;
wire n_1268;
wire n_7276;
wire n_8056;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_8739;
wire n_5043;
wire n_6747;
wire n_2025;
wire n_2357;
wire n_5583;
wire n_4654;
wire n_6433;
wire n_3640;
wire n_642;
wire n_995;
wire n_1159;
wire n_3481;
wire n_6640;
wire n_8856;
wire n_2250;
wire n_3033;
wire n_303;
wire n_6142;
wire n_5775;
wire n_6462;
wire n_7769;
wire n_2374;
wire n_416;
wire n_1681;
wire n_6034;
wire n_520;
wire n_418;
wire n_4597;
wire n_113;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_7233;
wire n_8732;
wire n_7602;
wire n_7034;
wire n_5220;
wire n_1618;
wire n_7390;
wire n_4867;
wire n_6870;
wire n_6221;
wire n_8231;
wire n_8185;
wire n_6279;
wire n_5061;
wire n_6775;
wire n_1653;
wire n_7881;
wire n_4063;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_6071;
wire n_2920;
wire n_773;
wire n_7598;
wire n_920;
wire n_1374;
wire n_8908;
wire n_2648;
wire n_3212;
wire n_8220;
wire n_6833;
wire n_6793;
wire n_1169;
wire n_6767;
wire n_6295;
wire n_1617;
wire n_3370;
wire n_3386;
wire n_335;
wire n_4721;
wire n_463;
wire n_3093;
wire n_8090;
wire n_8053;
wire n_848;
wire n_120;
wire n_274;
wire n_6385;
wire n_7426;
wire n_4247;
wire n_8137;
wire n_7045;
wire n_3169;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1806;
wire n_7984;
wire n_6788;
wire n_2023;
wire n_7014;
wire n_2720;
wire n_2204;
wire n_496;
wire n_8305;
wire n_4614;
wire n_177;
wire n_3360;
wire n_2087;
wire n_1636;
wire n_3956;
wire n_8163;
wire n_4001;
wire n_7220;
wire n_1323;
wire n_6709;
wire n_2627;
wire n_4422;
wire n_960;
wire n_6550;
wire n_6712;
wire n_7416;
wire n_6143;
wire n_778;
wire n_3004;
wire n_8841;
wire n_3870;
wire n_5177;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_6743;
wire n_4632;
wire n_1610;
wire n_3084;
wire n_5785;
wire n_2343;
wire n_793;
wire n_7465;
wire n_5967;
wire n_4546;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_6672;
wire n_2942;
wire n_4966;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_2515;
wire n_7936;
wire n_8966;
wire n_316;
wire n_6084;
wire n_1551;
wire n_4847;
wire n_4054;
wire n_8538;
wire n_7738;
wire n_2555;
wire n_3586;
wire n_3653;
wire n_8395;
wire n_5966;
wire n_2201;
wire n_725;
wire n_6634;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_8961;
wire n_7462;
wire n_4635;
wire n_368;
wire n_994;
wire n_5735;
wire n_7490;
wire n_2278;
wire n_7545;
wire n_1020;
wire n_8625;
wire n_1273;
wire n_7160;
wire n_7464;
wire n_8937;
wire n_4214;
wire n_6919;
wire n_3448;
wire n_7805;
wire n_617;
wire n_7115;
wire n_7295;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_7348;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_5360;
wire n_6681;
wire n_6104;
wire n_8179;
wire n_421;
wire n_3991;
wire n_6548;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_6993;
wire n_1095;
wire n_8511;
wire n_6973;
wire n_1270;
wire n_4405;
wire n_610;
wire n_4413;
wire n_1852;
wire n_7453;
wire n_8715;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_3670;
wire n_2381;
wire n_2052;
wire n_179;
wire n_4667;
wire n_5081;
wire n_517;
wire n_4182;
wire n_667;
wire n_3230;
wire n_8371;
wire n_8702;
wire n_8116;
wire n_1279;
wire n_1115;
wire n_7946;
wire n_8195;
wire n_1499;
wire n_8806;
wire n_504;
wire n_1409;
wire n_5877;
wire n_7681;
wire n_8845;
wire n_6018;
wire n_6619;
wire n_5189;
wire n_1503;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_8149;
wire n_3041;
wire n_4637;
wire n_2423;
wire n_8042;
wire n_603;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_8392;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_6718;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_4155;
wire n_6854;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_167;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_1216;
wire n_2716;
wire n_6032;
wire n_9047;
wire n_2452;
wire n_3650;
wire n_8968;
wire n_5446;
wire n_3010;
wire n_7855;
wire n_3043;
wire n_8050;
wire n_5224;
wire n_4590;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_2486;
wire n_3560;
wire n_3177;
wire n_4929;
wire n_5678;
wire n_6981;
wire n_122;
wire n_2220;
wire n_7065;
wire n_2577;
wire n_1262;
wire n_3238;
wire n_218;
wire n_3529;
wire n_4835;
wire n_2232;
wire n_4038;
wire n_6122;
wire n_2790;
wire n_7911;
wire n_6765;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_3784;
wire n_7330;
wire n_5437;
wire n_8883;
wire n_220;
wire n_8586;
wire n_4586;
wire n_1608;
wire n_7336;
wire n_2373;
wire n_1472;
wire n_7446;
wire n_3628;
wire n_8401;
wire n_7854;
wire n_5454;
wire n_800;
wire n_4734;
wire n_7493;
wire n_7357;
wire n_1491;
wire n_8756;
wire n_8737;
wire n_1840;
wire n_4434;
wire n_7923;
wire n_5307;
wire n_2244;
wire n_6439;
wire n_4290;
wire n_8602;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_8240;
wire n_7714;
wire n_1352;
wire n_5407;
wire n_2017;
wire n_8422;
wire n_3029;
wire n_3597;
wire n_5913;
wire n_7088;
wire n_1046;
wire n_2560;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_8878;
wire n_6406;
wire n_7440;
wire n_1102;
wire n_1963;
wire n_6945;
wire n_8112;
wire n_258;
wire n_3790;
wire n_7029;
wire n_2766;
wire n_260;
wire n_8593;
wire n_356;
wire n_3318;
wire n_4833;
wire n_5062;
wire n_6618;
wire n_6474;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_152;
wire n_4888;
wire n_7317;
wire n_776;
wire n_321;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_6000;
wire n_2782;
wire n_3977;
wire n_227;
wire n_8194;
wire n_8055;
wire n_8579;
wire n_6816;
wire n_8360;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_6425;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_7522;
wire n_6492;
wire n_2229;
wire n_8755;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_6046;
wire n_2099;
wire n_8251;
wire n_5323;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_464;
wire n_3245;
wire n_3075;
wire n_7046;
wire n_4007;
wire n_4949;
wire n_6852;
wire n_2642;
wire n_4239;
wire n_8677;
wire n_7468;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_2986;
wire n_5702;
wire n_6251;
wire n_3915;
wire n_2536;
wire n_139;
wire n_1633;
wire n_3489;
wire n_8108;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_5914;
wire n_2820;
wire n_2293;
wire n_5250;
wire n_3074;
wire n_6869;
wire n_3102;
wire n_5590;
wire n_2026;
wire n_1282;
wire n_5260;
wire n_8325;
wire n_7621;
wire n_7359;
wire n_8498;
wire n_550;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_275;
wire n_3377;
wire n_2727;
wire n_7924;
wire n_560;
wire n_4782;
wire n_1321;
wire n_7659;
wire n_2533;
wire n_569;
wire n_3530;
wire n_9005;
wire n_2869;
wire n_8875;
wire n_4378;
wire n_5349;
wire n_8274;
wire n_7153;
wire n_1235;
wire n_2759;
wire n_7836;
wire n_2361;
wire n_1292;
wire n_2266;
wire n_4876;
wire n_6146;
wire n_8504;
wire n_346;
wire n_7280;
wire n_5813;
wire n_790;
wire n_5833;
wire n_2901;
wire n_2611;
wire n_7886;
wire n_4358;
wire n_5616;
wire n_5805;
wire n_2653;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_299;
wire n_1248;
wire n_902;
wire n_2189;
wire n_2246;
wire n_6631;
wire n_4469;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_431;
wire n_5816;
wire n_3156;
wire n_8927;
wire n_672;
wire n_6228;
wire n_6711;
wire n_1941;
wire n_3483;
wire n_5416;
wire n_8946;
wire n_706;
wire n_1794;
wire n_1236;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_8017;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_8474;
wire n_3524;
wire n_7275;
wire n_8232;
wire n_489;
wire n_2885;
wire n_8795;
wire n_7195;
wire n_6102;
wire n_636;
wire n_8904;
wire n_6274;
wire n_8838;
wire n_3097;
wire n_7007;
wire n_660;
wire n_2062;
wire n_7070;
wire n_4539;
wire n_2975;
wire n_8382;
wire n_4421;
wire n_6072;
wire n_7610;
wire n_2839;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_2070;
wire n_7259;
wire n_1607;
wire n_1454;
wire n_6353;
wire n_4953;
wire n_6992;
wire n_2944;
wire n_2348;
wire n_8128;
wire n_6818;
wire n_3831;
wire n_869;
wire n_1154;
wire n_646;
wire n_528;
wire n_391;
wire n_1329;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5830;
wire n_5932;
wire n_3589;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_7539;
wire n_841;
wire n_1476;
wire n_3391;
wire n_8794;
wire n_7616;
wire n_508;
wire n_1800;
wire n_8189;
wire n_6498;
wire n_1463;
wire n_8481;
wire n_3458;
wire n_7775;
wire n_4505;
wire n_3190;
wire n_1562;
wire n_7930;
wire n_5558;
wire n_1826;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_8205;
wire n_5051;
wire n_5587;
wire n_6976;
wire n_6304;
wire n_5236;
wire n_853;
wire n_7640;
wire n_875;
wire n_5012;
wire n_1678;
wire n_661;
wire n_6864;
wire n_7969;
wire n_8605;
wire n_3787;
wire n_1256;
wire n_7548;
wire n_3585;
wire n_3565;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_5025;
wire n_933;
wire n_6998;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_3135;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_8000;
wire n_1217;
wire n_7197;
wire n_5645;
wire n_3990;
wire n_7393;
wire n_6917;
wire n_6937;
wire n_7591;
wire n_310;
wire n_1628;
wire n_5766;
wire n_2109;
wire n_7727;
wire n_7358;
wire n_988;
wire n_2796;
wire n_7324;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_4534;
wire n_1536;
wire n_6301;
wire n_1204;
wire n_1132;
wire n_6929;
wire n_233;
wire n_1327;
wire n_8719;
wire n_955;
wire n_8045;
wire n_7729;
wire n_246;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_8209;
wire n_769;
wire n_2380;
wire n_4786;
wire n_7565;
wire n_1120;
wire n_6699;
wire n_555;
wire n_4579;
wire n_7291;
wire n_7631;
wire n_669;
wire n_8784;
wire n_2290;
wire n_7382;
wire n_4811;
wire n_2048;
wire n_176;
wire n_114;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_2005;
wire n_4857;
wire n_7437;
wire n_6677;
wire n_3432;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_7618;
wire n_4282;
wire n_1196;
wire n_3493;
wire n_8769;
wire n_6764;
wire n_8575;
wire n_863;
wire n_3774;
wire n_5733;
wire n_6780;
wire n_8815;
wire n_2910;
wire n_6620;
wire n_6597;
wire n_748;
wire n_3268;
wire n_1785;
wire n_1147;
wire n_1754;
wire n_3057;
wire n_3701;
wire n_5148;
wire n_8261;
wire n_2584;
wire n_7673;
wire n_1812;
wire n_6830;
wire n_866;
wire n_8655;
wire n_7282;
wire n_2287;
wire n_452;
wire n_6586;
wire n_6333;
wire n_7139;
wire n_8745;
wire n_5791;
wire n_5727;
wire n_8086;
wire n_761;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_2492;
wire n_7953;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_5657;
wire n_174;
wire n_1173;
wire n_8901;
wire n_8695;
wire n_4974;
wire n_5975;
wire n_4911;
wire n_8173;
wire n_4436;
wire n_8363;
wire n_5119;
wire n_4569;
wire n_1174;
wire n_8665;
wire n_6510;
wire n_8282;
wire n_3334;
wire n_5938;
wire n_6237;
wire n_5602;
wire n_647;
wire n_5097;
wire n_844;
wire n_4985;
wire n_7751;
wire n_2117;
wire n_2234;
wire n_3823;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_7581;
wire n_888;
wire n_6360;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_236;
wire n_4858;
wire n_4678;
wire n_2649;
wire n_3556;
wire n_3836;
wire n_5579;
wire n_8835;
wire n_414;
wire n_1922;
wire n_5750;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_1215;
wire n_839;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_8493;
wire n_7346;
wire n_779;
wire n_1537;
wire n_2205;
wire n_4243;
wire n_7579;
wire n_4025;
wire n_7428;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_4059;
wire n_1509;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_8870;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_4313;
wire n_3309;
wire n_4142;
wire n_3671;
wire n_2015;
wire n_6475;
wire n_7283;
wire n_3982;
wire n_7699;
wire n_7015;
wire n_8507;
wire n_6314;
wire n_8415;
wire n_6103;
wire n_2609;
wire n_1161;
wire n_7249;
wire n_5546;
wire n_3796;
wire n_232;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_3840;
wire n_3461;
wire n_6680;
wire n_3408;
wire n_7985;
wire n_4246;
wire n_7432;
wire n_8365;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_228;
wire n_8893;
wire n_1525;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_4244;
wire n_2147;
wire n_592;
wire n_2503;
wire n_4049;
wire n_6752;
wire n_1156;
wire n_8976;
wire n_6426;
wire n_2600;
wire n_984;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_8502;
wire n_8244;
wire n_7612;
wire n_8156;
wire n_7494;
wire n_132;
wire n_868;
wire n_4353;
wire n_735;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_4787;
wire n_7736;
wire n_5633;
wire n_469;
wire n_1218;
wire n_5664;
wire n_7589;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7177;
wire n_7814;
wire n_357;
wire n_8660;
wire n_2429;
wire n_8479;
wire n_985;
wire n_2440;
wire n_6054;
wire n_3521;
wire n_8723;
wire n_802;
wire n_561;
wire n_8606;
wire n_980;
wire n_2681;
wire n_7843;
wire n_6235;
wire n_8235;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_116;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_6496;
wire n_3066;
wire n_7756;
wire n_2844;
wire n_8342;
wire n_8940;
wire n_2303;
wire n_1619;
wire n_2285;
wire n_8448;
wire n_5280;
wire n_8472;
wire n_7700;
wire n_4451;
wire n_4332;
wire n_810;
wire n_7555;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_3976;
wire n_7988;
wire n_8658;
wire n_3563;
wire n_6513;
wire n_7500;
wire n_2367;
wire n_201;
wire n_3198;
wire n_3495;
wire n_1034;
wire n_5925;
wire n_2909;
wire n_754;
wire n_6138;
wire n_5369;
wire n_8061;
wire n_8866;
wire n_975;
wire n_5730;
wire n_5576;
wire n_3359;
wire n_5272;
wire n_6330;
wire n_467;
wire n_3187;
wire n_3218;
wire n_8457;
wire n_6802;
wire n_582;
wire n_861;
wire n_6909;
wire n_7157;
wire n_6908;
wire n_857;
wire n_8237;
wire n_7411;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4336;
wire n_4201;
wire n_7266;
wire n_2221;
wire n_8046;
wire n_588;
wire n_7871;
wire n_5646;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_6477;
wire n_6263;
wire n_8073;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_6490;
wire n_2709;
wire n_8652;
wire n_8821;
wire n_534;
wire n_7198;
wire n_1578;
wire n_8335;
wire n_1861;
wire n_3955;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_5214;
wire n_203;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_207;
wire n_2079;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_8663;
wire n_3433;
wire n_4463;
wire n_7794;
wire n_205;
wire n_2185;
wire n_6038;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_2774;
wire n_3162;
wire n_1274;
wire n_8309;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_8945;
wire n_6605;
wire n_5032;
wire n_8964;
wire n_1899;
wire n_9032;
wire n_6313;
wire n_784;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_3965;
wire n_7145;
wire n_9041;
wire n_5859;
wire n_5380;
wire n_4500;
wire n_5065;
wire n_862;
wire n_5776;
wire n_8166;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_5644;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_2091;
wire n_8960;
wire n_5920;
wire n_2991;
wire n_5030;
wire n_4194;
wire n_7994;
wire n_1449;
wire n_4703;
wire n_8443;
wire n_361;
wire n_7349;
wire n_8215;
wire n_7715;
wire n_2419;
wire n_6180;
wire n_8683;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_2677;
wire n_3182;
wire n_5756;
wire n_3283;
wire n_5527;
wire n_6476;
wire n_8037;
wire n_1742;
wire n_4030;

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_14),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_37),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g118 ( 
.A(n_68),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_6),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_52),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_16),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_36),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_31),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_45),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

BUFx10_ASAP7_75t_L g128 ( 
.A(n_53),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_19),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_35),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_34),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_26),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_41),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_29),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_60),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_43),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_80),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_8),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_34),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_13),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_96),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_22),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_15),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_5),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_19),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_106),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_45),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_48),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_105),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_47),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_23),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_40),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_42),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_47),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_29),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_33),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_16),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_98),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_94),
.Y(n_168)
);

BUFx2_ASAP7_75t_SL g169 ( 
.A(n_59),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_43),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_30),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_51),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_56),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_102),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_76),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_17),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_55),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_17),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_35),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_42),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_0),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_0),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_41),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_2),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_13),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_8),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_4),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_20),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_71),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_111),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_11),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_95),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_85),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_14),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_52),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_75),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_25),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_90),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_77),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_33),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_38),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_1),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_57),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_2),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_93),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_48),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_64),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_74),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_50),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_39),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_51),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_10),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_78),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_3),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_49),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_113),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_135),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_117),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_117),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_156),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_116),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_128),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_137),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_139),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_153),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_143),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_115),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_123),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_117),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_117),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_117),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_194),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_117),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_117),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_140),
.B(n_1),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_117),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_162),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_235),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_228),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_230),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_228),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_231),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_225),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_236),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_237),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_240),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_233),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_226),
.B(n_131),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_233),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_240),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_R g284 ( 
.A(n_241),
.B(n_120),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_226),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_241),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_229),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_229),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_235),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_288),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_222),
.B1(n_205),
.B2(n_167),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_256),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_258),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_265),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_251),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_270),
.B(n_272),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_158),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_259),
.A2(n_244),
.B1(n_246),
.B2(n_129),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_276),
.A2(n_159),
.B1(n_141),
.B2(n_138),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_254),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_260),
.B(n_254),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_288),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_263),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_264),
.B(n_232),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_153),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_255),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_269),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_255),
.Y(n_324)
);

AND2x4_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_158),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_261),
.Y(n_326)
);

OAI21x1_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_213),
.B(n_249),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_284),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_288),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_267),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

BUFx8_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_273),
.B(n_131),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_285),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_285),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_289),
.A2(n_292),
.B(n_291),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g340 ( 
.A(n_289),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_287),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

OAI21x1_ASAP7_75t_L g346 ( 
.A1(n_257),
.A2(n_213),
.B(n_249),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_232),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_286),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_280),
.B(n_232),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_282),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_288),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_288),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_256),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_274),
.B(n_238),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_270),
.B(n_227),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_281),
.B(n_244),
.Y(n_357)
);

AND2x6_ASAP7_75t_L g358 ( 
.A(n_256),
.B(n_153),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_256),
.Y(n_359)
);

BUFx8_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_259),
.A2(n_246),
.B1(n_122),
.B2(n_129),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_288),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_256),
.A2(n_121),
.B(n_114),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_284),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_270),
.B(n_234),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_281),
.A2(n_130),
.B1(n_125),
.B2(n_124),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_256),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_274),
.B(n_238),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_274),
.B(n_238),
.Y(n_371)
);

BUFx8_ASAP7_75t_L g372 ( 
.A(n_274),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_288),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_259),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_256),
.B(n_171),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_256),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_270),
.Y(n_377)
);

OAI22x1_ASAP7_75t_R g378 ( 
.A1(n_259),
.A2(n_170),
.B1(n_164),
.B2(n_160),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_274),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_281),
.B(n_249),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_256),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_265),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_270),
.B(n_128),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_256),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_274),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_256),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_256),
.Y(n_387)
);

AOI22x1_ASAP7_75t_SL g388 ( 
.A1(n_259),
.A2(n_145),
.B1(n_202),
.B2(n_190),
.Y(n_388)
);

OA21x2_ASAP7_75t_L g389 ( 
.A1(n_256),
.A2(n_179),
.B(n_114),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_256),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_256),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_256),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_288),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_256),
.A2(n_147),
.B(n_127),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_270),
.B(n_234),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_256),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_256),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_256),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_256),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_256),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_256),
.B(n_171),
.Y(n_402)
);

CKINVDCx6p67_ASAP7_75t_R g403 ( 
.A(n_257),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_274),
.B(n_238),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_270),
.B(n_121),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_256),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_274),
.B(n_253),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_259),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_270),
.B(n_127),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_256),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_270),
.B(n_128),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

AO22x2_ASAP7_75t_L g413 ( 
.A1(n_388),
.A2(n_140),
.B1(n_223),
.B2(n_219),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_377),
.Y(n_414)
);

AO22x2_ASAP7_75t_L g415 ( 
.A1(n_388),
.A2(n_182),
.B1(n_223),
.B2(n_219),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_163),
.B1(n_221),
.B2(n_168),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_336),
.A2(n_196),
.B1(n_174),
.B2(n_175),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_336),
.A2(n_147),
.B1(n_179),
.B2(n_200),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_296),
.A2(n_136),
.B1(n_220),
.B2(n_218),
.Y(n_419)
);

NAND3x1_ASAP7_75t_L g420 ( 
.A(n_296),
.B(n_142),
.C(n_216),
.Y(n_420)
);

AO22x2_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_142),
.B1(n_216),
.B2(n_119),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_356),
.B(n_150),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_357),
.A2(n_197),
.B1(n_217),
.B2(n_178),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_332),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_362),
.A2(n_133),
.B1(n_215),
.B2(n_126),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_346),
.A2(n_154),
.B1(n_192),
.B2(n_165),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_346),
.A2(n_193),
.B1(n_203),
.B2(n_176),
.Y(n_427)
);

NOR2x1p5_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_157),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_L g429 ( 
.A1(n_367),
.A2(n_200),
.B1(n_214),
.B2(n_161),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g430 ( 
.A1(n_411),
.A2(n_182),
.B1(n_122),
.B2(n_212),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_356),
.B(n_157),
.Y(n_431)
);

OA22x2_ASAP7_75t_L g432 ( 
.A1(n_367),
.A2(n_186),
.B1(n_184),
.B2(n_183),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_333),
.B(n_149),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_298),
.Y(n_434)
);

OAI22xp33_ASAP7_75t_L g435 ( 
.A1(n_306),
.A2(n_118),
.B1(n_161),
.B2(n_214),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_339),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_332),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_346),
.A2(n_211),
.B1(n_209),
.B2(n_152),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_356),
.B(n_155),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g440 ( 
.A1(n_304),
.A2(n_201),
.B1(n_118),
.B2(n_169),
.Y(n_440)
);

OAI22xp33_ASAP7_75t_L g441 ( 
.A1(n_306),
.A2(n_180),
.B1(n_189),
.B2(n_191),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_298),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_304),
.A2(n_169),
.B1(n_128),
.B2(n_162),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_303),
.Y(n_444)
);

AO22x2_ASAP7_75t_L g445 ( 
.A1(n_344),
.A2(n_173),
.B1(n_172),
.B2(n_166),
.Y(n_445)
);

OR2x2_ASAP7_75t_L g446 ( 
.A(n_377),
.B(n_177),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_379),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_362),
.A2(n_208),
.B1(n_199),
.B2(n_134),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_366),
.B(n_119),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_332),
.Y(n_450)
);

OR2x6_ASAP7_75t_L g451 ( 
.A(n_343),
.B(n_132),
.Y(n_451)
);

AO22x2_ASAP7_75t_L g452 ( 
.A1(n_344),
.A2(n_134),
.B1(n_132),
.B2(n_144),
.Y(n_452)
);

OR2x6_ASAP7_75t_L g453 ( 
.A(n_343),
.B(n_144),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_366),
.B(n_148),
.Y(n_454)
);

OAI22xp33_ASAP7_75t_SL g455 ( 
.A1(n_328),
.A2(n_148),
.B1(n_212),
.B2(n_166),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_343),
.B(n_198),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_366),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_332),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_395),
.B(n_195),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_395),
.B(n_195),
.Y(n_460)
);

OAI22xp33_ASAP7_75t_L g461 ( 
.A1(n_343),
.A2(n_180),
.B1(n_172),
.B2(n_173),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_395),
.B(n_204),
.Y(n_462)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_326),
.Y(n_463)
);

BUFx10_ASAP7_75t_L g464 ( 
.A(n_301),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_405),
.B(n_204),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_315),
.B(n_183),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_405),
.B(n_206),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_300),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_206),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_409),
.B(n_328),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_409),
.B(n_365),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_340),
.B(n_162),
.Y(n_472)
);

BUFx10_ASAP7_75t_L g473 ( 
.A(n_382),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_304),
.A2(n_162),
.B1(n_207),
.B2(n_210),
.Y(n_474)
);

AO22x2_ASAP7_75t_L g475 ( 
.A1(n_409),
.A2(n_210),
.B1(n_207),
.B2(n_198),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_365),
.B(n_347),
.Y(n_476)
);

OAI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_304),
.A2(n_186),
.B1(n_184),
.B2(n_162),
.Y(n_477)
);

AO22x2_ASAP7_75t_L g478 ( 
.A1(n_348),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_350),
.B(n_162),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_304),
.A2(n_162),
.B1(n_252),
.B2(n_238),
.Y(n_480)
);

AO22x2_ASAP7_75t_L g481 ( 
.A1(n_348),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_305),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_325),
.A2(n_253),
.B1(n_252),
.B2(n_238),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_332),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_325),
.A2(n_253),
.B1(n_252),
.B2(n_238),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_300),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_374),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_325),
.A2(n_253),
.B1(n_252),
.B2(n_110),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_313),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_343),
.A2(n_253),
.B1(n_252),
.B2(n_20),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_313),
.Y(n_491)
);

OR2x2_ASAP7_75t_L g492 ( 
.A(n_350),
.B(n_12),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_325),
.A2(n_12),
.B1(n_18),
.B2(n_21),
.Y(n_493)
);

AO22x2_ASAP7_75t_L g494 ( 
.A1(n_348),
.A2(n_18),
.B1(n_21),
.B2(n_22),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_339),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_340),
.B(n_253),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_318),
.Y(n_497)
);

OAI22xp33_ASAP7_75t_L g498 ( 
.A1(n_343),
.A2(n_253),
.B1(n_252),
.B2(n_25),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_408),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_325),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_375),
.A2(n_253),
.B1(n_252),
.B2(n_63),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_350),
.B(n_252),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_375),
.A2(n_61),
.B1(n_104),
.B2(n_101),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_318),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_332),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_347),
.B(n_24),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_315),
.B(n_54),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_297),
.Y(n_508)
);

OR2x6_ASAP7_75t_L g509 ( 
.A(n_343),
.B(n_27),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_375),
.A2(n_402),
.B1(n_379),
.B2(n_385),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_297),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_320),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_320),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_347),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_375),
.A2(n_62),
.B1(n_100),
.B2(n_99),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_375),
.A2(n_107),
.B1(n_92),
.B2(n_89),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_321),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_315),
.B(n_27),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_379),
.B(n_88),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_297),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_345),
.B(n_28),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_402),
.A2(n_82),
.B1(n_81),
.B2(n_70),
.Y(n_522)
);

OAI22xp33_ASAP7_75t_L g523 ( 
.A1(n_345),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_402),
.A2(n_32),
.B1(n_36),
.B2(n_37),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_321),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_385),
.B(n_65),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_345),
.A2(n_354),
.B1(n_400),
.B2(n_399),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_305),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_SL g529 ( 
.A1(n_402),
.A2(n_46),
.B1(n_49),
.B2(n_334),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_402),
.A2(n_46),
.B1(n_385),
.B2(n_340),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_345),
.B(n_403),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_334),
.A2(n_410),
.B1(n_400),
.B2(n_399),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_354),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_369),
.A2(n_410),
.B1(n_392),
.B2(n_381),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_351),
.A2(n_349),
.B1(n_378),
.B2(n_345),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_369),
.A2(n_381),
.B1(n_392),
.B2(n_390),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_386),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_386),
.Y(n_538)
);

BUFx10_ASAP7_75t_L g539 ( 
.A(n_345),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_387),
.A2(n_390),
.B1(n_391),
.B2(n_331),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_345),
.B(n_349),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_378),
.A2(n_349),
.B1(n_387),
.B2(n_391),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_331),
.A2(n_302),
.B1(n_307),
.B2(n_324),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_299),
.Y(n_544)
);

OA22x2_ASAP7_75t_L g545 ( 
.A1(n_351),
.A2(n_327),
.B1(n_403),
.B2(n_384),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_331),
.A2(n_372),
.B1(n_360),
.B2(n_384),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_299),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_299),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_309),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_309),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_331),
.A2(n_372),
.B1(n_360),
.B2(n_319),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_309),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_360),
.A2(n_372),
.B1(n_319),
.B2(n_322),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_312),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_312),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_335),
.A2(n_364),
.B1(n_394),
.B2(n_389),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_312),
.B(n_406),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_314),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_314),
.B(n_397),
.Y(n_559)
);

INVxp33_ASAP7_75t_L g560 ( 
.A(n_364),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_SL g561 ( 
.A1(n_308),
.A2(n_324),
.B1(n_317),
.B2(n_307),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_302),
.B(n_308),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_317),
.B(n_359),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_314),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_319),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_364),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_360),
.A2(n_372),
.B1(n_361),
.B2(n_406),
.Y(n_567)
);

OAI22xp33_ASAP7_75t_L g568 ( 
.A1(n_322),
.A2(n_361),
.B1(n_406),
.B2(n_398),
.Y(n_568)
);

OAI22xp33_ASAP7_75t_L g569 ( 
.A1(n_322),
.A2(n_342),
.B1(n_384),
.B2(n_361),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_329),
.Y(n_570)
);

OAI22xp33_ASAP7_75t_L g571 ( 
.A1(n_329),
.A2(n_341),
.B1(n_342),
.B2(n_359),
.Y(n_571)
);

AO22x2_ASAP7_75t_L g572 ( 
.A1(n_335),
.A2(n_329),
.B1(n_398),
.B2(n_397),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_337),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_364),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_364),
.A2(n_389),
.B1(n_394),
.B2(n_335),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_337),
.B(n_342),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_337),
.A2(n_359),
.B1(n_341),
.B2(n_398),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_335),
.A2(n_376),
.B1(n_341),
.B2(n_397),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_338),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_316),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_389),
.A2(n_394),
.B1(n_339),
.B2(n_376),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_360),
.A2(n_372),
.B1(n_396),
.B2(n_376),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_338),
.A2(n_396),
.B1(n_339),
.B2(n_327),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_338),
.Y(n_584)
);

NAND2x1p5_ASAP7_75t_L g585 ( 
.A(n_339),
.B(n_327),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_396),
.B(n_363),
.Y(n_586)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_389),
.B(n_394),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_389),
.A2(n_394),
.B1(n_404),
.B2(n_407),
.Y(n_588)
);

AO22x2_ASAP7_75t_L g589 ( 
.A1(n_355),
.A2(n_407),
.B1(n_404),
.B2(n_371),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_355),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_310),
.A2(n_401),
.B1(n_373),
.B2(n_363),
.Y(n_591)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_370),
.B(n_371),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_310),
.B(n_401),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_310),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_310),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_352),
.B(n_401),
.Y(n_596)
);

INVx8_ASAP7_75t_L g597 ( 
.A(n_316),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_316),
.Y(n_598)
);

BUFx10_ASAP7_75t_L g599 ( 
.A(n_316),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_352),
.B(n_401),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_352),
.A2(n_373),
.B1(n_363),
.B2(n_370),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_352),
.A2(n_373),
.B1(n_363),
.B2(n_316),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_373),
.A2(n_358),
.B1(n_316),
.B2(n_311),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_295),
.B(n_311),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_295),
.A2(n_311),
.B1(n_368),
.B2(n_323),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_316),
.A2(n_358),
.B1(n_311),
.B2(n_323),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_R g607 ( 
.A1(n_316),
.A2(n_358),
.B1(n_311),
.B2(n_323),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_316),
.A2(n_358),
.B1(n_311),
.B2(n_323),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_295),
.B(n_311),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_295),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_295),
.B(n_323),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_393),
.A2(n_358),
.B1(n_323),
.B2(n_330),
.Y(n_612)
);

AND2x2_ASAP7_75t_SL g613 ( 
.A(n_295),
.B(n_323),
.Y(n_613)
);

OAI22xp33_ASAP7_75t_R g614 ( 
.A1(n_358),
.A2(n_295),
.B1(n_330),
.B2(n_353),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_330),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_358),
.A2(n_330),
.B1(n_353),
.B2(n_368),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_330),
.B(n_353),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_330),
.A2(n_353),
.B1(n_368),
.B2(n_393),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_330),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_358),
.A2(n_353),
.B1(n_368),
.B2(n_393),
.Y(n_620)
);

OAI22xp33_ASAP7_75t_L g621 ( 
.A1(n_353),
.A2(n_368),
.B1(n_393),
.B2(n_358),
.Y(n_621)
);

AO22x2_ASAP7_75t_L g622 ( 
.A1(n_353),
.A2(n_388),
.B1(n_336),
.B2(n_246),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_368),
.A2(n_380),
.B1(n_336),
.B2(n_357),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_368),
.A2(n_228),
.B1(n_261),
.B2(n_259),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_393),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_393),
.B(n_356),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_393),
.A2(n_388),
.B1(n_336),
.B2(n_246),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_339),
.Y(n_629)
);

AND2x2_ASAP7_75t_SL g630 ( 
.A(n_336),
.B(n_296),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_298),
.Y(n_632)
);

OAI22xp33_ASAP7_75t_L g633 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_298),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_356),
.B(n_366),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_L g636 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_636)
);

OAI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_336),
.A2(n_380),
.B1(n_235),
.B2(n_296),
.Y(n_637)
);

OA22x2_ASAP7_75t_L g638 ( 
.A1(n_367),
.A2(n_296),
.B1(n_362),
.B2(n_306),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_332),
.Y(n_640)
);

OAI22xp33_ASAP7_75t_L g641 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_641)
);

NOR2x1p5_ASAP7_75t_L g642 ( 
.A(n_403),
.B(n_233),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_332),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_L g644 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_644)
);

AO22x2_ASAP7_75t_L g645 ( 
.A1(n_388),
.A2(n_336),
.B1(n_246),
.B2(n_244),
.Y(n_645)
);

OA22x2_ASAP7_75t_L g646 ( 
.A1(n_367),
.A2(n_296),
.B1(n_362),
.B2(n_306),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_298),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_356),
.B(n_366),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_339),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_332),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_340),
.B(n_380),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_332),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_298),
.Y(n_654)
);

AO22x2_ASAP7_75t_L g655 ( 
.A1(n_388),
.A2(n_336),
.B1(n_246),
.B2(n_244),
.Y(n_655)
);

AO22x2_ASAP7_75t_L g656 ( 
.A1(n_388),
.A2(n_336),
.B1(n_246),
.B2(n_244),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_343),
.B(n_345),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_339),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_377),
.Y(n_660)
);

AO22x2_ASAP7_75t_L g661 ( 
.A1(n_388),
.A2(n_336),
.B1(n_246),
.B2(n_244),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_332),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_663)
);

OAI22xp33_ASAP7_75t_SL g664 ( 
.A1(n_336),
.A2(n_380),
.B1(n_235),
.B2(n_296),
.Y(n_664)
);

AO22x2_ASAP7_75t_L g665 ( 
.A1(n_388),
.A2(n_336),
.B1(n_246),
.B2(n_244),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_332),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_356),
.B(n_366),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_298),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_343),
.B(n_345),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_298),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_332),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_377),
.Y(n_674)
);

OAI22xp33_ASAP7_75t_SL g675 ( 
.A1(n_336),
.A2(n_380),
.B1(n_235),
.B2(n_296),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_326),
.Y(n_676)
);

OAI22xp33_ASAP7_75t_SL g677 ( 
.A1(n_336),
.A2(n_380),
.B1(n_235),
.B2(n_296),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_332),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_380),
.A2(n_336),
.B1(n_357),
.B2(n_346),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_336),
.A2(n_367),
.B1(n_380),
.B2(n_296),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_332),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_633),
.Y(n_682)
);

INVx4_ASAP7_75t_L g683 ( 
.A(n_613),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_544),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_623),
.B(n_636),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_557),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_576),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_652),
.B(n_562),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_544),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_547),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_609),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_635),
.B(n_648),
.Y(n_692)
);

AND2x6_ASAP7_75t_L g693 ( 
.A(n_436),
.B(n_495),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_547),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_548),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_463),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_434),
.B(n_468),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_641),
.B(n_644),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_650),
.B(n_680),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_SL g700 ( 
.A(n_630),
.B(n_464),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_434),
.B(n_468),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_657),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_638),
.A2(n_646),
.B1(n_545),
.B2(n_507),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_657),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_548),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_L g706 ( 
.A(n_615),
.B(n_531),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_628),
.B(n_639),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_550),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_614),
.A2(n_659),
.B1(n_669),
.B2(n_663),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_507),
.A2(n_518),
.B1(n_479),
.B2(n_673),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_550),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_679),
.B(n_470),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_552),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_609),
.Y(n_714)
);

BUFx4f_ASAP7_75t_L g715 ( 
.A(n_670),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_497),
.B(n_504),
.Y(n_716)
);

XOR2xp5_ASAP7_75t_L g717 ( 
.A(n_624),
.B(n_433),
.Y(n_717)
);

NAND2xp33_ASAP7_75t_SL g718 ( 
.A(n_535),
.B(n_471),
.Y(n_718)
);

INVx4_ASAP7_75t_SL g719 ( 
.A(n_581),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_552),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_554),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_554),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_614),
.A2(n_575),
.B1(n_592),
.B2(n_667),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_497),
.B(n_504),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_555),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_539),
.B(n_457),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_555),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_573),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_414),
.B(n_674),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_512),
.B(n_513),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_573),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_SL g732 ( 
.A(n_464),
.B(n_473),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_660),
.B(n_476),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_429),
.A2(n_502),
.B1(n_466),
.B2(n_521),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_600),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_539),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_579),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_579),
.Y(n_738)
);

CKINVDCx11_ASAP7_75t_R g739 ( 
.A(n_473),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_559),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_466),
.A2(n_477),
.B1(n_435),
.B2(n_563),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_559),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_512),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_513),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_517),
.B(n_525),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_525),
.B(n_533),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_533),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_SL g749 ( 
.A(n_492),
.B(n_506),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_537),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_514),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_537),
.Y(n_752)
);

AOI22xp33_ASAP7_75t_SL g753 ( 
.A1(n_637),
.A2(n_664),
.B1(n_675),
.B2(n_677),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_465),
.B(n_467),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_538),
.B(n_632),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_538),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_632),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_446),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_670),
.Y(n_759)
);

INVx3_ASAP7_75t_L g760 ( 
.A(n_600),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_519),
.B(n_526),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_604),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_634),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_634),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_469),
.B(n_459),
.Y(n_765)
);

INVxp67_ASAP7_75t_R g766 ( 
.A(n_626),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_668),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_611),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_519),
.B(n_526),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_668),
.B(n_671),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_671),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_530),
.A2(n_523),
.B1(n_540),
.B2(n_510),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_436),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_508),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_495),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_442),
.B(n_486),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_478),
.A2(n_481),
.B1(n_494),
.B2(n_574),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_617),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_629),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_444),
.B(n_423),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_629),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_489),
.B(n_491),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_532),
.B(n_536),
.C(n_647),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_654),
.B(n_590),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_451),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_649),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_541),
.B(n_553),
.Y(n_787)
);

BUFx4f_ASAP7_75t_L g788 ( 
.A(n_541),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_590),
.B(n_534),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_511),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_561),
.B(n_543),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_444),
.B(n_417),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_416),
.B(n_439),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_605),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_649),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_567),
.B(n_582),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_527),
.B(n_418),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_658),
.Y(n_798)
);

BUFx10_ASAP7_75t_L g799 ( 
.A(n_642),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_520),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_549),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_SL g802 ( 
.A(n_428),
.B(n_460),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_419),
.B(n_449),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_454),
.B(n_658),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_558),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_564),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_412),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_676),
.B(n_451),
.Y(n_808)
);

AOI22xp5_ASAP7_75t_L g809 ( 
.A1(n_589),
.A2(n_474),
.B1(n_607),
.B2(n_432),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_426),
.B(n_427),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_565),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_487),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_570),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_584),
.Y(n_814)
);

OR2x2_ASAP7_75t_L g815 ( 
.A(n_453),
.B(n_456),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_422),
.B(n_431),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_441),
.A2(n_421),
.B1(n_430),
.B2(n_589),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_421),
.A2(n_430),
.B1(n_560),
.B2(n_456),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_453),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_577),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_586),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_572),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_568),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_607),
.A2(n_622),
.B1(n_448),
.B2(n_475),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_569),
.Y(n_825)
);

AND3x2_ASAP7_75t_L g826 ( 
.A(n_499),
.B(n_462),
.C(n_528),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_509),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_572),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_475),
.B(n_445),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_438),
.B(n_546),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_585),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_455),
.B(n_425),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_597),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_447),
.B(n_463),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_440),
.B(n_509),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_571),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_566),
.B(n_472),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_424),
.B(n_681),
.Y(n_838)
);

BUFx6f_ASAP7_75t_SL g839 ( 
.A(n_580),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_443),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_594),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_595),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_551),
.B(n_529),
.Y(n_843)
);

INVx8_ASAP7_75t_L g844 ( 
.A(n_597),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_490),
.A2(n_498),
.B1(n_461),
.B2(n_587),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_437),
.B(n_678),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_610),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_608),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_610),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_478),
.A2(n_481),
.B1(n_494),
.B2(n_640),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_619),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_450),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_619),
.B(n_556),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_458),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_484),
.B(n_672),
.Y(n_855)
);

AND2x6_ASAP7_75t_L g856 ( 
.A(n_583),
.B(n_501),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_505),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_643),
.B(n_666),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_651),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_653),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_662),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_608),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_601),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_591),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_496),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_593),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_596),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_482),
.B(n_524),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_578),
.A2(n_588),
.B1(n_622),
.B2(n_515),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_618),
.B(n_602),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_480),
.Y(n_871)
);

AO22x2_ASAP7_75t_L g872 ( 
.A1(n_578),
.A2(n_420),
.B1(n_627),
.B2(n_445),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_616),
.Y(n_873)
);

BUFx10_ASAP7_75t_L g874 ( 
.A(n_625),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_612),
.B(n_500),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_625),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_483),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_485),
.Y(n_878)
);

NAND3xp33_ASAP7_75t_L g879 ( 
.A(n_488),
.B(n_503),
.C(n_522),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_620),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_603),
.Y(n_881)
);

BUFx8_ASAP7_75t_SL g882 ( 
.A(n_645),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_606),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_580),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_598),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_598),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_452),
.B(n_621),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_599),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_452),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_599),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_542),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_516),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_542),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_493),
.B(n_627),
.C(n_665),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_413),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_645),
.B(n_655),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_655),
.A2(n_656),
.B1(n_661),
.B2(n_665),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_656),
.A2(n_661),
.B1(n_413),
.B2(n_415),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_415),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_631),
.B(n_357),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_557),
.Y(n_901)
);

INVx4_ASAP7_75t_SL g902 ( 
.A(n_581),
.Y(n_902)
);

AOI22xp33_ASAP7_75t_L g903 ( 
.A1(n_631),
.A2(n_636),
.B1(n_641),
.B2(n_633),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_557),
.Y(n_904)
);

NOR3xp33_ASAP7_75t_L g905 ( 
.A(n_631),
.B(n_636),
.C(n_633),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_544),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_557),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_613),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_652),
.B(n_562),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_544),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_414),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_557),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_631),
.A2(n_636),
.B1(n_641),
.B2(n_633),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_652),
.B(n_562),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_L g915 ( 
.A(n_615),
.B(n_343),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_544),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_613),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_544),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_631),
.B(n_357),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_652),
.B(n_562),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_613),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_557),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_L g923 ( 
.A1(n_631),
.A2(n_636),
.B1(n_641),
.B2(n_633),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_544),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_600),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_464),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_557),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_631),
.B(n_357),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_557),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_613),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_544),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_544),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_544),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_623),
.B(n_631),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_652),
.B(n_562),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_652),
.B(n_562),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_557),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_660),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_652),
.B(n_562),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_623),
.B(n_631),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_544),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_600),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_557),
.Y(n_943)
);

INVx8_ASAP7_75t_L g944 ( 
.A(n_657),
.Y(n_944)
);

AND2x6_ASAP7_75t_L g945 ( 
.A(n_436),
.B(n_495),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_557),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_613),
.Y(n_947)
);

AND3x2_ASAP7_75t_L g948 ( 
.A(n_531),
.B(n_336),
.C(n_328),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_544),
.Y(n_949)
);

XNOR2xp5_ASAP7_75t_L g950 ( 
.A(n_630),
.B(n_631),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_557),
.Y(n_951)
);

BUFx8_ASAP7_75t_SL g952 ( 
.A(n_487),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_557),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_613),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_557),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_623),
.B(n_631),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_635),
.B(n_648),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_544),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_L g959 ( 
.A1(n_631),
.A2(n_636),
.B1(n_641),
.B2(n_633),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_544),
.Y(n_960)
);

NAND2xp33_ASAP7_75t_SL g961 ( 
.A(n_531),
.B(n_343),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_544),
.Y(n_962)
);

INVxp67_ASAP7_75t_SL g963 ( 
.A(n_605),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_544),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_635),
.B(n_648),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_660),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_660),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_631),
.B(n_357),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_544),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_544),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_652),
.B(n_562),
.Y(n_971)
);

BUFx4f_ASAP7_75t_L g972 ( 
.A(n_657),
.Y(n_972)
);

BUFx10_ASAP7_75t_L g973 ( 
.A(n_476),
.Y(n_973)
);

OAI22xp33_ASAP7_75t_SL g974 ( 
.A1(n_509),
.A2(n_336),
.B1(n_639),
.B2(n_628),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_613),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_544),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_414),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_519),
.B(n_526),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_557),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_600),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_464),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_557),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_L g983 ( 
.A1(n_631),
.A2(n_636),
.B1(n_641),
.B2(n_633),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_557),
.Y(n_984)
);

AND2x6_ASAP7_75t_L g985 ( 
.A(n_436),
.B(n_495),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_544),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_557),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_623),
.B(n_631),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_600),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_600),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_544),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_544),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_600),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_652),
.B(n_562),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_557),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_544),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_623),
.B(n_631),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_414),
.Y(n_998)
);

INVx4_ASAP7_75t_L g999 ( 
.A(n_613),
.Y(n_999)
);

BUFx2_ASAP7_75t_L g1000 ( 
.A(n_635),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_631),
.B(n_357),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_557),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_557),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_652),
.B(n_562),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_652),
.B(n_562),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_652),
.B(n_562),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_623),
.B(n_631),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_631),
.A2(n_636),
.B1(n_641),
.B2(n_633),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_600),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_600),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_652),
.B(n_562),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_557),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_635),
.B(n_648),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_628),
.B(n_659),
.C(n_639),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_623),
.B(n_631),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_557),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_623),
.B(n_631),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_544),
.Y(n_1018)
);

AND2x6_ASAP7_75t_L g1019 ( 
.A(n_436),
.B(n_495),
.Y(n_1019)
);

AND2x6_ASAP7_75t_L g1020 ( 
.A(n_436),
.B(n_495),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_900),
.B(n_919),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_744),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_754),
.B(n_692),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_761),
.B(n_978),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_744),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_748),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_748),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_754),
.B(n_765),
.Y(n_1028)
);

INVx3_ASAP7_75t_L g1029 ( 
.A(n_693),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_750),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_903),
.A2(n_923),
.B1(n_959),
.B2(n_913),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_750),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_690),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_761),
.B(n_978),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_752),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_752),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_944),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_763),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_763),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_761),
.B(n_978),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_761),
.B(n_978),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_692),
.B(n_957),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_957),
.B(n_965),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_764),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_928),
.B(n_968),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_965),
.B(n_1013),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_905),
.A2(n_682),
.B1(n_699),
.B2(n_983),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_690),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1001),
.A2(n_1008),
.B1(n_698),
.B2(n_950),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_690),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_977),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_695),
.Y(n_1052)
);

NOR3xp33_ASAP7_75t_L g1053 ( 
.A(n_803),
.B(n_909),
.C(n_688),
.Y(n_1053)
);

AND3x4_ASAP7_75t_L g1054 ( 
.A(n_893),
.B(n_975),
.C(n_954),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_765),
.B(n_1013),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_954),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_695),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_695),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_844),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_764),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_914),
.B(n_920),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_767),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_767),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_771),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_950),
.A2(n_685),
.B1(n_940),
.B2(n_934),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_771),
.Y(n_1066)
);

AND2x4_ASAP7_75t_L g1067 ( 
.A(n_740),
.B(n_735),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_743),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_743),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_693),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_746),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_740),
.B(n_735),
.Y(n_1072)
);

BUFx10_ASAP7_75t_L g1073 ( 
.A(n_729),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_944),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_746),
.Y(n_1075)
);

INVx5_ASAP7_75t_L g1076 ( 
.A(n_693),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_756),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_705),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_756),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_757),
.Y(n_1080)
);

INVx3_ASAP7_75t_R g1081 ( 
.A(n_815),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_757),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_954),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_705),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_833),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_684),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_944),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_684),
.Y(n_1088)
);

NAND2x1_ASAP7_75t_L g1089 ( 
.A(n_736),
.B(n_683),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_735),
.B(n_760),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_975),
.Y(n_1091)
);

INVx4_ASAP7_75t_L g1092 ( 
.A(n_844),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_708),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_816),
.B(n_769),
.Y(n_1094)
);

OAI221xp5_ASAP7_75t_L g1095 ( 
.A1(n_793),
.A2(n_935),
.B1(n_971),
.B2(n_939),
.C(n_936),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_833),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_700),
.B(n_994),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_708),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_735),
.B(n_760),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_693),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_901),
.B(n_904),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_689),
.Y(n_1103)
);

NAND3x1_ASAP7_75t_L g1104 ( 
.A(n_868),
.B(n_824),
.C(n_829),
.Y(n_1104)
);

AND2x4_ASAP7_75t_L g1105 ( 
.A(n_760),
.B(n_925),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_693),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_689),
.Y(n_1107)
);

AO22x2_ASAP7_75t_L g1108 ( 
.A1(n_1014),
.A2(n_988),
.B1(n_997),
.B2(n_956),
.Y(n_1108)
);

INVxp67_ASAP7_75t_L g1109 ( 
.A(n_911),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1006),
.B(n_1011),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1000),
.B(n_703),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_760),
.B(n_925),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_711),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_1000),
.B(n_686),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_711),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_686),
.B(n_687),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_925),
.B(n_942),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_833),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_694),
.Y(n_1119)
);

INVx8_ASAP7_75t_L g1120 ( 
.A(n_844),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_713),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_998),
.B(n_973),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_901),
.B(n_904),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_907),
.B(n_912),
.Y(n_1124)
);

INVxp67_ASAP7_75t_SL g1125 ( 
.A(n_736),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_733),
.B(n_751),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_907),
.B(n_912),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_844),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_713),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_938),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_694),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_710),
.A2(n_1015),
.B1(n_1017),
.B2(n_1007),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_683),
.B(n_917),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_721),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_833),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_975),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_938),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_720),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_720),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_925),
.B(n_942),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_908),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_686),
.B(n_687),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_833),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_722),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_942),
.B(n_980),
.Y(n_1145)
);

AO22x2_ASAP7_75t_L g1146 ( 
.A1(n_1014),
.A2(n_719),
.B1(n_902),
.B2(n_894),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_942),
.B(n_980),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_966),
.Y(n_1148)
);

BUFx4_ASAP7_75t_L g1149 ( 
.A(n_895),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_952),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_722),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_725),
.Y(n_1152)
);

INVx3_ASAP7_75t_R g1153 ( 
.A(n_815),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_725),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_SL g1155 ( 
.A(n_683),
.B(n_917),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_736),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_721),
.Y(n_1157)
);

INVx4_ASAP7_75t_L g1158 ( 
.A(n_844),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_737),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_718),
.A2(n_723),
.B1(n_709),
.B2(n_712),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_683),
.B(n_917),
.Y(n_1161)
);

INVx8_ASAP7_75t_L g1162 ( 
.A(n_944),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_908),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_727),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_739),
.Y(n_1165)
);

AND2x4_ASAP7_75t_L g1166 ( 
.A(n_980),
.B(n_989),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_922),
.B(n_927),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_892),
.A2(n_974),
.B1(n_707),
.B2(n_810),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_727),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_980),
.B(n_989),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_728),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_728),
.Y(n_1172)
);

AND2x6_ASAP7_75t_L g1173 ( 
.A(n_908),
.B(n_930),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_731),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_966),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_944),
.Y(n_1176)
);

INVx4_ASAP7_75t_L g1177 ( 
.A(n_736),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_989),
.B(n_990),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_736),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_989),
.B(n_990),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_731),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_715),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_906),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_906),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_737),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_910),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_910),
.Y(n_1187)
);

NOR2x1p5_ASAP7_75t_L g1188 ( 
.A(n_926),
.B(n_981),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_916),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_693),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_916),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_926),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_918),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_758),
.B(n_973),
.Y(n_1194)
);

INVx5_ASAP7_75t_L g1195 ( 
.A(n_693),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_990),
.B(n_993),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_922),
.B(n_927),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_945),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_812),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_967),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_918),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_945),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_973),
.B(n_780),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_924),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_967),
.Y(n_1205)
);

INVxp33_ASAP7_75t_L g1206 ( 
.A(n_808),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_908),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_953),
.B(n_955),
.Y(n_1208)
);

NAND3x1_ASAP7_75t_L g1209 ( 
.A(n_824),
.B(n_829),
.C(n_832),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_953),
.B(n_955),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_738),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_924),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_981),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_738),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_979),
.B(n_982),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_709),
.A2(n_917),
.B1(n_999),
.B2(n_921),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_979),
.B(n_982),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_786),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_931),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_921),
.A2(n_999),
.B1(n_734),
.B2(n_723),
.Y(n_1220)
);

INVxp67_ASAP7_75t_L g1221 ( 
.A(n_895),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_931),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_990),
.B(n_993),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_993),
.B(n_1009),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_932),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_715),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_932),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_908),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_945),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_973),
.B(n_792),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_715),
.Y(n_1231)
);

INVx8_ASAP7_75t_L g1232 ( 
.A(n_839),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_995),
.B(n_1002),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_972),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_786),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_972),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_691),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_786),
.Y(n_1238)
);

OR2x4_ASAP7_75t_L g1239 ( 
.A(n_834),
.B(n_835),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_933),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_691),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_933),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_687),
.B(n_929),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_941),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_941),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_949),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_795),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_949),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_691),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_921),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_958),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_921),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_795),
.Y(n_1253)
);

OAI221xp5_ASAP7_75t_L g1254 ( 
.A1(n_753),
.A2(n_749),
.B1(n_717),
.B2(n_802),
.C(n_897),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_929),
.B(n_937),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_R g1256 ( 
.A(n_696),
.B(n_732),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_958),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_999),
.B(n_972),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_L g1259 ( 
.A(n_930),
.B(n_947),
.Y(n_1259)
);

BUFx6f_ASAP7_75t_L g1260 ( 
.A(n_691),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_893),
.B(n_785),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_960),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_929),
.B(n_937),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_960),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_795),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_999),
.A2(n_879),
.B1(n_892),
.B2(n_853),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_798),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_945),
.Y(n_1268)
);

NAND2x1p5_ASAP7_75t_L g1269 ( 
.A(n_930),
.B(n_947),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_785),
.B(n_819),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_819),
.B(n_889),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_798),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_993),
.B(n_1009),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_995),
.B(n_1002),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_962),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_962),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_889),
.B(n_948),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_691),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_798),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_759),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_759),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_827),
.B(n_894),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_773),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_930),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_964),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_773),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_799),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_964),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_945),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_930),
.B(n_947),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_899),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_714),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_937),
.B(n_943),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_714),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_714),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_969),
.Y(n_1297)
);

NAND3xp33_ASAP7_75t_L g1298 ( 
.A(n_783),
.B(n_741),
.C(n_879),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1003),
.B(n_1012),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_969),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1003),
.B(n_1012),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1009),
.B(n_1010),
.Y(n_1302)
);

AO22x2_ASAP7_75t_L g1303 ( 
.A1(n_719),
.A2(n_902),
.B1(n_822),
.B2(n_896),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1010),
.B(n_702),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_943),
.B(n_946),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_947),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_899),
.Y(n_1307)
);

OAI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_817),
.A2(n_818),
.B(n_772),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_783),
.A2(n_856),
.B1(n_797),
.B2(n_772),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_891),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_714),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1010),
.B(n_702),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_775),
.Y(n_1313)
);

INVx3_ASAP7_75t_L g1314 ( 
.A(n_945),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_943),
.B(n_946),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_970),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_947),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_784),
.B(n_974),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_799),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_775),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_779),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_946),
.B(n_951),
.Y(n_1322)
);

OAI221xp5_ASAP7_75t_L g1323 ( 
.A1(n_717),
.A2(n_898),
.B1(n_891),
.B2(n_869),
.C(n_845),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_SL g1324 ( 
.A(n_799),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_970),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_840),
.B(n_776),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_799),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_779),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_L g1329 ( 
.A(n_782),
.B(n_826),
.Y(n_1329)
);

INVxp33_ASAP7_75t_L g1330 ( 
.A(n_882),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_976),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_856),
.A2(n_830),
.B1(n_820),
.B2(n_843),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_848),
.Y(n_1333)
);

INVx5_ASAP7_75t_L g1334 ( 
.A(n_945),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_976),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_714),
.Y(n_1336)
);

NOR2xp33_ASAP7_75t_L g1337 ( 
.A(n_778),
.B(n_726),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_951),
.B(n_984),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_951),
.B(n_984),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_778),
.B(n_762),
.Y(n_1340)
);

AO22x2_ASAP7_75t_L g1341 ( 
.A1(n_719),
.A2(n_902),
.B1(n_822),
.B2(n_828),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_781),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_702),
.B(n_704),
.Y(n_1343)
);

INVx8_ASAP7_75t_L g1344 ( 
.A(n_839),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_985),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_986),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_848),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_759),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_984),
.B(n_987),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_SL g1350 ( 
.A1(n_850),
.A2(n_809),
.B1(n_887),
.B2(n_791),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_986),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_991),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_987),
.B(n_1016),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_987),
.B(n_1016),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1016),
.B(n_766),
.Y(n_1355)
);

INVx8_ASAP7_75t_L g1356 ( 
.A(n_839),
.Y(n_1356)
);

AND2x6_ASAP7_75t_L g1357 ( 
.A(n_796),
.B(n_885),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_759),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_991),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_992),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_762),
.B(n_768),
.Y(n_1361)
);

INVx8_ASAP7_75t_L g1362 ( 
.A(n_985),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_787),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_992),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_781),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_996),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_996),
.Y(n_1367)
);

AOI22x1_ASAP7_75t_L g1368 ( 
.A1(n_866),
.A2(n_867),
.B1(n_823),
.B2(n_825),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_759),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_848),
.Y(n_1370)
);

INVx4_ASAP7_75t_L g1371 ( 
.A(n_778),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1018),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_778),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_821),
.B(n_804),
.Y(n_1374)
);

INVx5_ASAP7_75t_L g1375 ( 
.A(n_985),
.Y(n_1375)
);

INVx2_ASAP7_75t_SL g1376 ( 
.A(n_704),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_872),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_704),
.Y(n_1378)
);

AO22x2_ASAP7_75t_L g1379 ( 
.A1(n_719),
.A2(n_902),
.B1(n_828),
.B2(n_796),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_821),
.B(n_697),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_766),
.B(n_881),
.Y(n_1381)
);

AO22x2_ASAP7_75t_L g1382 ( 
.A1(n_828),
.A2(n_796),
.B1(n_777),
.B2(n_848),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1018),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_778),
.Y(n_1384)
);

INVx2_ASAP7_75t_SL g1385 ( 
.A(n_847),
.Y(n_1385)
);

BUFx4f_ASAP7_75t_L g1386 ( 
.A(n_787),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_881),
.B(n_883),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_985),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_762),
.B(n_768),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_851),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_762),
.B(n_768),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_851),
.Y(n_1392)
);

NAND2x1p5_ASAP7_75t_L g1393 ( 
.A(n_768),
.B(n_788),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_851),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_849),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_849),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_847),
.Y(n_1397)
);

INVxp33_ASAP7_75t_SL g1398 ( 
.A(n_872),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_701),
.B(n_716),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_806),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_883),
.B(n_820),
.Y(n_1401)
);

NAND2x1p5_ASAP7_75t_L g1402 ( 
.A(n_788),
.B(n_862),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_806),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_806),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_788),
.B(n_742),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_724),
.B(n_730),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_L g1407 ( 
.A(n_985),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_862),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_745),
.B(n_747),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_811),
.Y(n_1410)
);

INVx1_ASAP7_75t_SL g1411 ( 
.A(n_872),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_873),
.B(n_789),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_787),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_862),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_787),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_985),
.Y(n_1416)
);

NOR2xp33_ASAP7_75t_L g1417 ( 
.A(n_862),
.B(n_755),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_811),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_SL g1419 ( 
.A(n_796),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_770),
.B(n_866),
.Y(n_1420)
);

INVx1_ASAP7_75t_SL g1421 ( 
.A(n_872),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_742),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_811),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_813),
.Y(n_1424)
);

NAND2x1p5_ASAP7_75t_L g1425 ( 
.A(n_885),
.B(n_886),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_SL g1426 ( 
.A(n_961),
.B(n_809),
.Y(n_1426)
);

BUFx6f_ASAP7_75t_SL g1427 ( 
.A(n_873),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_813),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_813),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_876),
.B(n_884),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_876),
.B(n_884),
.Y(n_1431)
);

AND2x6_ASAP7_75t_L g1432 ( 
.A(n_885),
.B(n_831),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_863),
.B(n_864),
.C(n_915),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_814),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_985),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_856),
.A2(n_863),
.B1(n_794),
.B2(n_963),
.Y(n_1436)
);

AND2x6_ASAP7_75t_L g1437 ( 
.A(n_885),
.B(n_831),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_856),
.A2(n_864),
.B1(n_871),
.B2(n_875),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_871),
.B(n_880),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_814),
.Y(n_1440)
);

AND2x4_ASAP7_75t_L g1441 ( 
.A(n_888),
.B(n_890),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_814),
.Y(n_1442)
);

AND2x6_ASAP7_75t_L g1443 ( 
.A(n_888),
.B(n_890),
.Y(n_1443)
);

AND2x6_ASAP7_75t_L g1444 ( 
.A(n_823),
.B(n_825),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_886),
.B(n_842),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_777),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_SL g1447 ( 
.A(n_886),
.B(n_880),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_867),
.B(n_1020),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1019),
.B(n_1020),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_774),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_774),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_790),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_874),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_790),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_800),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_SL g1456 ( 
.A1(n_777),
.A2(n_856),
.B1(n_706),
.B2(n_870),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_877),
.B(n_878),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_800),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_L g1459 ( 
.A(n_877),
.B(n_878),
.C(n_836),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_801),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_836),
.A2(n_886),
.B1(n_837),
.B2(n_854),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_801),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1019),
.B(n_1020),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_841),
.B(n_842),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_854),
.B(n_857),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_805),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_805),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_841),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_857),
.Y(n_1469)
);

BUFx6f_ASAP7_75t_L g1470 ( 
.A(n_1019),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_859),
.A2(n_860),
.B1(n_865),
.B2(n_852),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_859),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_1019),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1019),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1019),
.B(n_1020),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_860),
.A2(n_865),
.B1(n_807),
.B2(n_852),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_874),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_861),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_807),
.B(n_852),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_861),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_807),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_807),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_852),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1019),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_777),
.B(n_838),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1020),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_846),
.B(n_858),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_855),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1020),
.Y(n_1489)
);

INVx4_ASAP7_75t_L g1490 ( 
.A(n_1020),
.Y(n_1490)
);

INVx4_ASAP7_75t_L g1491 ( 
.A(n_874),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_874),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_856),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_856),
.B(n_761),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_690),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_761),
.B(n_978),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_744),
.Y(n_1497)
);

BUFx6f_ASAP7_75t_L g1498 ( 
.A(n_833),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_744),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_900),
.B(n_919),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_754),
.B(n_692),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_954),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_754),
.B(n_765),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_900),
.B(n_919),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_744),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1394),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_L g1507 ( 
.A(n_1491),
.B(n_1250),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1033),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1021),
.A2(n_1500),
.B1(n_1504),
.B2(n_1045),
.Y(n_1509)
);

NOR2x2_ASAP7_75t_L g1510 ( 
.A(n_1452),
.B(n_1460),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_SL g1511 ( 
.A(n_1326),
.B(n_1126),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1031),
.A2(n_1047),
.B1(n_1065),
.B2(n_1049),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1049),
.B(n_1387),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1387),
.B(n_1042),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1042),
.B(n_1043),
.Y(n_1515)
);

NOR2xp67_ASAP7_75t_L g1516 ( 
.A(n_1298),
.B(n_1284),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1173),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1043),
.B(n_1046),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_L g1519 ( 
.A(n_1095),
.B(n_1061),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1053),
.B(n_1110),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1394),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1033),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1309),
.A2(n_1160),
.B1(n_1456),
.B2(n_1436),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1073),
.B(n_1028),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1046),
.B(n_1108),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1108),
.B(n_1412),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1048),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1051),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1068),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1048),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_SL g1531 ( 
.A(n_1073),
.B(n_1503),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1108),
.B(n_1160),
.Y(n_1532)
);

NOR2xp67_ASAP7_75t_L g1533 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1108),
.B(n_1412),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1319),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_SL g1536 ( 
.A(n_1073),
.B(n_1200),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1490),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1399),
.B(n_1406),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1409),
.B(n_1132),
.Y(n_1539)
);

AOI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1308),
.A2(n_1323),
.B1(n_1254),
.B2(n_1266),
.C(n_1309),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1380),
.B(n_1023),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1050),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1050),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1023),
.B(n_1501),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1120),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1436),
.B(n_1116),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1052),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1501),
.B(n_1439),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1052),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1220),
.A2(n_1350),
.B1(n_1102),
.B2(n_1308),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1439),
.B(n_1116),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1068),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1142),
.B(n_1243),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1350),
.A2(n_1168),
.B1(n_1318),
.B2(n_1332),
.Y(n_1554)
);

AOI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1209),
.A2(n_1097),
.B1(n_1419),
.B2(n_1417),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1426),
.A2(n_1427),
.B1(n_1459),
.B2(n_1146),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1054),
.A2(n_1438),
.B1(n_1386),
.B2(n_1457),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1069),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1142),
.B(n_1243),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1069),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1255),
.B(n_1263),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1255),
.B(n_1263),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1294),
.B(n_1315),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1294),
.B(n_1315),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1057),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_SL g1566 ( 
.A(n_1073),
.B(n_1055),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1056),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1057),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1058),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_SL g1570 ( 
.A1(n_1239),
.A2(n_1054),
.B1(n_1398),
.B2(n_1282),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1427),
.A2(n_1146),
.B1(n_1419),
.B2(n_1438),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1058),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1071),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1494),
.B(n_1024),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1071),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1401),
.B(n_1420),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1203),
.B(n_1230),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1209),
.A2(n_1419),
.B1(n_1104),
.B2(n_1216),
.Y(n_1578)
);

NOR2xp33_ASAP7_75t_L g1579 ( 
.A(n_1206),
.B(n_1239),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1401),
.B(n_1374),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1070),
.B(n_1076),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1427),
.A2(n_1146),
.B1(n_1444),
.B2(n_1111),
.Y(n_1582)
);

BUFx6f_ASAP7_75t_L g1583 ( 
.A(n_1070),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1104),
.A2(n_1381),
.B1(n_1329),
.B2(n_1386),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1457),
.A2(n_1386),
.B1(n_1368),
.B2(n_1488),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1075),
.Y(n_1586)
);

BUFx5_ASAP7_75t_L g1587 ( 
.A(n_1357),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1070),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1239),
.B(n_1199),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1114),
.B(n_1444),
.Y(n_1590)
);

NOR2x1p5_ASAP7_75t_L g1591 ( 
.A(n_1182),
.B(n_1226),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1130),
.B(n_1137),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1056),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1114),
.B(n_1444),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1494),
.B(n_1024),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1495),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1146),
.A2(n_1444),
.B1(n_1111),
.B2(n_1493),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1444),
.B(n_1381),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1444),
.B(n_1355),
.Y(n_1599)
);

BUFx6f_ASAP7_75t_L g1600 ( 
.A(n_1070),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1444),
.B(n_1355),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1075),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1094),
.B(n_1194),
.C(n_1277),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1077),
.B(n_1079),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1083),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1130),
.B(n_1137),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1077),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1327),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1493),
.A2(n_1415),
.B1(n_1413),
.B2(n_1494),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1079),
.B(n_1080),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1446),
.B(n_1494),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1080),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1082),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1082),
.B(n_1305),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1446),
.B(n_1141),
.Y(n_1615)
);

INVx5_ASAP7_75t_L g1616 ( 
.A(n_1362),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1322),
.B(n_1338),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1495),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1339),
.B(n_1349),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1353),
.B(n_1354),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1205),
.B(n_1109),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1101),
.B(n_1123),
.Y(n_1622)
);

NOR2xp67_ASAP7_75t_L g1623 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1413),
.A2(n_1415),
.B1(n_1433),
.B2(n_1368),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1083),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1124),
.B(n_1127),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1167),
.B(n_1197),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1413),
.A2(n_1415),
.B1(n_1054),
.B2(n_1155),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1208),
.B(n_1210),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1141),
.B(n_1163),
.Y(n_1630)
);

O2A1O1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1221),
.A2(n_1310),
.B(n_1405),
.C(n_1377),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1390),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1390),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1433),
.A2(n_1382),
.B1(n_1485),
.B2(n_1217),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1091),
.B(n_1136),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1392),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1382),
.A2(n_1485),
.B1(n_1233),
.B2(n_1274),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1292),
.A2(n_1307),
.B(n_1472),
.C(n_1461),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1215),
.B(n_1299),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1448),
.A2(n_1391),
.B(n_1487),
.Y(n_1640)
);

O2A1O1Ixp5_ASAP7_75t_L g1641 ( 
.A1(n_1447),
.A2(n_1471),
.B(n_1291),
.C(n_1476),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1392),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1301),
.B(n_1086),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1205),
.B(n_1256),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1218),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1086),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1070),
.A2(n_1195),
.B(n_1076),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1649)
);

O2A1O1Ixp5_ASAP7_75t_L g1650 ( 
.A1(n_1465),
.A2(n_1089),
.B(n_1383),
.C(n_1340),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1107),
.B(n_1119),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1218),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1107),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1382),
.A2(n_1363),
.B1(n_1025),
.B2(n_1026),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1261),
.A2(n_1259),
.B1(n_1271),
.B2(n_1337),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1235),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1119),
.B(n_1131),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1235),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1131),
.B(n_1138),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1238),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1662)
);

AND2x6_ASAP7_75t_SL g1663 ( 
.A(n_1270),
.B(n_1343),
.Y(n_1663)
);

O2A1O1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1122),
.A2(n_1151),
.B(n_1152),
.C(n_1144),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1238),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1477),
.B(n_1304),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1411),
.A2(n_1421),
.B1(n_1154),
.B2(n_1164),
.C(n_1152),
.Y(n_1667)
);

AND2x4_ASAP7_75t_SL g1668 ( 
.A(n_1250),
.B(n_1252),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1151),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1382),
.A2(n_1363),
.B1(n_1025),
.B2(n_1026),
.Y(n_1670)
);

NAND2x1_ASAP7_75t_L g1671 ( 
.A(n_1357),
.B(n_1432),
.Y(n_1671)
);

O2A1O1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1154),
.A2(n_1169),
.B(n_1171),
.C(n_1164),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1247),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1169),
.B(n_1171),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1173),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1247),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1172),
.B(n_1174),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1678)
);

NOR2xp67_ASAP7_75t_L g1679 ( 
.A(n_1284),
.B(n_1306),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_SL g1680 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1172),
.A2(n_1181),
.B(n_1183),
.C(n_1174),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1181),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1304),
.B(n_1312),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1163),
.B(n_1207),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1183),
.B(n_1184),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1173),
.Y(n_1686)
);

AND2x6_ASAP7_75t_SL g1687 ( 
.A(n_1343),
.B(n_1024),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1184),
.Y(n_1688)
);

AOI22x1_ASAP7_75t_L g1689 ( 
.A1(n_1383),
.A2(n_1063),
.B1(n_1064),
.B2(n_1060),
.Y(n_1689)
);

INVxp67_ASAP7_75t_SL g1690 ( 
.A(n_1395),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1070),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1186),
.B(n_1187),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1186),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1076),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1253),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_SL g1696 ( 
.A(n_1312),
.B(n_1148),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1187),
.B(n_1189),
.Y(n_1697)
);

INVx4_ASAP7_75t_L g1698 ( 
.A(n_1120),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1067),
.A2(n_1072),
.B(n_1441),
.C(n_1191),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1076),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1363),
.A2(n_1303),
.B1(n_1379),
.B2(n_1422),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1379),
.A2(n_1191),
.B1(n_1193),
.B2(n_1189),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1193),
.B(n_1201),
.Y(n_1703)
);

AO22x2_ASAP7_75t_L g1704 ( 
.A1(n_1250),
.A2(n_1252),
.B1(n_1379),
.B2(n_1204),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1201),
.B(n_1204),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1091),
.B(n_1136),
.Y(n_1706)
);

BUFx3_ASAP7_75t_L g1707 ( 
.A(n_1173),
.Y(n_1707)
);

NOR2xp33_ASAP7_75t_L g1708 ( 
.A(n_1502),
.B(n_1175),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1422),
.B(n_1451),
.C(n_1450),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_SL g1710 ( 
.A1(n_1379),
.A2(n_1252),
.B1(n_1250),
.B2(n_1182),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1363),
.A2(n_1303),
.B1(n_1357),
.B2(n_1228),
.Y(n_1711)
);

AND2x6_ASAP7_75t_SL g1712 ( 
.A(n_1343),
.B(n_1024),
.Y(n_1712)
);

AOI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1303),
.A2(n_1222),
.B1(n_1225),
.B2(n_1219),
.C(n_1212),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1212),
.B(n_1219),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1222),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1207),
.B(n_1060),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1022),
.A2(n_1030),
.B1(n_1032),
.B2(n_1027),
.Y(n_1717)
);

INVxp67_ASAP7_75t_L g1718 ( 
.A(n_1502),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_SL g1720 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1227),
.B(n_1240),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1022),
.A2(n_1030),
.B1(n_1032),
.B2(n_1027),
.Y(n_1723)
);

INVx2_ASAP7_75t_SL g1724 ( 
.A(n_1076),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1240),
.B(n_1242),
.Y(n_1725)
);

NAND2x1p5_ASAP7_75t_L g1726 ( 
.A(n_1076),
.B(n_1195),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1063),
.B(n_1064),
.Y(n_1727)
);

BUFx3_ASAP7_75t_L g1728 ( 
.A(n_1173),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1333),
.B(n_1347),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1242),
.B(n_1244),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_L g1731 ( 
.A(n_1306),
.B(n_1317),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1195),
.Y(n_1732)
);

AND2x4_ASAP7_75t_SL g1733 ( 
.A(n_1252),
.B(n_1059),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1244),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1735)
);

AND2x6_ASAP7_75t_SL g1736 ( 
.A(n_1343),
.B(n_1034),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1253),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1067),
.B(n_1072),
.Y(n_1738)
);

NOR2xp67_ASAP7_75t_SL g1739 ( 
.A(n_1195),
.B(n_1334),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1245),
.B(n_1246),
.Y(n_1740)
);

OR2x6_ASAP7_75t_L g1741 ( 
.A(n_1133),
.B(n_1161),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1333),
.B(n_1347),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1265),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_L g1745 ( 
.A(n_1162),
.B(n_1232),
.Y(n_1745)
);

INVx8_ASAP7_75t_L g1746 ( 
.A(n_1120),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1035),
.A2(n_1036),
.B1(n_1039),
.B2(n_1038),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_L g1748 ( 
.A(n_1317),
.B(n_1370),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1303),
.A2(n_1357),
.B1(n_1040),
.B2(n_1041),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1035),
.A2(n_1036),
.B1(n_1039),
.B2(n_1038),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1265),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1264),
.B(n_1275),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1264),
.B(n_1275),
.Y(n_1756)
);

INVx2_ASAP7_75t_SL g1757 ( 
.A(n_1195),
.Y(n_1757)
);

O2A1O1Ixp5_ASAP7_75t_L g1758 ( 
.A1(n_1089),
.A2(n_1469),
.B(n_1286),
.C(n_1289),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1317),
.B(n_1370),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1276),
.A2(n_1289),
.B1(n_1297),
.B2(n_1286),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1276),
.A2(n_1300),
.B(n_1316),
.C(n_1297),
.Y(n_1761)
);

NAND2xp33_ASAP7_75t_L g1762 ( 
.A(n_1162),
.B(n_1232),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1133),
.B(n_1161),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1300),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1267),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1267),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1150),
.Y(n_1767)
);

NAND2xp33_ASAP7_75t_L g1768 ( 
.A(n_1162),
.B(n_1232),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1195),
.A2(n_1375),
.B(n_1334),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1408),
.B(n_1317),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1316),
.Y(n_1771)
);

NAND2xp33_ASAP7_75t_L g1772 ( 
.A(n_1162),
.B(n_1232),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1408),
.B(n_1192),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1044),
.A2(n_1066),
.B1(n_1497),
.B2(n_1062),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1325),
.B(n_1331),
.Y(n_1775)
);

BUFx3_ASAP7_75t_L g1776 ( 
.A(n_1173),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1213),
.B(n_1081),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1325),
.Y(n_1778)
);

NOR2x1_ASAP7_75t_R g1779 ( 
.A(n_1165),
.B(n_1182),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1272),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1331),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1272),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1279),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1335),
.B(n_1346),
.Y(n_1784)
);

INVx4_ASAP7_75t_L g1785 ( 
.A(n_1120),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1081),
.B(n_1153),
.Y(n_1786)
);

NOR2xp67_ASAP7_75t_L g1787 ( 
.A(n_1177),
.B(n_1371),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1395),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1153),
.B(n_1226),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1090),
.B(n_1099),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1090),
.B(n_1099),
.Y(n_1791)
);

INVxp67_ASAP7_75t_L g1792 ( 
.A(n_1311),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1414),
.B(n_1226),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1279),
.Y(n_1794)
);

O2A1O1Ixp33_ASAP7_75t_L g1795 ( 
.A1(n_1335),
.A2(n_1351),
.B(n_1352),
.C(n_1346),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_SL g1796 ( 
.A(n_1090),
.B(n_1099),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1090),
.B(n_1099),
.Y(n_1797)
);

AND2x4_ASAP7_75t_SL g1798 ( 
.A(n_1059),
.B(n_1092),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1078),
.B(n_1084),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1105),
.B(n_1112),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1359),
.B(n_1360),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_1133),
.B(n_1161),
.Y(n_1805)
);

NAND2xp33_ASAP7_75t_SL g1806 ( 
.A(n_1324),
.B(n_1414),
.Y(n_1806)
);

O2A1O1Ixp5_ASAP7_75t_L g1807 ( 
.A1(n_1469),
.A2(n_1372),
.B(n_1364),
.C(n_1367),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1366),
.B(n_1367),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1372),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1490),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1105),
.B(n_1112),
.Y(n_1811)
);

NOR2xp33_ASAP7_75t_L g1812 ( 
.A(n_1231),
.B(n_1234),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1396),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1044),
.A2(n_1505),
.B1(n_1497),
.B2(n_1066),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1396),
.B(n_1062),
.Y(n_1815)
);

NOR3x1_ASAP7_75t_L g1816 ( 
.A(n_1376),
.B(n_1378),
.C(n_1149),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1078),
.B(n_1084),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1105),
.B(n_1112),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1423),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_1288),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1324),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1499),
.Y(n_1822)
);

AO22x1_ASAP7_75t_L g1823 ( 
.A1(n_1357),
.A2(n_1173),
.B1(n_1414),
.B2(n_1443),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1452),
.A2(n_1462),
.B1(n_1460),
.B2(n_1467),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1487),
.B(n_1385),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1385),
.B(n_1397),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1397),
.B(n_1093),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1093),
.B(n_1098),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1098),
.B(n_1113),
.Y(n_1830)
);

NOR2x2_ASAP7_75t_L g1831 ( 
.A(n_1462),
.B(n_1149),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1357),
.A2(n_1041),
.B1(n_1034),
.B2(n_1496),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1336),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1113),
.B(n_1115),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1105),
.B(n_1112),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1115),
.B(n_1121),
.Y(n_1836)
);

AO22x1_ASAP7_75t_L g1837 ( 
.A1(n_1357),
.A2(n_1414),
.B1(n_1443),
.B2(n_1125),
.Y(n_1837)
);

AOI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1034),
.A2(n_1496),
.B1(n_1040),
.B2(n_1041),
.Y(n_1838)
);

NAND2x1_ASAP7_75t_L g1839 ( 
.A(n_1432),
.B(n_1437),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1121),
.B(n_1129),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1129),
.B(n_1134),
.Y(n_1841)
);

NOR2xp33_ASAP7_75t_L g1842 ( 
.A(n_1231),
.B(n_1234),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1134),
.B(n_1157),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1450),
.B(n_1454),
.C(n_1451),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_SL g1845 ( 
.A(n_1117),
.B(n_1140),
.Y(n_1845)
);

O2A1O1Ixp33_ASAP7_75t_L g1846 ( 
.A1(n_1454),
.A2(n_1455),
.B(n_1467),
.C(n_1466),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1157),
.B(n_1159),
.Y(n_1847)
);

OR2x6_ASAP7_75t_L g1848 ( 
.A(n_1258),
.B(n_1393),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_SL g1849 ( 
.A(n_1117),
.B(n_1140),
.Y(n_1849)
);

INVx3_ASAP7_75t_L g1850 ( 
.A(n_1490),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1159),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_SL g1852 ( 
.A(n_1117),
.B(n_1140),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1334),
.A2(n_1375),
.B(n_1362),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1185),
.B(n_1211),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1185),
.B(n_1211),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1214),
.B(n_1455),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1214),
.B(n_1458),
.Y(n_1857)
);

INVxp67_ASAP7_75t_SL g1858 ( 
.A(n_1269),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1423),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1376),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1034),
.B(n_1040),
.Y(n_1861)
);

AOI22xp33_ASAP7_75t_L g1862 ( 
.A1(n_1458),
.A2(n_1466),
.B1(n_1468),
.B2(n_1234),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1269),
.B(n_1258),
.Y(n_1863)
);

OAI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1449),
.A2(n_1475),
.B(n_1463),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1400),
.B(n_1403),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1231),
.B(n_1236),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1400),
.B(n_1403),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1429),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1040),
.B(n_1041),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1361),
.A2(n_1389),
.B(n_1287),
.Y(n_1870)
);

OR2x6_ASAP7_75t_L g1871 ( 
.A(n_1258),
.B(n_1393),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1404),
.B(n_1410),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1269),
.B(n_1361),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1429),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1117),
.B(n_1140),
.Y(n_1875)
);

AND2x4_ASAP7_75t_L g1876 ( 
.A(n_1496),
.B(n_1145),
.Y(n_1876)
);

OAI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1236),
.A2(n_1402),
.B1(n_1037),
.B2(n_1176),
.Y(n_1877)
);

NOR2xp67_ASAP7_75t_L g1878 ( 
.A(n_1177),
.B(n_1371),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1404),
.B(n_1410),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1418),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1418),
.Y(n_1881)
);

NOR2x2_ASAP7_75t_L g1882 ( 
.A(n_1483),
.B(n_1283),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1468),
.A2(n_1236),
.B1(n_1464),
.B2(n_1341),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1464),
.A2(n_1341),
.B1(n_1478),
.B2(n_1480),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1464),
.A2(n_1341),
.B1(n_1478),
.B2(n_1480),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1496),
.A2(n_1341),
.B1(n_1178),
.B2(n_1196),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1424),
.B(n_1428),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1434),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1424),
.B(n_1428),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1440),
.B(n_1430),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_SL g1891 ( 
.A(n_1037),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1371),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1280),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1434),
.B(n_1442),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1440),
.B(n_1430),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1430),
.B(n_1431),
.Y(n_1896)
);

INVx1_ASAP7_75t_SL g1897 ( 
.A(n_1280),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1402),
.B(n_1371),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1145),
.B(n_1147),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1442),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1324),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1402),
.B(n_1384),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1384),
.B(n_1378),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1384),
.B(n_1441),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1393),
.B(n_1389),
.C(n_1361),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1283),
.Y(n_1906)
);

INVx3_ASAP7_75t_L g1907 ( 
.A(n_1334),
.Y(n_1907)
);

BUFx6f_ASAP7_75t_L g1908 ( 
.A(n_1334),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1287),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1384),
.B(n_1441),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1145),
.B(n_1147),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1145),
.B(n_1147),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1313),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1313),
.Y(n_1914)
);

A2O1A1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1441),
.A2(n_1302),
.B(n_1180),
.C(n_1178),
.Y(n_1915)
);

AOI21xp5_ASAP7_75t_L g1916 ( 
.A1(n_1375),
.A2(n_1362),
.B(n_1445),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1430),
.B(n_1431),
.Y(n_1917)
);

INVx4_ASAP7_75t_L g1918 ( 
.A(n_1120),
.Y(n_1918)
);

NOR3xp33_ASAP7_75t_L g1919 ( 
.A(n_1147),
.B(n_1302),
.C(n_1285),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1188),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1320),
.B(n_1321),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1431),
.B(n_1464),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1320),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1431),
.B(n_1321),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1328),
.B(n_1342),
.Y(n_1925)
);

INVx4_ASAP7_75t_L g1926 ( 
.A(n_1375),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1373),
.B(n_1166),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1328),
.B(n_1342),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1365),
.B(n_1166),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1375),
.A2(n_1176),
.B1(n_1037),
.B2(n_1087),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1365),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1481),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1389),
.B(n_1492),
.Y(n_1934)
);

OAI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1484),
.A2(n_1483),
.B(n_1486),
.Y(n_1935)
);

O2A1O1Ixp5_ASAP7_75t_L g1936 ( 
.A1(n_1492),
.A2(n_1445),
.B(n_1481),
.C(n_1482),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1166),
.B(n_1170),
.Y(n_1937)
);

CKINVDCx5p33_ASAP7_75t_R g1938 ( 
.A(n_1188),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1170),
.B(n_1178),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1074),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1482),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1170),
.B(n_1178),
.Y(n_1942)
);

AND2x6_ASAP7_75t_SL g1943 ( 
.A(n_1180),
.B(n_1196),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1373),
.B(n_1180),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1375),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1373),
.B(n_1180),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1196),
.B(n_1223),
.Y(n_1947)
);

OR2x2_ASAP7_75t_L g1948 ( 
.A(n_1373),
.B(n_1453),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1479),
.Y(n_1949)
);

BUFx6f_ASAP7_75t_L g1950 ( 
.A(n_1407),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1407),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1074),
.A2(n_1176),
.B1(n_1087),
.B2(n_1296),
.Y(n_1952)
);

INVx5_ASAP7_75t_L g1953 ( 
.A(n_1362),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1373),
.B(n_1280),
.Y(n_1954)
);

AOI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1196),
.A2(n_1285),
.B1(n_1224),
.B2(n_1223),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1479),
.Y(n_1956)
);

INVx3_ASAP7_75t_L g1957 ( 
.A(n_1362),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1223),
.B(n_1273),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1281),
.B(n_1358),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1445),
.A2(n_1425),
.B(n_1486),
.Y(n_1960)
);

NAND2x1p5_ASAP7_75t_L g1961 ( 
.A(n_1491),
.B(n_1029),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1281),
.B(n_1358),
.Y(n_1962)
);

AOI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1223),
.A2(n_1302),
.B1(n_1273),
.B2(n_1224),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1029),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1074),
.A2(n_1087),
.B1(n_1296),
.B2(n_1260),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1224),
.B(n_1302),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1224),
.B(n_1285),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1479),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1484),
.A2(n_1479),
.B(n_1445),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1273),
.B(n_1285),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1237),
.A2(n_1293),
.B1(n_1348),
.B2(n_1241),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1273),
.B(n_1489),
.Y(n_1972)
);

NAND2xp33_ASAP7_75t_L g1973 ( 
.A(n_1344),
.B(n_1356),
.Y(n_1973)
);

BUFx3_ASAP7_75t_L g1974 ( 
.A(n_1344),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1029),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1432),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1281),
.B(n_1358),
.Y(n_1977)
);

INVx4_ASAP7_75t_L g1978 ( 
.A(n_1059),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1029),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1369),
.B(n_1348),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1453),
.B(n_1443),
.Y(n_1981)
);

INVx2_ASAP7_75t_L g1982 ( 
.A(n_1100),
.Y(n_1982)
);

NOR3xp33_ASAP7_75t_L g1983 ( 
.A(n_1491),
.B(n_1177),
.C(n_1388),
.Y(n_1983)
);

INVx2_ASAP7_75t_L g1984 ( 
.A(n_1100),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1432),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1432),
.Y(n_1986)
);

INVxp33_ASAP7_75t_L g1987 ( 
.A(n_1237),
.Y(n_1987)
);

INVx3_ASAP7_75t_L g1988 ( 
.A(n_1407),
.Y(n_1988)
);

NOR2xp33_ASAP7_75t_L g1989 ( 
.A(n_1369),
.B(n_1348),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_L g1990 ( 
.A1(n_1237),
.A2(n_1293),
.B1(n_1249),
.B2(n_1260),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1443),
.B(n_1491),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1473),
.B(n_1489),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1369),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1443),
.B(n_1432),
.Y(n_1994)
);

INVx2_ASAP7_75t_SL g1995 ( 
.A(n_1100),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1432),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1330),
.B(n_1278),
.Y(n_1997)
);

AND3x1_ASAP7_75t_L g1998 ( 
.A(n_1100),
.B(n_1229),
.C(n_1345),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1443),
.B(n_1437),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1443),
.B(n_1437),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1437),
.B(n_1237),
.Y(n_2001)
);

BUFx3_ASAP7_75t_L g2002 ( 
.A(n_1344),
.Y(n_2002)
);

AOI21xp5_ASAP7_75t_L g2003 ( 
.A1(n_1425),
.A2(n_1268),
.B(n_1229),
.Y(n_2003)
);

INVx2_ASAP7_75t_L g2004 ( 
.A(n_1106),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1237),
.B(n_1278),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1437),
.B(n_1278),
.Y(n_2006)
);

OAI22xp5_ASAP7_75t_SL g2007 ( 
.A1(n_1241),
.A2(n_1295),
.B1(n_1293),
.B2(n_1296),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1437),
.B(n_1278),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1437),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1106),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1241),
.B(n_1278),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1059),
.B(n_1128),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1241),
.B(n_1348),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1241),
.B(n_1260),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1249),
.B(n_1293),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1106),
.Y(n_2016)
);

INVxp67_ASAP7_75t_L g2017 ( 
.A(n_1249),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1249),
.A2(n_1293),
.B1(n_1348),
.B2(n_1260),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1425),
.A2(n_1268),
.B(n_1345),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1249),
.B(n_1296),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1260),
.B(n_1295),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1156),
.B(n_1179),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1473),
.B(n_1489),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1295),
.B(n_1296),
.Y(n_2024)
);

NOR2xp33_ASAP7_75t_L g2025 ( 
.A(n_1295),
.B(n_1179),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1156),
.B(n_1179),
.Y(n_2026)
);

AND2x6_ASAP7_75t_SL g2027 ( 
.A(n_1344),
.B(n_1356),
.Y(n_2027)
);

INVx5_ASAP7_75t_L g2028 ( 
.A(n_1407),
.Y(n_2028)
);

BUFx6f_ASAP7_75t_L g2029 ( 
.A(n_1407),
.Y(n_2029)
);

AND2x4_ASAP7_75t_L g2030 ( 
.A(n_1092),
.B(n_1128),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1156),
.B(n_1179),
.Y(n_2031)
);

NAND2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1106),
.B(n_1268),
.Y(n_2032)
);

INVx8_ASAP7_75t_L g2033 ( 
.A(n_1416),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1295),
.B(n_1473),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1190),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1156),
.B(n_1179),
.Y(n_2036)
);

BUFx3_ASAP7_75t_L g2037 ( 
.A(n_1344),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1156),
.B(n_1416),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1416),
.B(n_1435),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1416),
.B(n_1435),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1190),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1190),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_1092),
.B(n_1158),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_1190),
.A2(n_1268),
.B(n_1345),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1198),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1416),
.B(n_1435),
.Y(n_2046)
);

NAND2x1p5_ASAP7_75t_L g2047 ( 
.A(n_1198),
.B(n_1229),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1356),
.A2(n_1435),
.B1(n_1474),
.B2(n_1470),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1435),
.B(n_1474),
.Y(n_2049)
);

INVxp67_ASAP7_75t_L g2050 ( 
.A(n_1085),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_SL g2051 ( 
.A(n_1356),
.B(n_1085),
.C(n_1498),
.Y(n_2051)
);

NOR2x1p5_ASAP7_75t_L g2052 ( 
.A(n_1092),
.B(n_1158),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1470),
.B(n_1474),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1470),
.B(n_1474),
.Y(n_2054)
);

AOI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1198),
.A2(n_1229),
.B(n_1290),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1198),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_1202),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1470),
.B(n_1474),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1470),
.B(n_1202),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1202),
.B(n_1314),
.Y(n_2060)
);

INVx2_ASAP7_75t_SL g2061 ( 
.A(n_1202),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1356),
.B(n_1085),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1085),
.B(n_1498),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_1085),
.B(n_1096),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1498),
.B(n_1096),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_1290),
.B(n_1388),
.Y(n_2066)
);

INVx2_ASAP7_75t_SL g2067 ( 
.A(n_1290),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1096),
.B(n_1118),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1290),
.B(n_1388),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_1314),
.A2(n_1388),
.B(n_1345),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1314),
.Y(n_2071)
);

OAI22xp5_ASAP7_75t_L g2072 ( 
.A1(n_1128),
.A2(n_1158),
.B1(n_1314),
.B2(n_1135),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1096),
.B(n_1118),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1096),
.B(n_1118),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1118),
.B(n_1498),
.Y(n_2075)
);

AND2x6_ASAP7_75t_SL g2076 ( 
.A(n_1118),
.B(n_1135),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1135),
.A2(n_1143),
.B1(n_1498),
.B2(n_903),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1135),
.B(n_1143),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1135),
.B(n_1143),
.Y(n_2079)
);

BUFx4_ASAP7_75t_L g2080 ( 
.A(n_1143),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1143),
.B(n_1021),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_L g2082 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1021),
.A2(n_919),
.B(n_928),
.C(n_900),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1394),
.Y(n_2084)
);

AOI22xp33_ASAP7_75t_L g2085 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2089)
);

O2A1O1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1021),
.A2(n_919),
.B(n_928),
.C(n_900),
.Y(n_2090)
);

NOR2xp67_ASAP7_75t_L g2091 ( 
.A(n_1298),
.B(n_1284),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1326),
.B(n_343),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_SL g2094 ( 
.A1(n_1031),
.A2(n_630),
.B1(n_336),
.B2(n_900),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1394),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_1047),
.B(n_1065),
.Y(n_2097)
);

INVx5_ASAP7_75t_L g2098 ( 
.A(n_1362),
.Y(n_2098)
);

OAI22xp33_ASAP7_75t_L g2099 ( 
.A1(n_1049),
.A2(n_1045),
.B1(n_1500),
.B2(n_1021),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1326),
.B(n_343),
.Y(n_2103)
);

NOR2xp67_ASAP7_75t_L g2104 ( 
.A(n_1298),
.B(n_1284),
.Y(n_2104)
);

BUFx3_ASAP7_75t_L g2105 ( 
.A(n_1173),
.Y(n_2105)
);

AND2x6_ASAP7_75t_SL g2106 ( 
.A(n_1061),
.B(n_900),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2107)
);

OAI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1049),
.A2(n_903),
.B1(n_923),
.B2(n_913),
.Y(n_2108)
);

AOI22xp33_ASAP7_75t_L g2109 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1394),
.Y(n_2111)
);

AOI22xp33_ASAP7_75t_L g2112 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1326),
.B(n_343),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2115)
);

AOI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2116)
);

NOR2xp33_ASAP7_75t_L g2117 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1326),
.B(n_343),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1394),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2121)
);

INVx8_ASAP7_75t_L g2122 ( 
.A(n_1120),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2125)
);

AND2x2_ASAP7_75t_SL g2126 ( 
.A(n_1021),
.B(n_903),
.Y(n_2126)
);

NOR2xp67_ASAP7_75t_L g2127 ( 
.A(n_1298),
.B(n_1284),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1326),
.B(n_343),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1033),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1394),
.Y(n_2130)
);

AOI22xp5_ASAP7_75t_L g2131 ( 
.A1(n_1021),
.A2(n_919),
.B1(n_928),
.B2(n_900),
.Y(n_2131)
);

NAND2xp5_ASAP7_75t_L g2132 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1394),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2139)
);

OR2x6_ASAP7_75t_L g2140 ( 
.A(n_1133),
.B(n_1161),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1033),
.Y(n_2141)
);

INVx2_ASAP7_75t_SL g2142 ( 
.A(n_1070),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1394),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2144)
);

OR2x6_ASAP7_75t_L g2145 ( 
.A(n_1133),
.B(n_1161),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1031),
.A2(n_915),
.B(n_769),
.Y(n_2146)
);

AOI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1021),
.A2(n_919),
.B1(n_928),
.B2(n_900),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_SL g2150 ( 
.A(n_1326),
.B(n_343),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1033),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2153)
);

INVx2_ASAP7_75t_SL g2154 ( 
.A(n_1070),
.Y(n_2154)
);

NOR2xp33_ASAP7_75t_L g2155 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2155)
);

AOI22xp33_ASAP7_75t_L g2156 ( 
.A1(n_1021),
.A2(n_682),
.B1(n_699),
.B2(n_905),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_1021),
.B(n_1045),
.Y(n_2157)
);

NAND3xp33_ASAP7_75t_L g2158 ( 
.A(n_1021),
.B(n_919),
.C(n_900),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_1605),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1807),
.Y(n_2160)
);

BUFx3_ASAP7_75t_L g2161 ( 
.A(n_1517),
.Y(n_2161)
);

INVx3_ASAP7_75t_L g2162 ( 
.A(n_1926),
.Y(n_2162)
);

AND2x2_ASAP7_75t_SL g2163 ( 
.A(n_1532),
.B(n_2126),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1807),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1936),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2117),
.B(n_2123),
.Y(n_2166)
);

AND2x6_ASAP7_75t_SL g2167 ( 
.A(n_1519),
.B(n_2149),
.Y(n_2167)
);

AND2x4_ASAP7_75t_L g2168 ( 
.A(n_1848),
.B(n_1871),
.Y(n_2168)
);

INVx5_ASAP7_75t_L g2169 ( 
.A(n_2076),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1936),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1529),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1690),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1690),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1529),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1788),
.Y(n_2175)
);

INVx3_ASAP7_75t_L g2176 ( 
.A(n_1926),
.Y(n_2176)
);

INVx2_ASAP7_75t_SL g2177 ( 
.A(n_2080),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1788),
.Y(n_2178)
);

INVx5_ASAP7_75t_L g2179 ( 
.A(n_2076),
.Y(n_2179)
);

INVx5_ASAP7_75t_L g2180 ( 
.A(n_1583),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1672),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1672),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2131),
.B(n_2147),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1681),
.Y(n_2184)
);

BUFx3_ASAP7_75t_L g2185 ( 
.A(n_1517),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2131),
.B(n_2147),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1681),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_1605),
.Y(n_2188)
);

INVxp67_ASAP7_75t_SL g2189 ( 
.A(n_2080),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1761),
.Y(n_2190)
);

BUFx2_ASAP7_75t_L g2191 ( 
.A(n_1704),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1761),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1552),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_R g2194 ( 
.A(n_1820),
.B(n_1767),
.Y(n_2194)
);

BUFx3_ASAP7_75t_L g2195 ( 
.A(n_1517),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1741),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2085),
.B(n_2095),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1795),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_1552),
.Y(n_2199)
);

BUFx6f_ASAP7_75t_L g2200 ( 
.A(n_1741),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1558),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_1795),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_SL g2203 ( 
.A(n_2099),
.B(n_2126),
.Y(n_2203)
);

BUFx6f_ASAP7_75t_L g2204 ( 
.A(n_1741),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_1675),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2149),
.B(n_2155),
.Y(n_2206)
);

BUFx2_ASAP7_75t_L g2207 ( 
.A(n_1704),
.Y(n_2207)
);

INVx4_ASAP7_75t_L g2208 ( 
.A(n_1668),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1558),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1758),
.Y(n_2210)
);

AOI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2155),
.A2(n_2099),
.B1(n_2094),
.B2(n_2126),
.Y(n_2211)
);

OR2x2_ASAP7_75t_L g2212 ( 
.A(n_1526),
.B(n_1534),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_1560),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2085),
.B(n_2095),
.Y(n_2214)
);

BUFx2_ASAP7_75t_L g2215 ( 
.A(n_1704),
.Y(n_2215)
);

INVxp67_ASAP7_75t_L g2216 ( 
.A(n_1708),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2100),
.B(n_2109),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1560),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_L g2219 ( 
.A(n_1509),
.B(n_2094),
.C(n_2158),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2158),
.A2(n_1509),
.B1(n_2108),
.B2(n_2097),
.Y(n_2220)
);

NOR2xp33_ASAP7_75t_L g2221 ( 
.A(n_2082),
.B(n_2086),
.Y(n_2221)
);

HB1xp67_ASAP7_75t_L g2222 ( 
.A(n_1625),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_1583),
.Y(n_2223)
);

OR2x6_ASAP7_75t_L g2224 ( 
.A(n_2140),
.B(n_2145),
.Y(n_2224)
);

BUFx6f_ASAP7_75t_L g2225 ( 
.A(n_1741),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1573),
.Y(n_2226)
);

BUFx12f_ASAP7_75t_L g2227 ( 
.A(n_2027),
.Y(n_2227)
);

INVxp67_ASAP7_75t_L g2228 ( 
.A(n_1625),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1573),
.Y(n_2229)
);

INVx3_ASAP7_75t_L g2230 ( 
.A(n_1583),
.Y(n_2230)
);

BUFx3_ASAP7_75t_L g2231 ( 
.A(n_1675),
.Y(n_2231)
);

BUFx8_ASAP7_75t_SL g2232 ( 
.A(n_1535),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1758),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_1741),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_1848),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_1575),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1760),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_1741),
.Y(n_2238)
);

AND2x4_ASAP7_75t_L g2239 ( 
.A(n_1848),
.B(n_1871),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1760),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_1805),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2100),
.B(n_2109),
.Y(n_2242)
);

NOR2xp33_ASAP7_75t_L g2243 ( 
.A(n_2082),
.B(n_2086),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2112),
.B(n_2116),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1575),
.Y(n_2245)
);

BUFx4f_ASAP7_75t_L g2246 ( 
.A(n_1746),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1848),
.B(n_1871),
.Y(n_2247)
);

BUFx2_ASAP7_75t_L g2248 ( 
.A(n_1704),
.Y(n_2248)
);

AO22x2_ASAP7_75t_L g2249 ( 
.A1(n_1523),
.A2(n_1532),
.B1(n_1557),
.B2(n_2108),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1805),
.Y(n_2250)
);

BUFx8_ASAP7_75t_L g2251 ( 
.A(n_1891),
.Y(n_2251)
);

HB1xp67_ASAP7_75t_L g2252 ( 
.A(n_1567),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_1704),
.Y(n_2253)
);

BUFx3_ASAP7_75t_L g2254 ( 
.A(n_1675),
.Y(n_2254)
);

OR2x2_ASAP7_75t_SL g2255 ( 
.A(n_2087),
.B(n_2088),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1586),
.Y(n_2256)
);

AOI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2097),
.A2(n_1512),
.B1(n_2116),
.B2(n_2112),
.Y(n_2257)
);

OR2x2_ASAP7_75t_L g2258 ( 
.A(n_1526),
.B(n_1534),
.Y(n_2258)
);

INVx3_ASAP7_75t_L g2259 ( 
.A(n_1583),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1586),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1602),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_1567),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1602),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1607),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_1607),
.Y(n_2265)
);

INVx2_ASAP7_75t_SL g2266 ( 
.A(n_1848),
.Y(n_2266)
);

INVxp67_ASAP7_75t_L g2267 ( 
.A(n_1635),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_2087),
.B(n_2088),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1612),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2156),
.B(n_1538),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_1612),
.Y(n_2271)
);

A2O1A1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_2083),
.A2(n_2090),
.B(n_1540),
.C(n_1512),
.Y(n_2272)
);

AND2x4_ASAP7_75t_L g2273 ( 
.A(n_1848),
.B(n_1871),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_1686),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1613),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1613),
.Y(n_2276)
);

BUFx3_ASAP7_75t_L g2277 ( 
.A(n_1686),
.Y(n_2277)
);

INVx2_ASAP7_75t_SL g2278 ( 
.A(n_1871),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2156),
.B(n_1538),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1646),
.Y(n_2280)
);

CKINVDCx20_ASAP7_75t_R g2281 ( 
.A(n_1821),
.Y(n_2281)
);

INVx3_ASAP7_75t_SL g2282 ( 
.A(n_1831),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1646),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_1653),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_1653),
.Y(n_2285)
);

BUFx4f_ASAP7_75t_SL g2286 ( 
.A(n_1535),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1669),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_1686),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2097),
.A2(n_1540),
.B1(n_1550),
.B2(n_2089),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2083),
.B(n_2090),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_1669),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_1805),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_1682),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_1525),
.B(n_1532),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1539),
.B(n_1563),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_1682),
.Y(n_2296)
);

AOI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2089),
.A2(n_2093),
.B1(n_2102),
.B2(n_2101),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1546),
.B(n_1525),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_1546),
.B(n_1597),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_1688),
.Y(n_2300)
);

INVx4_ASAP7_75t_L g2301 ( 
.A(n_1668),
.Y(n_2301)
);

AOI21x1_ASAP7_75t_L g2302 ( 
.A1(n_1539),
.A2(n_1837),
.B(n_1516),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2093),
.B(n_2101),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1688),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_1563),
.B(n_1580),
.Y(n_2305)
);

INVx2_ASAP7_75t_L g2306 ( 
.A(n_1693),
.Y(n_2306)
);

INVx2_ASAP7_75t_SL g2307 ( 
.A(n_1871),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_L g2308 ( 
.A1(n_1550),
.A2(n_2107),
.B1(n_2110),
.B2(n_2102),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_1693),
.Y(n_2309)
);

CKINVDCx20_ASAP7_75t_R g2310 ( 
.A(n_1901),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1520),
.B(n_1555),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1563),
.B(n_1580),
.Y(n_2312)
);

INVx4_ASAP7_75t_L g2313 ( 
.A(n_1668),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_1546),
.B(n_1597),
.Y(n_2314)
);

INVx3_ASAP7_75t_L g2315 ( 
.A(n_1805),
.Y(n_2315)
);

BUFx6f_ASAP7_75t_L g2316 ( 
.A(n_1805),
.Y(n_2316)
);

BUFx3_ASAP7_75t_L g2317 ( 
.A(n_1707),
.Y(n_2317)
);

O2A1O1Ixp33_ASAP7_75t_L g2318 ( 
.A1(n_2107),
.A2(n_2110),
.B(n_2115),
.C(n_2114),
.Y(n_2318)
);

INVx2_ASAP7_75t_L g2319 ( 
.A(n_1715),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2114),
.B(n_2115),
.Y(n_2320)
);

INVx2_ASAP7_75t_SL g2321 ( 
.A(n_1805),
.Y(n_2321)
);

BUFx3_ASAP7_75t_L g2322 ( 
.A(n_1707),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2120),
.A2(n_2124),
.B1(n_2125),
.B2(n_2121),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1715),
.Y(n_2324)
);

INVx3_ASAP7_75t_L g2325 ( 
.A(n_1583),
.Y(n_2325)
);

NOR2x1_ASAP7_75t_L g2326 ( 
.A(n_1709),
.B(n_1844),
.Y(n_2326)
);

INVx4_ASAP7_75t_SL g2327 ( 
.A(n_2007),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_1637),
.B(n_1523),
.Y(n_2328)
);

AOI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_2120),
.A2(n_2124),
.B1(n_2125),
.B2(n_2121),
.Y(n_2329)
);

NAND3xp33_ASAP7_75t_SL g2330 ( 
.A(n_2137),
.B(n_2148),
.C(n_2138),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_SL g2331 ( 
.A(n_1555),
.B(n_1603),
.Y(n_2331)
);

BUFx12f_ASAP7_75t_L g2332 ( 
.A(n_2027),
.Y(n_2332)
);

INVx4_ASAP7_75t_L g2333 ( 
.A(n_1746),
.Y(n_2333)
);

BUFx3_ASAP7_75t_L g2334 ( 
.A(n_1707),
.Y(n_2334)
);

AND2x4_ASAP7_75t_L g2335 ( 
.A(n_1832),
.B(n_1919),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_1576),
.B(n_1513),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1576),
.B(n_1513),
.Y(n_2337)
);

BUFx4f_ASAP7_75t_SL g2338 ( 
.A(n_1535),
.Y(n_2338)
);

INVx2_ASAP7_75t_SL g2339 ( 
.A(n_2140),
.Y(n_2339)
);

BUFx6f_ASAP7_75t_L g2340 ( 
.A(n_2140),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_2140),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2132),
.B(n_2134),
.Y(n_2342)
);

BUFx4f_ASAP7_75t_L g2343 ( 
.A(n_1746),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1734),
.Y(n_2344)
);

BUFx3_ASAP7_75t_L g2345 ( 
.A(n_1728),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1551),
.B(n_2132),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_1551),
.B(n_2134),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_1734),
.Y(n_2348)
);

BUFx8_ASAP7_75t_L g2349 ( 
.A(n_1891),
.Y(n_2349)
);

AOI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_2135),
.A2(n_2137),
.B1(n_2138),
.B2(n_2136),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_1637),
.B(n_1634),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1764),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_1771),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_1593),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_2135),
.B(n_2136),
.Y(n_2355)
);

BUFx2_ASAP7_75t_L g2356 ( 
.A(n_2140),
.Y(n_2356)
);

INVx2_ASAP7_75t_SL g2357 ( 
.A(n_2145),
.Y(n_2357)
);

BUFx3_ASAP7_75t_L g2358 ( 
.A(n_1728),
.Y(n_2358)
);

BUFx3_ASAP7_75t_L g2359 ( 
.A(n_1728),
.Y(n_2359)
);

BUFx3_ASAP7_75t_L g2360 ( 
.A(n_1776),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_1832),
.B(n_1919),
.Y(n_2361)
);

HB1xp67_ASAP7_75t_L g2362 ( 
.A(n_1593),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1771),
.Y(n_2363)
);

BUFx6f_ASAP7_75t_L g2364 ( 
.A(n_2140),
.Y(n_2364)
);

OR2x6_ASAP7_75t_L g2365 ( 
.A(n_2145),
.B(n_1837),
.Y(n_2365)
);

AND2x4_ASAP7_75t_L g2366 ( 
.A(n_1574),
.B(n_1595),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_1778),
.Y(n_2367)
);

AND2x6_ASAP7_75t_L g2368 ( 
.A(n_1776),
.B(n_2105),
.Y(n_2368)
);

BUFx3_ASAP7_75t_L g2369 ( 
.A(n_1776),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1778),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1781),
.Y(n_2371)
);

BUFx6f_ASAP7_75t_L g2372 ( 
.A(n_2145),
.Y(n_2372)
);

BUFx2_ASAP7_75t_L g2373 ( 
.A(n_2145),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1781),
.Y(n_2374)
);

AND2x6_ASAP7_75t_SL g2375 ( 
.A(n_1579),
.B(n_1777),
.Y(n_2375)
);

AND3x2_ASAP7_75t_SL g2376 ( 
.A(n_1571),
.B(n_1578),
.C(n_1554),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1809),
.Y(n_2377)
);

INVx3_ASAP7_75t_L g2378 ( 
.A(n_1583),
.Y(n_2378)
);

INVx3_ASAP7_75t_L g2379 ( 
.A(n_2145),
.Y(n_2379)
);

INVx4_ASAP7_75t_L g2380 ( 
.A(n_1746),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_1809),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_1554),
.B(n_1557),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_1934),
.Y(n_2383)
);

OR2x2_ASAP7_75t_SL g2384 ( 
.A(n_2139),
.B(n_2144),
.Y(n_2384)
);

INVx2_ASAP7_75t_L g2385 ( 
.A(n_1813),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_1701),
.Y(n_2386)
);

NAND2x1p5_ASAP7_75t_L g2387 ( 
.A(n_1671),
.B(n_1739),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2139),
.B(n_2144),
.Y(n_2388)
);

BUFx6f_ASAP7_75t_L g2389 ( 
.A(n_1671),
.Y(n_2389)
);

AOI22xp33_ASAP7_75t_L g2390 ( 
.A1(n_2148),
.A2(n_2153),
.B1(n_2157),
.B2(n_2151),
.Y(n_2390)
);

OR2x6_ASAP7_75t_L g2391 ( 
.A(n_1823),
.B(n_1763),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_1813),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_1844),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1506),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_1506),
.Y(n_2395)
);

AND2x4_ASAP7_75t_SL g2396 ( 
.A(n_2051),
.B(n_1583),
.Y(n_2396)
);

NOR2xp67_ASAP7_75t_L g2397 ( 
.A(n_1905),
.B(n_1541),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2105),
.Y(n_2398)
);

BUFx3_ASAP7_75t_L g2399 ( 
.A(n_2105),
.Y(n_2399)
);

INVx2_ASAP7_75t_L g2400 ( 
.A(n_1941),
.Y(n_2400)
);

BUFx6f_ASAP7_75t_L g2401 ( 
.A(n_1763),
.Y(n_2401)
);

HB1xp67_ASAP7_75t_L g2402 ( 
.A(n_1934),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_1934),
.Y(n_2403)
);

BUFx2_ASAP7_75t_L g2404 ( 
.A(n_1701),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_1521),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_1510),
.Y(n_2406)
);

BUFx3_ASAP7_75t_L g2407 ( 
.A(n_1615),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1521),
.Y(n_2408)
);

AOI22xp5_ASAP7_75t_L g2409 ( 
.A1(n_2151),
.A2(n_2153),
.B1(n_2157),
.B2(n_1577),
.Y(n_2409)
);

HB1xp67_ASAP7_75t_L g2410 ( 
.A(n_1702),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2084),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2084),
.Y(n_2412)
);

AND2x6_ASAP7_75t_L g2413 ( 
.A(n_2012),
.B(n_2030),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_1941),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2096),
.Y(n_2415)
);

INVx1_ASAP7_75t_SL g2416 ( 
.A(n_1882),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_1603),
.B(n_1577),
.Y(n_2417)
);

CKINVDCx20_ASAP7_75t_R g2418 ( 
.A(n_1608),
.Y(n_2418)
);

INVx4_ASAP7_75t_L g2419 ( 
.A(n_1746),
.Y(n_2419)
);

AO22x1_ASAP7_75t_L g2420 ( 
.A1(n_1816),
.A2(n_1858),
.B1(n_1507),
.B2(n_1983),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2096),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2111),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2111),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1541),
.B(n_1553),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2119),
.Y(n_2425)
);

BUFx6f_ASAP7_75t_L g2426 ( 
.A(n_1763),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_1941),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2119),
.Y(n_2428)
);

INVx2_ASAP7_75t_SL g2429 ( 
.A(n_1863),
.Y(n_2429)
);

CKINVDCx8_ASAP7_75t_R g2430 ( 
.A(n_1687),
.Y(n_2430)
);

BUFx12f_ASAP7_75t_L g2431 ( 
.A(n_1608),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_1702),
.Y(n_2432)
);

AND2x4_ASAP7_75t_L g2433 ( 
.A(n_1574),
.B(n_1595),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_1886),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1553),
.B(n_1559),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2130),
.Y(n_2436)
);

INVx5_ASAP7_75t_L g2437 ( 
.A(n_1600),
.Y(n_2437)
);

BUFx6f_ASAP7_75t_L g2438 ( 
.A(n_1600),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1559),
.B(n_1561),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_1561),
.B(n_1562),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_SL g2441 ( 
.A(n_1655),
.B(n_1584),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_1600),
.Y(n_2442)
);

INVx3_ASAP7_75t_L g2443 ( 
.A(n_1600),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_1562),
.B(n_1564),
.Y(n_2444)
);

AOI22xp33_ASAP7_75t_L g2445 ( 
.A1(n_1570),
.A2(n_1511),
.B1(n_1556),
.B2(n_1518),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_1689),
.Y(n_2446)
);

OR2x6_ASAP7_75t_L g2447 ( 
.A(n_1823),
.B(n_1916),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2130),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2106),
.B(n_1514),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2133),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1564),
.B(n_1548),
.Y(n_2451)
);

HB1xp67_ASAP7_75t_L g2452 ( 
.A(n_1615),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1548),
.B(n_1614),
.Y(n_2453)
);

AND2x4_ASAP7_75t_L g2454 ( 
.A(n_1574),
.B(n_1595),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2133),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_1689),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_1863),
.Y(n_2457)
);

INVx2_ASAP7_75t_L g2458 ( 
.A(n_2143),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_1634),
.B(n_1640),
.Y(n_2459)
);

AOI22xp33_ASAP7_75t_L g2460 ( 
.A1(n_1570),
.A2(n_1556),
.B1(n_1518),
.B2(n_1544),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_2143),
.Y(n_2461)
);

INVx3_ASAP7_75t_L g2462 ( 
.A(n_1600),
.Y(n_2462)
);

INVxp67_ASAP7_75t_SL g2463 ( 
.A(n_1709),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_1600),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_1615),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_1691),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1880),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_1655),
.B(n_1584),
.Y(n_2468)
);

CKINVDCx5p33_ASAP7_75t_R g2469 ( 
.A(n_1608),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_1880),
.Y(n_2470)
);

INVx2_ASAP7_75t_SL g2471 ( 
.A(n_1863),
.Y(n_2471)
);

BUFx2_ASAP7_75t_L g2472 ( 
.A(n_1886),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1881),
.Y(n_2473)
);

OAI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_2146),
.A2(n_1650),
.B(n_1641),
.Y(n_2474)
);

INVx2_ASAP7_75t_SL g2475 ( 
.A(n_1507),
.Y(n_2475)
);

AOI22xp33_ASAP7_75t_SL g2476 ( 
.A1(n_2106),
.A2(n_2146),
.B1(n_1585),
.B2(n_2007),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_1881),
.Y(n_2477)
);

OR2x2_ASAP7_75t_L g2478 ( 
.A(n_1640),
.B(n_1598),
.Y(n_2478)
);

NOR2x1p5_ASAP7_75t_L g2479 ( 
.A(n_1974),
.B(n_2002),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_1932),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2092),
.B(n_2103),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_1574),
.B(n_1595),
.Y(n_2482)
);

INVxp67_ASAP7_75t_L g2483 ( 
.A(n_1706),
.Y(n_2483)
);

NAND2x1p5_ASAP7_75t_L g2484 ( 
.A(n_1739),
.B(n_1616),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_1614),
.B(n_2081),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_1822),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1822),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_1711),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_1932),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_1819),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_1846),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1846),
.Y(n_2492)
);

AND3x1_ASAP7_75t_SL g2493 ( 
.A(n_1591),
.B(n_1713),
.C(n_1976),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_1819),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2081),
.B(n_1617),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_1617),
.B(n_1619),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_1619),
.B(n_1620),
.Y(n_2497)
);

AND2x6_ASAP7_75t_L g2498 ( 
.A(n_2012),
.B(n_2030),
.Y(n_2498)
);

AOI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_1589),
.A2(n_1515),
.B1(n_1544),
.B2(n_1516),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_1620),
.B(n_1514),
.Y(n_2500)
);

BUFx6f_ASAP7_75t_L g2501 ( 
.A(n_1691),
.Y(n_2501)
);

INVx3_ASAP7_75t_L g2502 ( 
.A(n_1691),
.Y(n_2502)
);

AND2x4_ASAP7_75t_L g2503 ( 
.A(n_1574),
.B(n_1595),
.Y(n_2503)
);

INVx2_ASAP7_75t_SL g2504 ( 
.A(n_1873),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_SL g2505 ( 
.A(n_2113),
.B(n_2118),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_1604),
.Y(n_2506)
);

AND2x2_ASAP7_75t_L g2507 ( 
.A(n_1582),
.B(n_1611),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_1643),
.B(n_1622),
.Y(n_2508)
);

BUFx2_ASAP7_75t_L g2509 ( 
.A(n_1711),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_1582),
.B(n_1611),
.Y(n_2510)
);

BUFx4f_ASAP7_75t_L g2511 ( 
.A(n_1746),
.Y(n_2511)
);

CKINVDCx5p33_ASAP7_75t_R g2512 ( 
.A(n_1920),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_1819),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_1610),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_1610),
.Y(n_2515)
);

AND2x4_ASAP7_75t_L g2516 ( 
.A(n_1915),
.B(n_1870),
.Y(n_2516)
);

NOR2x1p5_ASAP7_75t_L g2517 ( 
.A(n_1974),
.B(n_2002),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_1648),
.Y(n_2518)
);

AO21x2_ASAP7_75t_L g2519 ( 
.A1(n_1905),
.A2(n_1870),
.B(n_2091),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_1648),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1649),
.Y(n_2521)
);

INVxp67_ASAP7_75t_L g2522 ( 
.A(n_1528),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_1691),
.Y(n_2523)
);

AOI22xp33_ASAP7_75t_L g2524 ( 
.A1(n_1515),
.A2(n_1578),
.B1(n_1571),
.B2(n_2128),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_1649),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1859),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_1643),
.B(n_1622),
.Y(n_2527)
);

INVx4_ASAP7_75t_L g2528 ( 
.A(n_2122),
.Y(n_2528)
);

AND2x2_ASAP7_75t_SL g2529 ( 
.A(n_1745),
.B(n_1762),
.Y(n_2529)
);

BUFx3_ASAP7_75t_L g2530 ( 
.A(n_1974),
.Y(n_2530)
);

AOI22xp33_ASAP7_75t_L g2531 ( 
.A1(n_2150),
.A2(n_2091),
.B1(n_2127),
.B2(n_2104),
.Y(n_2531)
);

BUFx8_ASAP7_75t_SL g2532 ( 
.A(n_1938),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_1626),
.B(n_1627),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_1651),
.Y(n_2534)
);

BUFx3_ASAP7_75t_L g2535 ( 
.A(n_2002),
.Y(n_2535)
);

BUFx6f_ASAP7_75t_L g2536 ( 
.A(n_1691),
.Y(n_2536)
);

NAND2x1p5_ASAP7_75t_L g2537 ( 
.A(n_1616),
.B(n_1953),
.Y(n_2537)
);

CKINVDCx5p33_ASAP7_75t_R g2538 ( 
.A(n_1773),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_1611),
.B(n_1710),
.Y(n_2539)
);

BUFx6f_ASAP7_75t_L g2540 ( 
.A(n_1694),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_2104),
.A2(n_2127),
.B1(n_1598),
.B2(n_1524),
.Y(n_2541)
);

INVx4_ASAP7_75t_L g2542 ( 
.A(n_2122),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_1969),
.Y(n_2543)
);

INVx3_ASAP7_75t_L g2544 ( 
.A(n_1694),
.Y(n_2544)
);

INVxp67_ASAP7_75t_SL g2545 ( 
.A(n_1651),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_1626),
.B(n_1627),
.Y(n_2546)
);

NOR2xp33_ASAP7_75t_L g2547 ( 
.A(n_1528),
.B(n_1599),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_1657),
.Y(n_2548)
);

BUFx6f_ASAP7_75t_L g2549 ( 
.A(n_1694),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_1657),
.Y(n_2550)
);

BUFx6f_ASAP7_75t_L g2551 ( 
.A(n_1694),
.Y(n_2551)
);

OR2x2_ASAP7_75t_L g2552 ( 
.A(n_1654),
.B(n_1670),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_1969),
.Y(n_2553)
);

AOI22xp33_ASAP7_75t_L g2554 ( 
.A1(n_1531),
.A2(n_1566),
.B1(n_1869),
.B2(n_1861),
.Y(n_2554)
);

BUFx4f_ASAP7_75t_L g2555 ( 
.A(n_2122),
.Y(n_2555)
);

CKINVDCx5p33_ASAP7_75t_R g2556 ( 
.A(n_1997),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1659),
.Y(n_2557)
);

INVx5_ASAP7_75t_L g2558 ( 
.A(n_1694),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_1599),
.B(n_1601),
.Y(n_2559)
);

HB1xp67_ASAP7_75t_L g2560 ( 
.A(n_1993),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_1629),
.B(n_1639),
.Y(n_2561)
);

AO21x2_ASAP7_75t_L g2562 ( 
.A1(n_1990),
.A2(n_1983),
.B(n_1935),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_1859),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1659),
.Y(n_2564)
);

HB1xp67_ASAP7_75t_L g2565 ( 
.A(n_1993),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_1661),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_1661),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_1662),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_L g2569 ( 
.A(n_1629),
.B(n_1639),
.Y(n_2569)
);

INVx2_ASAP7_75t_SL g2570 ( 
.A(n_1873),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_1662),
.Y(n_2571)
);

OR2x2_ASAP7_75t_L g2572 ( 
.A(n_1654),
.B(n_1670),
.Y(n_2572)
);

BUFx4f_ASAP7_75t_L g2573 ( 
.A(n_2122),
.Y(n_2573)
);

BUFx2_ASAP7_75t_L g2574 ( 
.A(n_1751),
.Y(n_2574)
);

INVx2_ASAP7_75t_L g2575 ( 
.A(n_1859),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_1826),
.B(n_1716),
.Y(n_2576)
);

OR2x6_ASAP7_75t_L g2577 ( 
.A(n_1916),
.B(n_1853),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_1674),
.Y(n_2578)
);

INVx3_ASAP7_75t_L g2579 ( 
.A(n_1694),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_1674),
.Y(n_2580)
);

CKINVDCx5p33_ASAP7_75t_R g2581 ( 
.A(n_1891),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_1677),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_1677),
.Y(n_2583)
);

BUFx3_ASAP7_75t_L g2584 ( 
.A(n_2037),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_1685),
.Y(n_2585)
);

INVxp67_ASAP7_75t_SL g2586 ( 
.A(n_1685),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_1692),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_1692),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_1826),
.B(n_1716),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_1697),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_1697),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_SL g2592 ( 
.A(n_1699),
.B(n_1638),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_SL g2593 ( 
.A(n_1638),
.B(n_1585),
.Y(n_2593)
);

AND2x6_ASAP7_75t_L g2594 ( 
.A(n_2012),
.B(n_2030),
.Y(n_2594)
);

INVx4_ASAP7_75t_L g2595 ( 
.A(n_2122),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_1703),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_1703),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_1716),
.B(n_1705),
.Y(n_2598)
);

BUFx3_ASAP7_75t_L g2599 ( 
.A(n_2037),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_1868),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_1705),
.B(n_1714),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_1710),
.B(n_1751),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_1630),
.B(n_1684),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_1630),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_1868),
.Y(n_2605)
);

OR2x6_ASAP7_75t_L g2606 ( 
.A(n_1853),
.B(n_1960),
.Y(n_2606)
);

BUFx2_ASAP7_75t_L g2607 ( 
.A(n_1713),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_1714),
.B(n_1721),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_SL g2609 ( 
.A1(n_1718),
.A2(n_1601),
.B1(n_1594),
.B2(n_1590),
.Y(n_2609)
);

INVx1_ASAP7_75t_L g2610 ( 
.A(n_1721),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_1868),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_1722),
.Y(n_2612)
);

INVx2_ASAP7_75t_L g2613 ( 
.A(n_1874),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_1722),
.Y(n_2614)
);

INVxp67_ASAP7_75t_SL g2615 ( 
.A(n_1725),
.Y(n_2615)
);

OR2x2_ASAP7_75t_L g2616 ( 
.A(n_1590),
.B(n_1594),
.Y(n_2616)
);

OR2x2_ASAP7_75t_SL g2617 ( 
.A(n_1873),
.B(n_1991),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_1725),
.B(n_1730),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_1874),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_1730),
.B(n_1735),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_1874),
.Y(n_2621)
);

OR2x2_ASAP7_75t_L g2622 ( 
.A(n_1628),
.B(n_1624),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_1735),
.B(n_1740),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_1740),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_1742),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_1742),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_1888),
.Y(n_2627)
);

INVx4_ASAP7_75t_L g2628 ( 
.A(n_2122),
.Y(n_2628)
);

AOI22xp33_ASAP7_75t_L g2629 ( 
.A1(n_1861),
.A2(n_1869),
.B1(n_1876),
.B2(n_1947),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_1888),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_1749),
.B(n_1750),
.Y(n_2631)
);

INVx2_ASAP7_75t_SL g2632 ( 
.A(n_2028),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_1749),
.B(n_1750),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_L g2634 ( 
.A(n_1752),
.B(n_1755),
.Y(n_2634)
);

INVx2_ASAP7_75t_SL g2635 ( 
.A(n_2028),
.Y(n_2635)
);

INVx2_ASAP7_75t_L g2636 ( 
.A(n_1888),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_1899),
.B(n_1963),
.Y(n_2637)
);

HB1xp67_ASAP7_75t_L g2638 ( 
.A(n_1718),
.Y(n_2638)
);

HB1xp67_ASAP7_75t_L g2639 ( 
.A(n_1890),
.Y(n_2639)
);

BUFx3_ASAP7_75t_L g2640 ( 
.A(n_2037),
.Y(n_2640)
);

INVx3_ASAP7_75t_L g2641 ( 
.A(n_1732),
.Y(n_2641)
);

BUFx5_ASAP7_75t_L g2642 ( 
.A(n_1976),
.Y(n_2642)
);

BUFx6f_ASAP7_75t_L g2643 ( 
.A(n_1732),
.Y(n_2643)
);

INVx5_ASAP7_75t_L g2644 ( 
.A(n_1732),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_1752),
.B(n_1755),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_1891),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_SL g2647 ( 
.A(n_1624),
.B(n_1628),
.Y(n_2647)
);

NOR2x1_ASAP7_75t_L g2648 ( 
.A(n_2052),
.B(n_1973),
.Y(n_2648)
);

AOI22xp5_ASAP7_75t_L g2649 ( 
.A1(n_1866),
.A2(n_1838),
.B1(n_1842),
.B2(n_1812),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_1508),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_1756),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_1756),
.Y(n_2652)
);

BUFx2_ASAP7_75t_L g2653 ( 
.A(n_1943),
.Y(n_2653)
);

NOR2xp33_ASAP7_75t_L g2654 ( 
.A(n_1630),
.B(n_1684),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_1861),
.A2(n_1869),
.B1(n_1876),
.B2(n_1947),
.Y(n_2655)
);

INVx5_ASAP7_75t_L g2656 ( 
.A(n_1732),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_1732),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_1899),
.B(n_1963),
.Y(n_2658)
);

NOR2xp33_ASAP7_75t_L g2659 ( 
.A(n_1684),
.B(n_1866),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_1943),
.Y(n_2660)
);

NAND2xp5_ASAP7_75t_L g2661 ( 
.A(n_1775),
.B(n_1784),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_1800),
.B(n_1802),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_1508),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_1800),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_1802),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_1803),
.B(n_1804),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1803),
.Y(n_2667)
);

INVx4_ASAP7_75t_L g2668 ( 
.A(n_1978),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_1732),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_1786),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_1804),
.Y(n_2671)
);

INVxp33_ASAP7_75t_SL g2672 ( 
.A(n_1779),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_1894),
.B(n_1884),
.Y(n_2673)
);

INVx4_ASAP7_75t_L g2674 ( 
.A(n_1978),
.Y(n_2674)
);

BUFx3_ASAP7_75t_L g2675 ( 
.A(n_1892),
.Y(n_2675)
);

NOR2xp33_ASAP7_75t_L g2676 ( 
.A(n_1896),
.B(n_1917),
.Y(n_2676)
);

AND2x4_ASAP7_75t_L g2677 ( 
.A(n_1899),
.B(n_1876),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_1808),
.B(n_1815),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_1732),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_1894),
.B(n_1884),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_1808),
.B(n_1815),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_1865),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_1865),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_1885),
.B(n_1609),
.Y(n_2684)
);

AOI221xp5_ASAP7_75t_L g2685 ( 
.A1(n_1631),
.A2(n_1644),
.B1(n_1621),
.B2(n_1664),
.C(n_1606),
.Y(n_2685)
);

HB1xp67_ASAP7_75t_L g2686 ( 
.A(n_1890),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_1867),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_1861),
.A2(n_1869),
.B1(n_1876),
.B2(n_1947),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_1867),
.Y(n_2689)
);

AOI22xp5_ASAP7_75t_L g2690 ( 
.A1(n_1838),
.A2(n_1910),
.B1(n_1904),
.B2(n_1609),
.Y(n_2690)
);

INVx2_ASAP7_75t_SL g2691 ( 
.A(n_2028),
.Y(n_2691)
);

AND2x4_ASAP7_75t_L g2692 ( 
.A(n_1899),
.B(n_1876),
.Y(n_2692)
);

NAND2x1p5_ASAP7_75t_L g2693 ( 
.A(n_1616),
.B(n_1953),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_1872),
.Y(n_2694)
);

BUFx12f_ASAP7_75t_L g2695 ( 
.A(n_1687),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_1895),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_1824),
.B(n_1895),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_1948),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_1508),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_1872),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_1879),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_1856),
.B(n_1857),
.Y(n_2702)
);

AND2x4_ASAP7_75t_L g2703 ( 
.A(n_1899),
.B(n_1864),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_1861),
.A2(n_1869),
.B1(n_1591),
.B2(n_1696),
.Y(n_2704)
);

INVx5_ASAP7_75t_L g2705 ( 
.A(n_1908),
.Y(n_2705)
);

INVx2_ASAP7_75t_L g2706 ( 
.A(n_1522),
.Y(n_2706)
);

INVx2_ASAP7_75t_SL g2707 ( 
.A(n_2028),
.Y(n_2707)
);

BUFx6f_ASAP7_75t_L g2708 ( 
.A(n_1908),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_1522),
.Y(n_2709)
);

INVx5_ASAP7_75t_L g2710 ( 
.A(n_1908),
.Y(n_2710)
);

BUFx6f_ASAP7_75t_L g2711 ( 
.A(n_1908),
.Y(n_2711)
);

CKINVDCx5p33_ASAP7_75t_R g2712 ( 
.A(n_1789),
.Y(n_2712)
);

INVx3_ASAP7_75t_L g2713 ( 
.A(n_1908),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_1857),
.B(n_1896),
.Y(n_2714)
);

NAND3xp33_ASAP7_75t_L g2715 ( 
.A(n_1631),
.B(n_1862),
.C(n_1664),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_1892),
.Y(n_2716)
);

CKINVDCx16_ASAP7_75t_R g2717 ( 
.A(n_1972),
.Y(n_2717)
);

AO22x1_ASAP7_75t_L g2718 ( 
.A1(n_1816),
.A2(n_1858),
.B1(n_1965),
.B2(n_1770),
.Y(n_2718)
);

INVx2_ASAP7_75t_SL g2719 ( 
.A(n_2028),
.Y(n_2719)
);

INVx1_ASAP7_75t_SL g2720 ( 
.A(n_1893),
.Y(n_2720)
);

BUFx8_ASAP7_75t_L g2721 ( 
.A(n_1587),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_1877),
.B(n_1748),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_1522),
.Y(n_2723)
);

BUFx6f_ASAP7_75t_L g2724 ( 
.A(n_1908),
.Y(n_2724)
);

INVx5_ASAP7_75t_L g2725 ( 
.A(n_1616),
.Y(n_2725)
);

BUFx6f_ASAP7_75t_L g2726 ( 
.A(n_1839),
.Y(n_2726)
);

INVx2_ASAP7_75t_SL g2727 ( 
.A(n_2028),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_1879),
.Y(n_2728)
);

BUFx6f_ASAP7_75t_L g2729 ( 
.A(n_1839),
.Y(n_2729)
);

AND3x1_ASAP7_75t_L g2730 ( 
.A(n_2051),
.B(n_1793),
.C(n_1959),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_1885),
.B(n_1883),
.Y(n_2731)
);

INVxp67_ASAP7_75t_L g2732 ( 
.A(n_1729),
.Y(n_2732)
);

INVxp67_ASAP7_75t_SL g2733 ( 
.A(n_1990),
.Y(n_2733)
);

HB1xp67_ASAP7_75t_L g2734 ( 
.A(n_1948),
.Y(n_2734)
);

BUFx2_ASAP7_75t_L g2735 ( 
.A(n_1663),
.Y(n_2735)
);

OAI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_1650),
.A2(n_1641),
.B(n_2044),
.Y(n_2736)
);

BUFx3_ASAP7_75t_L g2737 ( 
.A(n_1940),
.Y(n_2737)
);

BUFx3_ASAP7_75t_L g2738 ( 
.A(n_1940),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_1527),
.Y(n_2739)
);

NOR2xp67_ASAP7_75t_L g2740 ( 
.A(n_2028),
.B(n_1949),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_1887),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_1887),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_1527),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_1917),
.B(n_1825),
.Y(n_2744)
);

AOI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_1666),
.A2(n_1729),
.B1(n_1743),
.B2(n_1536),
.Y(n_2745)
);

AND2x4_ASAP7_75t_L g2746 ( 
.A(n_1864),
.B(n_1972),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_1889),
.Y(n_2747)
);

BUFx6f_ASAP7_75t_L g2748 ( 
.A(n_1961),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_1825),
.B(n_1922),
.Y(n_2749)
);

BUFx6f_ASAP7_75t_L g2750 ( 
.A(n_1961),
.Y(n_2750)
);

BUFx2_ASAP7_75t_L g2751 ( 
.A(n_1663),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_1922),
.B(n_1727),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_1894),
.B(n_1527),
.Y(n_2753)
);

BUFx2_ASAP7_75t_L g2754 ( 
.A(n_1587),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_1948),
.Y(n_2755)
);

BUFx4f_ASAP7_75t_L g2756 ( 
.A(n_2012),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_1889),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_1530),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_L g2759 ( 
.A1(n_1743),
.A2(n_1680),
.B1(n_1683),
.B2(n_1678),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_1587),
.Y(n_2760)
);

BUFx2_ASAP7_75t_L g2761 ( 
.A(n_1587),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1727),
.B(n_1799),
.Y(n_2762)
);

OR2x6_ASAP7_75t_L g2763 ( 
.A(n_1960),
.B(n_1647),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_1727),
.B(n_1799),
.Y(n_2764)
);

AND2x4_ASAP7_75t_L g2765 ( 
.A(n_1972),
.B(n_1533),
.Y(n_2765)
);

CKINVDCx20_ASAP7_75t_R g2766 ( 
.A(n_1806),
.Y(n_2766)
);

BUFx6f_ASAP7_75t_L g2767 ( 
.A(n_1961),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_1971),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_1530),
.Y(n_2769)
);

CKINVDCx8_ASAP7_75t_R g2770 ( 
.A(n_1712),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_1862),
.A2(n_1956),
.B1(n_1968),
.B2(n_1949),
.Y(n_2771)
);

AND2x4_ASAP7_75t_L g2772 ( 
.A(n_1533),
.B(n_1623),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_1956),
.A2(n_1968),
.B1(n_1939),
.B2(n_1942),
.Y(n_2773)
);

HB1xp67_ASAP7_75t_L g2774 ( 
.A(n_1971),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_1530),
.Y(n_2775)
);

OR2x6_ASAP7_75t_L g2776 ( 
.A(n_1647),
.B(n_1769),
.Y(n_2776)
);

INVx2_ASAP7_75t_L g2777 ( 
.A(n_1542),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_1542),
.Y(n_2778)
);

AND2x4_ASAP7_75t_L g2779 ( 
.A(n_1623),
.B(n_1679),
.Y(n_2779)
);

INVx2_ASAP7_75t_L g2780 ( 
.A(n_1542),
.Y(n_2780)
);

AND2x4_ASAP7_75t_L g2781 ( 
.A(n_1679),
.B(n_1731),
.Y(n_2781)
);

NOR2xp67_ASAP7_75t_L g2782 ( 
.A(n_2028),
.B(n_1988),
.Y(n_2782)
);

CKINVDCx20_ASAP7_75t_R g2783 ( 
.A(n_1940),
.Y(n_2783)
);

AND2x4_ASAP7_75t_L g2784 ( 
.A(n_1731),
.B(n_2012),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_1799),
.B(n_1817),
.Y(n_2785)
);

INVx2_ASAP7_75t_L g2786 ( 
.A(n_1543),
.Y(n_2786)
);

HB1xp67_ASAP7_75t_L g2787 ( 
.A(n_2018),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_1543),
.Y(n_2788)
);

AND2x4_ASAP7_75t_L g2789 ( 
.A(n_2030),
.B(n_2043),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_L g2790 ( 
.A(n_1817),
.B(n_1717),
.Y(n_2790)
);

OR2x2_ASAP7_75t_L g2791 ( 
.A(n_1883),
.B(n_1991),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_1817),
.B(n_1717),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_SL g2793 ( 
.A(n_1877),
.B(n_1759),
.Y(n_2793)
);

AOI21x1_ASAP7_75t_L g2794 ( 
.A1(n_2044),
.A2(n_2070),
.B(n_2055),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_R g2795 ( 
.A(n_1768),
.B(n_1772),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_1543),
.Y(n_2796)
);

BUFx12f_ASAP7_75t_SL g2797 ( 
.A(n_1545),
.Y(n_2797)
);

AND2x4_ASAP7_75t_L g2798 ( 
.A(n_2030),
.B(n_2043),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_1793),
.A2(n_1720),
.B1(n_1738),
.B2(n_1719),
.Y(n_2799)
);

INVx5_ASAP7_75t_L g2800 ( 
.A(n_1616),
.Y(n_2800)
);

INVx2_ASAP7_75t_SL g2801 ( 
.A(n_1961),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_1937),
.B(n_1939),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_L g2803 ( 
.A(n_1723),
.B(n_1747),
.Y(n_2803)
);

BUFx2_ASAP7_75t_L g2804 ( 
.A(n_1587),
.Y(n_2804)
);

BUFx3_ASAP7_75t_L g2805 ( 
.A(n_1992),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_1770),
.B(n_2077),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_1547),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_1723),
.B(n_1747),
.Y(n_2808)
);

INVx1_ASAP7_75t_SL g2809 ( 
.A(n_1893),
.Y(n_2809)
);

AND2x6_ASAP7_75t_L g2810 ( 
.A(n_2043),
.B(n_1537),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_1547),
.Y(n_2811)
);

AND2x4_ASAP7_75t_L g2812 ( 
.A(n_2043),
.B(n_1988),
.Y(n_2812)
);

AND2x4_ASAP7_75t_L g2813 ( 
.A(n_2043),
.B(n_1988),
.Y(n_2813)
);

O2A1O1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2272),
.A2(n_1592),
.B(n_2077),
.C(n_1860),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2211),
.A2(n_1774),
.B1(n_1814),
.B2(n_1753),
.Y(n_2815)
);

NOR2x1_ASAP7_75t_L g2816 ( 
.A(n_2330),
.B(n_2018),
.Y(n_2816)
);

INVx1_ASAP7_75t_SL g2817 ( 
.A(n_2720),
.Y(n_2817)
);

AOI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2166),
.A2(n_1902),
.B1(n_1898),
.B2(n_1790),
.Y(n_2818)
);

OR2x6_ASAP7_75t_SL g2819 ( 
.A(n_2219),
.B(n_2581),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_2409),
.B(n_1937),
.Y(n_2820)
);

OAI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_2211),
.A2(n_1774),
.B1(n_1814),
.B2(n_1753),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2577),
.A2(n_1733),
.B(n_2003),
.Y(n_2822)
);

AOI21xp5_ASAP7_75t_L g2823 ( 
.A1(n_2577),
.A2(n_1733),
.B(n_2003),
.Y(n_2823)
);

AO32x1_ASAP7_75t_L g2824 ( 
.A1(n_2160),
.A2(n_1930),
.A3(n_1965),
.B1(n_1667),
.B2(n_2067),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_SL g2825 ( 
.A(n_2409),
.B(n_1942),
.Y(n_2825)
);

OR2x6_ASAP7_75t_L g2826 ( 
.A(n_2577),
.B(n_1930),
.Y(n_2826)
);

BUFx2_ASAP7_75t_L g2827 ( 
.A(n_2401),
.Y(n_2827)
);

NOR2xp67_ASAP7_75t_SL g2828 ( 
.A(n_2169),
.B(n_2179),
.Y(n_2828)
);

BUFx6f_ASAP7_75t_L g2829 ( 
.A(n_2530),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2308),
.B(n_1958),
.Y(n_2830)
);

INVx2_ASAP7_75t_SL g2831 ( 
.A(n_2737),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2577),
.A2(n_1733),
.B(n_2019),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2166),
.B(n_1958),
.Y(n_2833)
);

INVx5_ASAP7_75t_L g2834 ( 
.A(n_2169),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2308),
.B(n_1966),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2171),
.Y(n_2836)
);

AOI21xp5_ASAP7_75t_L g2837 ( 
.A1(n_2606),
.A2(n_2019),
.B(n_2072),
.Y(n_2837)
);

AOI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2257),
.A2(n_1791),
.B1(n_1797),
.B2(n_1796),
.Y(n_2838)
);

NAND3xp33_ASAP7_75t_L g2839 ( 
.A(n_2219),
.B(n_1667),
.C(n_1955),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2298),
.B(n_2539),
.Y(n_2840)
);

OAI21xp5_ASAP7_75t_L g2841 ( 
.A1(n_2272),
.A2(n_2070),
.B(n_2055),
.Y(n_2841)
);

AOI221xp5_ASAP7_75t_L g2842 ( 
.A1(n_2203),
.A2(n_1792),
.B1(n_1833),
.B2(n_1860),
.C(n_1929),
.Y(n_2842)
);

AOI21xp5_ASAP7_75t_L g2843 ( 
.A1(n_2606),
.A2(n_2072),
.B(n_1999),
.Y(n_2843)
);

INVx2_ASAP7_75t_L g2844 ( 
.A(n_2480),
.Y(n_2844)
);

O2A1O1Ixp5_ASAP7_75t_L g2845 ( 
.A1(n_2331),
.A2(n_2049),
.B(n_1994),
.C(n_2000),
.Y(n_2845)
);

NOR2xp33_ASAP7_75t_L g2846 ( 
.A(n_2206),
.B(n_1966),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2297),
.B(n_1970),
.Y(n_2847)
);

AO32x1_ASAP7_75t_L g2848 ( 
.A1(n_2160),
.A2(n_2061),
.A3(n_1964),
.B1(n_1975),
.B2(n_2067),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2480),
.Y(n_2849)
);

INVx4_ASAP7_75t_L g2850 ( 
.A(n_2169),
.Y(n_2850)
);

NOR3xp33_ASAP7_75t_L g2851 ( 
.A(n_2417),
.B(n_1811),
.C(n_1801),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2480),
.Y(n_2852)
);

BUFx8_ASAP7_75t_L g2853 ( 
.A(n_2431),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2297),
.B(n_1970),
.Y(n_2854)
);

AO32x1_ASAP7_75t_L g2855 ( 
.A1(n_2160),
.A2(n_2061),
.A3(n_2067),
.B1(n_1995),
.B2(n_1975),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2171),
.Y(n_2856)
);

NOR2xp33_ASAP7_75t_L g2857 ( 
.A(n_2206),
.B(n_1779),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2294),
.B(n_1924),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2323),
.B(n_2329),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2323),
.B(n_2329),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2390),
.B(n_1792),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2171),
.Y(n_2862)
);

INVx5_ASAP7_75t_L g2863 ( 
.A(n_2169),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2390),
.B(n_2221),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2489),
.Y(n_2865)
);

AND2x2_ASAP7_75t_L g2866 ( 
.A(n_2298),
.B(n_1921),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_L g2867 ( 
.A(n_2221),
.B(n_1833),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_L g2868 ( 
.A(n_2243),
.B(n_1929),
.Y(n_2868)
);

AOI21xp5_ASAP7_75t_L g2869 ( 
.A1(n_2606),
.A2(n_1726),
.B(n_1581),
.Y(n_2869)
);

OA22x2_ASAP7_75t_L g2870 ( 
.A1(n_2289),
.A2(n_1952),
.B1(n_1985),
.B2(n_1986),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2318),
.B(n_1981),
.Y(n_2871)
);

NOR2xp33_ASAP7_75t_L g2872 ( 
.A(n_2167),
.B(n_1818),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2171),
.Y(n_2873)
);

NOR2xp33_ASAP7_75t_L g2874 ( 
.A(n_2167),
.B(n_1835),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2606),
.A2(n_1726),
.B(n_1581),
.Y(n_2875)
);

AOI21xp5_ASAP7_75t_L g2876 ( 
.A1(n_2606),
.A2(n_1726),
.B(n_1581),
.Y(n_2876)
);

O2A1O1Ixp33_ASAP7_75t_L g2877 ( 
.A1(n_2417),
.A2(n_1933),
.B(n_1967),
.C(n_1911),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2474),
.A2(n_1581),
.B(n_1588),
.Y(n_2878)
);

O2A1O1Ixp5_ASAP7_75t_L g2879 ( 
.A1(n_2331),
.A2(n_1981),
.B(n_2026),
.C(n_2031),
.Y(n_2879)
);

A2O1A1Ixp33_ASAP7_75t_L g2880 ( 
.A1(n_2257),
.A2(n_1959),
.B(n_1962),
.C(n_1977),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2174),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2289),
.A2(n_2350),
.B1(n_2382),
.B2(n_2607),
.Y(n_2882)
);

A2O1A1Ixp33_ASAP7_75t_L g2883 ( 
.A1(n_2318),
.A2(n_1962),
.B(n_1977),
.C(n_1903),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2243),
.B(n_1924),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_SL g2885 ( 
.A(n_2350),
.B(n_1955),
.Y(n_2885)
);

INVxp67_ASAP7_75t_L g2886 ( 
.A(n_2522),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2174),
.Y(n_2887)
);

OAI22xp5_ASAP7_75t_L g2888 ( 
.A1(n_2382),
.A2(n_1897),
.B1(n_2048),
.B2(n_1827),
.Y(n_2888)
);

NAND2xp5_ASAP7_75t_L g2889 ( 
.A(n_2268),
.B(n_1927),
.Y(n_2889)
);

HB1xp67_ASAP7_75t_L g2890 ( 
.A(n_2252),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2268),
.B(n_1944),
.Y(n_2891)
);

AOI33xp33_ASAP7_75t_L g2892 ( 
.A1(n_2406),
.A2(n_1897),
.A3(n_1851),
.B1(n_1931),
.B2(n_1909),
.B3(n_1913),
.Y(n_2892)
);

OAI21xp33_ASAP7_75t_L g2893 ( 
.A1(n_2203),
.A2(n_1827),
.B(n_1828),
.Y(n_2893)
);

AOI21x1_ASAP7_75t_L g2894 ( 
.A1(n_2420),
.A2(n_2311),
.B(n_2593),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2303),
.B(n_1946),
.Y(n_2895)
);

BUFx3_ASAP7_75t_L g2896 ( 
.A(n_2251),
.Y(n_2896)
);

AOI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2533),
.A2(n_1700),
.B(n_1588),
.Y(n_2897)
);

NOR2x1_ASAP7_75t_L g2898 ( 
.A(n_2330),
.B(n_2052),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_SL g2899 ( 
.A(n_2556),
.B(n_1952),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2303),
.B(n_1921),
.Y(n_2900)
);

OR2x6_ASAP7_75t_L g2901 ( 
.A(n_2224),
.B(n_1545),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2298),
.B(n_1921),
.Y(n_2902)
);

AOI21xp5_ASAP7_75t_L g2903 ( 
.A1(n_2533),
.A2(n_1724),
.B(n_1700),
.Y(n_2903)
);

A2O1A1Ixp33_ASAP7_75t_L g2904 ( 
.A1(n_2220),
.A2(n_1980),
.B(n_1989),
.C(n_2062),
.Y(n_2904)
);

A2O1A1Ixp33_ASAP7_75t_SL g2905 ( 
.A1(n_2449),
.A2(n_2014),
.B(n_2005),
.C(n_2025),
.Y(n_2905)
);

AOI21xp5_ASAP7_75t_L g2906 ( 
.A1(n_2546),
.A2(n_1757),
.B(n_1724),
.Y(n_2906)
);

NAND3xp33_ASAP7_75t_L g2907 ( 
.A(n_2220),
.B(n_1849),
.C(n_1845),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_2726),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2174),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2382),
.A2(n_2607),
.B1(n_2214),
.B2(n_2217),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2320),
.B(n_2342),
.Y(n_2911)
);

BUFx12f_ASAP7_75t_L g2912 ( 
.A(n_2469),
.Y(n_2912)
);

BUFx6f_ASAP7_75t_L g2913 ( 
.A(n_2530),
.Y(n_2913)
);

HB1xp67_ASAP7_75t_L g2914 ( 
.A(n_2252),
.Y(n_2914)
);

OAI22xp5_ASAP7_75t_L g2915 ( 
.A1(n_2607),
.A2(n_2214),
.B1(n_2217),
.B2(n_2197),
.Y(n_2915)
);

INVxp67_ASAP7_75t_L g2916 ( 
.A(n_2522),
.Y(n_2916)
);

AOI21xp5_ASAP7_75t_L g2917 ( 
.A1(n_2546),
.A2(n_2569),
.B(n_2561),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2569),
.A2(n_2497),
.B(n_2496),
.Y(n_2918)
);

NOR2xp33_ASAP7_75t_L g2919 ( 
.A(n_2342),
.B(n_1852),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2346),
.B(n_1909),
.Y(n_2920)
);

BUFx2_ASAP7_75t_L g2921 ( 
.A(n_2401),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2174),
.Y(n_2922)
);

NAND2xp5_ASAP7_75t_L g2923 ( 
.A(n_2346),
.B(n_1913),
.Y(n_2923)
);

OAI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2197),
.A2(n_2048),
.B1(n_1828),
.B2(n_1998),
.Y(n_2924)
);

INVx2_ASAP7_75t_L g2925 ( 
.A(n_2489),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2347),
.B(n_1931),
.Y(n_2926)
);

BUFx6f_ASAP7_75t_L g2927 ( 
.A(n_2530),
.Y(n_2927)
);

BUFx2_ASAP7_75t_L g2928 ( 
.A(n_2401),
.Y(n_2928)
);

OAI21x1_ASAP7_75t_L g2929 ( 
.A1(n_2794),
.A2(n_1935),
.B(n_1985),
.Y(n_2929)
);

BUFx6f_ASAP7_75t_L g2930 ( 
.A(n_2530),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2347),
.B(n_1980),
.Y(n_2931)
);

OAI22x1_ASAP7_75t_L g2932 ( 
.A1(n_2593),
.A2(n_1989),
.B1(n_2009),
.B2(n_1986),
.Y(n_2932)
);

AOI22xp33_ASAP7_75t_L g2933 ( 
.A1(n_2242),
.A2(n_1912),
.B1(n_1875),
.B2(n_1587),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_2355),
.B(n_1954),
.Y(n_2934)
);

OAI21xp5_ASAP7_75t_L g2935 ( 
.A1(n_2290),
.A2(n_2069),
.B(n_2060),
.Y(n_2935)
);

AO32x2_ASAP7_75t_L g2936 ( 
.A1(n_2429),
.A2(n_2471),
.A3(n_2457),
.B1(n_2570),
.B2(n_2504),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2556),
.B(n_1992),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2508),
.A2(n_2142),
.B(n_1945),
.Y(n_2938)
);

BUFx2_ASAP7_75t_L g2939 ( 
.A(n_2401),
.Y(n_2939)
);

OR2x2_ASAP7_75t_L g2940 ( 
.A(n_2294),
.B(n_2011),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2527),
.A2(n_2154),
.B(n_2142),
.Y(n_2941)
);

NOR2xp33_ASAP7_75t_SL g2942 ( 
.A(n_2169),
.B(n_1545),
.Y(n_2942)
);

OAI21xp5_ASAP7_75t_L g2943 ( 
.A1(n_2290),
.A2(n_2244),
.B(n_2242),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2355),
.B(n_1987),
.Y(n_2944)
);

BUFx6f_ASAP7_75t_L g2945 ( 
.A(n_2535),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2388),
.B(n_1954),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2193),
.Y(n_2947)
);

AOI21xp5_ASAP7_75t_L g2948 ( 
.A1(n_2527),
.A2(n_2154),
.B(n_2142),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2388),
.B(n_1906),
.Y(n_2949)
);

AOI21xp5_ASAP7_75t_L g2950 ( 
.A1(n_2763),
.A2(n_1810),
.B(n_1537),
.Y(n_2950)
);

AOI22xp33_ASAP7_75t_L g2951 ( 
.A1(n_2244),
.A2(n_1587),
.B1(n_1992),
.B2(n_2023),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2193),
.Y(n_2952)
);

AOI21xp5_ASAP7_75t_L g2953 ( 
.A1(n_2763),
.A2(n_1810),
.B(n_1537),
.Y(n_2953)
);

OR2x2_ASAP7_75t_L g2954 ( 
.A(n_2294),
.B(n_2011),
.Y(n_2954)
);

INVx2_ASAP7_75t_L g2955 ( 
.A(n_2489),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2193),
.Y(n_2956)
);

AOI21xp5_ASAP7_75t_L g2957 ( 
.A1(n_2763),
.A2(n_1810),
.B(n_1537),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2763),
.A2(n_1850),
.B(n_1798),
.Y(n_2958)
);

HB1xp67_ASAP7_75t_L g2959 ( 
.A(n_2262),
.Y(n_2959)
);

AND2x2_ASAP7_75t_L g2960 ( 
.A(n_2539),
.B(n_1906),
.Y(n_2960)
);

AOI21xp5_ASAP7_75t_L g2961 ( 
.A1(n_2763),
.A2(n_1850),
.B(n_1798),
.Y(n_2961)
);

A2O1A1Ixp33_ASAP7_75t_L g2962 ( 
.A1(n_2311),
.A2(n_2073),
.B(n_2068),
.C(n_2064),
.Y(n_2962)
);

AOI21x1_ASAP7_75t_L g2963 ( 
.A1(n_2420),
.A2(n_1996),
.B(n_2022),
.Y(n_2963)
);

OAI21xp5_ASAP7_75t_L g2964 ( 
.A1(n_2183),
.A2(n_2186),
.B(n_2715),
.Y(n_2964)
);

BUFx12f_ASAP7_75t_L g2965 ( 
.A(n_2469),
.Y(n_2965)
);

O2A1O1Ixp33_ASAP7_75t_SL g2966 ( 
.A1(n_2189),
.A2(n_2001),
.B(n_2006),
.C(n_2008),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_SL g2967 ( 
.A(n_2685),
.B(n_2270),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2802),
.B(n_1906),
.Y(n_2968)
);

INVx1_ASAP7_75t_SL g2969 ( 
.A(n_2720),
.Y(n_2969)
);

AOI21xp5_ASAP7_75t_L g2970 ( 
.A1(n_2763),
.A2(n_1850),
.B(n_1798),
.Y(n_2970)
);

AOI21x1_ASAP7_75t_L g2971 ( 
.A1(n_2420),
.A2(n_2075),
.B(n_2065),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_SL g2972 ( 
.A(n_2685),
.B(n_2023),
.Y(n_2972)
);

O2A1O1Ixp33_ASAP7_75t_L g2973 ( 
.A1(n_2183),
.A2(n_2001),
.B(n_2006),
.C(n_2008),
.Y(n_2973)
);

NOR2xp33_ASAP7_75t_L g2974 ( 
.A(n_2538),
.B(n_2039),
.Y(n_2974)
);

INVx3_ASAP7_75t_L g2975 ( 
.A(n_2726),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2193),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2199),
.Y(n_2977)
);

AOI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2186),
.A2(n_2449),
.B1(n_2270),
.B2(n_2279),
.Y(n_2978)
);

A2O1A1Ixp33_ASAP7_75t_L g2979 ( 
.A1(n_2715),
.A2(n_2073),
.B(n_2034),
.C(n_2023),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2802),
.B(n_1914),
.Y(n_2980)
);

BUFx2_ASAP7_75t_L g2981 ( 
.A(n_2401),
.Y(n_2981)
);

AOI21xp5_ASAP7_75t_L g2982 ( 
.A1(n_2756),
.A2(n_2592),
.B(n_2736),
.Y(n_2982)
);

O2A1O1Ixp5_ASAP7_75t_L g2983 ( 
.A1(n_2592),
.A2(n_2063),
.B(n_2078),
.C(n_2053),
.Y(n_2983)
);

AOI21xp5_ASAP7_75t_L g2984 ( 
.A1(n_2756),
.A2(n_1850),
.B(n_2098),
.Y(n_2984)
);

AO21x1_ASAP7_75t_L g2985 ( 
.A1(n_2647),
.A2(n_2045),
.B(n_2010),
.Y(n_2985)
);

AOI21xp5_ASAP7_75t_L g2986 ( 
.A1(n_2756),
.A2(n_1616),
.B(n_2098),
.Y(n_2986)
);

OAI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2460),
.A2(n_1998),
.B1(n_1978),
.B2(n_1698),
.Y(n_2987)
);

AOI21xp5_ASAP7_75t_L g2988 ( 
.A1(n_2756),
.A2(n_2736),
.B(n_2615),
.Y(n_2988)
);

OAI22xp5_ASAP7_75t_SL g2989 ( 
.A1(n_2476),
.A2(n_2017),
.B1(n_2034),
.B2(n_2021),
.Y(n_2989)
);

BUFx2_ASAP7_75t_L g2990 ( 
.A(n_2401),
.Y(n_2990)
);

AOI21xp5_ASAP7_75t_L g2991 ( 
.A1(n_2756),
.A2(n_2098),
.B(n_1953),
.Y(n_2991)
);

HB1xp67_ASAP7_75t_L g2992 ( 
.A(n_2262),
.Y(n_2992)
);

BUFx2_ASAP7_75t_L g2993 ( 
.A(n_2401),
.Y(n_2993)
);

INVx2_ASAP7_75t_L g2994 ( 
.A(n_2489),
.Y(n_2994)
);

AOI21xp33_ASAP7_75t_L g2995 ( 
.A1(n_2279),
.A2(n_2069),
.B(n_2060),
.Y(n_2995)
);

OAI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2460),
.A2(n_1978),
.B1(n_1698),
.B2(n_1785),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2199),
.Y(n_2997)
);

NOR2xp33_ASAP7_75t_L g2998 ( 
.A(n_2538),
.B(n_2039),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_L g2999 ( 
.A(n_2676),
.B(n_1914),
.Y(n_2999)
);

OAI22xp5_ASAP7_75t_L g3000 ( 
.A1(n_2445),
.A2(n_1978),
.B1(n_1918),
.B2(n_1698),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2199),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2160),
.Y(n_3002)
);

BUFx2_ASAP7_75t_L g3003 ( 
.A(n_2401),
.Y(n_3003)
);

AND2x2_ASAP7_75t_SL g3004 ( 
.A(n_2163),
.B(n_1545),
.Y(n_3004)
);

BUFx3_ASAP7_75t_L g3005 ( 
.A(n_2251),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2199),
.Y(n_3006)
);

OAI22xp5_ASAP7_75t_L g3007 ( 
.A1(n_2445),
.A2(n_1545),
.B1(n_1918),
.B2(n_1785),
.Y(n_3007)
);

NOR2x1p5_ASAP7_75t_SL g3008 ( 
.A(n_2794),
.B(n_1587),
.Y(n_3008)
);

BUFx8_ASAP7_75t_L g3009 ( 
.A(n_2431),
.Y(n_3009)
);

NOR3xp33_ASAP7_75t_L g3010 ( 
.A(n_2441),
.B(n_2040),
.C(n_2046),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2547),
.B(n_2040),
.Y(n_3011)
);

OAI22xp5_ASAP7_75t_L g3012 ( 
.A1(n_2328),
.A2(n_1918),
.B1(n_1785),
.B2(n_1698),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_2676),
.B(n_1914),
.Y(n_3013)
);

AOI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2328),
.A2(n_2468),
.B1(n_2441),
.B2(n_2547),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_SL g3015 ( 
.A(n_2649),
.B(n_1587),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2424),
.B(n_1923),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2424),
.B(n_1923),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2495),
.B(n_1923),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2201),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2201),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_L g3021 ( 
.A(n_2495),
.B(n_1900),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_SL g3022 ( 
.A(n_2649),
.B(n_1587),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2499),
.B(n_1787),
.Y(n_3023)
);

NAND3xp33_ASAP7_75t_L g3024 ( 
.A(n_2468),
.B(n_2059),
.C(n_1841),
.Y(n_3024)
);

INVx2_ASAP7_75t_SL g3025 ( 
.A(n_2737),
.Y(n_3025)
);

INVx2_ASAP7_75t_L g3026 ( 
.A(n_2201),
.Y(n_3026)
);

A2O1A1Ixp33_ASAP7_75t_L g3027 ( 
.A1(n_2328),
.A2(n_1878),
.B(n_1787),
.C(n_2017),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2336),
.B(n_1900),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2201),
.Y(n_3029)
);

CKINVDCx11_ASAP7_75t_R g3030 ( 
.A(n_2418),
.Y(n_3030)
);

AOI21xp5_ASAP7_75t_L g3031 ( 
.A1(n_2545),
.A2(n_2586),
.B(n_2165),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2209),
.Y(n_3032)
);

AND2x2_ASAP7_75t_L g3033 ( 
.A(n_2539),
.B(n_1645),
.Y(n_3033)
);

NOR2xp33_ASAP7_75t_L g3034 ( 
.A(n_2375),
.B(n_2046),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2603),
.B(n_1645),
.Y(n_3035)
);

AO21x1_ASAP7_75t_L g3036 ( 
.A1(n_2647),
.A2(n_2045),
.B(n_2010),
.Y(n_3036)
);

OAI22xp5_ASAP7_75t_L g3037 ( 
.A1(n_2169),
.A2(n_1918),
.B1(n_1785),
.B2(n_1843),
.Y(n_3037)
);

OAI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_2169),
.A2(n_1829),
.B1(n_1830),
.B2(n_1834),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2209),
.Y(n_3039)
);

BUFx6f_ASAP7_75t_L g3040 ( 
.A(n_2535),
.Y(n_3040)
);

OR2x6_ASAP7_75t_L g3041 ( 
.A(n_2224),
.B(n_2033),
.Y(n_3041)
);

BUFx2_ASAP7_75t_SL g3042 ( 
.A(n_2169),
.Y(n_3042)
);

OAI21xp5_ASAP7_75t_L g3043 ( 
.A1(n_2397),
.A2(n_2059),
.B(n_2066),
.Y(n_3043)
);

BUFx4f_ASAP7_75t_L g3044 ( 
.A(n_2227),
.Y(n_3044)
);

BUFx4f_ASAP7_75t_L g3045 ( 
.A(n_2227),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_2336),
.B(n_1547),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_L g3047 ( 
.A(n_2337),
.B(n_1549),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_L g3048 ( 
.A(n_2337),
.B(n_1549),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2209),
.Y(n_3049)
);

O2A1O1Ixp5_ASAP7_75t_L g3050 ( 
.A1(n_2481),
.A2(n_2058),
.B(n_2053),
.C(n_2054),
.Y(n_3050)
);

HB1xp67_ASAP7_75t_L g3051 ( 
.A(n_2354),
.Y(n_3051)
);

CKINVDCx14_ASAP7_75t_R g3052 ( 
.A(n_2194),
.Y(n_3052)
);

AND2x2_ASAP7_75t_L g3053 ( 
.A(n_2603),
.B(n_1645),
.Y(n_3053)
);

BUFx8_ASAP7_75t_SL g3054 ( 
.A(n_2232),
.Y(n_3054)
);

AOI21x1_ASAP7_75t_L g3055 ( 
.A1(n_2446),
.A2(n_1878),
.B(n_2015),
.Y(n_3055)
);

AOI22xp5_ASAP7_75t_L g3056 ( 
.A1(n_2406),
.A2(n_2066),
.B1(n_2054),
.B2(n_2058),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_SL g3057 ( 
.A(n_2499),
.B(n_1950),
.Y(n_3057)
);

A2O1A1Ixp33_ASAP7_75t_L g3058 ( 
.A1(n_2476),
.A2(n_2038),
.B(n_2050),
.C(n_1988),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_2209),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2485),
.B(n_1549),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_SL g3061 ( 
.A(n_2745),
.B(n_1950),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_2213),
.Y(n_3062)
);

AOI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2586),
.A2(n_2098),
.B(n_1953),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_2603),
.B(n_1652),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_L g3065 ( 
.A(n_2485),
.B(n_1565),
.Y(n_3065)
);

A2O1A1Ixp33_ASAP7_75t_L g3066 ( 
.A1(n_2326),
.A2(n_2038),
.B(n_2050),
.C(n_2020),
.Y(n_3066)
);

OAI21xp5_ASAP7_75t_L g3067 ( 
.A1(n_2397),
.A2(n_2066),
.B(n_1982),
.Y(n_3067)
);

BUFx6f_ASAP7_75t_L g3068 ( 
.A(n_2535),
.Y(n_3068)
);

NOR2xp33_ASAP7_75t_SL g3069 ( 
.A(n_2179),
.B(n_1616),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2375),
.B(n_1712),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2500),
.B(n_2453),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2745),
.B(n_1950),
.Y(n_3072)
);

AOI21xp5_ASAP7_75t_L g3073 ( 
.A1(n_2165),
.A2(n_2170),
.B(n_2529),
.Y(n_3073)
);

NAND2x1p5_ASAP7_75t_L g3074 ( 
.A(n_2179),
.B(n_1616),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2751),
.B(n_1950),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_2213),
.Y(n_3076)
);

BUFx3_ASAP7_75t_L g3077 ( 
.A(n_2251),
.Y(n_3077)
);

OAI22xp5_ASAP7_75t_L g3078 ( 
.A1(n_2179),
.A2(n_1855),
.B1(n_1829),
.B2(n_1830),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_L g3079 ( 
.A1(n_2165),
.A2(n_2170),
.B(n_2529),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_2751),
.B(n_1950),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2500),
.B(n_1565),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2165),
.A2(n_2170),
.B(n_2529),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2213),
.Y(n_3083)
);

OAI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2179),
.A2(n_1843),
.B1(n_1836),
.B2(n_1855),
.Y(n_3084)
);

OR2x6_ASAP7_75t_L g3085 ( 
.A(n_2224),
.B(n_2033),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2218),
.Y(n_3086)
);

OAI22x1_ASAP7_75t_L g3087 ( 
.A1(n_2282),
.A2(n_2020),
.B1(n_2013),
.B2(n_2015),
.Y(n_3087)
);

A2O1A1Ixp33_ASAP7_75t_SL g3088 ( 
.A1(n_2531),
.A2(n_1907),
.B(n_1979),
.C(n_1982),
.Y(n_3088)
);

INVx2_ASAP7_75t_L g3089 ( 
.A(n_2218),
.Y(n_3089)
);

AOI21xp5_ASAP7_75t_L g3090 ( 
.A1(n_2170),
.A2(n_1907),
.B(n_2033),
.Y(n_3090)
);

AOI21xp5_ASAP7_75t_L g3091 ( 
.A1(n_2678),
.A2(n_1907),
.B(n_2033),
.Y(n_3091)
);

A2O1A1Ixp33_ASAP7_75t_L g3092 ( 
.A1(n_2326),
.A2(n_2024),
.B(n_2013),
.C(n_2021),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2453),
.B(n_1565),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2726),
.Y(n_3094)
);

NOR2xp33_ASAP7_75t_L g3095 ( 
.A(n_2216),
.B(n_1736),
.Y(n_3095)
);

O2A1O1Ixp33_ASAP7_75t_L g3096 ( 
.A1(n_2282),
.A2(n_2024),
.B(n_2036),
.C(n_1964),
.Y(n_3096)
);

BUFx2_ASAP7_75t_L g3097 ( 
.A(n_2401),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2416),
.A2(n_2035),
.B1(n_2071),
.B2(n_2016),
.Y(n_3098)
);

NAND2xp5_ASAP7_75t_SL g3099 ( 
.A(n_2735),
.B(n_1950),
.Y(n_3099)
);

OAI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2481),
.A2(n_2004),
.B(n_1979),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2218),
.Y(n_3101)
);

AOI21xp5_ASAP7_75t_L g3102 ( 
.A1(n_2678),
.A2(n_2681),
.B(n_2447),
.Y(n_3102)
);

OAI22xp5_ASAP7_75t_L g3103 ( 
.A1(n_2179),
.A2(n_2282),
.B1(n_2783),
.B2(n_2249),
.Y(n_3103)
);

OR2x2_ASAP7_75t_L g3104 ( 
.A(n_2212),
.B(n_1925),
.Y(n_3104)
);

AOI21xp5_ASAP7_75t_L g3105 ( 
.A1(n_2681),
.A2(n_2033),
.B(n_2036),
.Y(n_3105)
);

AND2x2_ASAP7_75t_L g3106 ( 
.A(n_2507),
.B(n_1794),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2218),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_2305),
.B(n_1568),
.Y(n_3108)
);

AOI21xp5_ASAP7_75t_L g3109 ( 
.A1(n_2447),
.A2(n_2608),
.B(n_2601),
.Y(n_3109)
);

HB1xp67_ASAP7_75t_L g3110 ( 
.A(n_2354),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2305),
.B(n_1568),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_2447),
.A2(n_1951),
.B(n_2029),
.Y(n_3112)
);

AOI21xp33_ASAP7_75t_L g3113 ( 
.A1(n_2459),
.A2(n_2035),
.B(n_1964),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2507),
.B(n_1794),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_SL g3115 ( 
.A(n_2179),
.B(n_2029),
.Y(n_3115)
);

A2O1A1Ixp33_ASAP7_75t_L g3116 ( 
.A1(n_2735),
.A2(n_1975),
.B(n_2061),
.C(n_1995),
.Y(n_3116)
);

O2A1O1Ixp33_ASAP7_75t_L g3117 ( 
.A1(n_2282),
.A2(n_1995),
.B(n_2079),
.C(n_2074),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2312),
.B(n_1568),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2251),
.Y(n_3119)
);

CKINVDCx20_ASAP7_75t_R g3120 ( 
.A(n_2194),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2312),
.B(n_1569),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2216),
.B(n_1736),
.Y(n_3122)
);

OR2x6_ASAP7_75t_L g3123 ( 
.A(n_2224),
.B(n_1957),
.Y(n_3123)
);

BUFx4f_ASAP7_75t_L g3124 ( 
.A(n_2227),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2226),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2226),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2451),
.B(n_1569),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_2447),
.A2(n_2608),
.B(n_2601),
.Y(n_3128)
);

INVx1_ASAP7_75t_L g3129 ( 
.A(n_2226),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2451),
.B(n_1569),
.Y(n_3130)
);

BUFx6f_ASAP7_75t_L g3131 ( 
.A(n_2535),
.Y(n_3131)
);

AOI22xp5_ASAP7_75t_L g3132 ( 
.A1(n_2416),
.A2(n_1982),
.B1(n_2071),
.B2(n_2057),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2226),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_L g3134 ( 
.A(n_2584),
.Y(n_3134)
);

O2A1O1Ixp33_ASAP7_75t_L g3135 ( 
.A1(n_2505),
.A2(n_2793),
.B(n_2722),
.C(n_2267),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2229),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2559),
.B(n_1572),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2559),
.B(n_1572),
.Y(n_3138)
);

AOI22xp33_ASAP7_75t_L g3139 ( 
.A1(n_2335),
.A2(n_2071),
.B1(n_2057),
.B2(n_2056),
.Y(n_3139)
);

OA22x2_ASAP7_75t_L g3140 ( 
.A1(n_2759),
.A2(n_2079),
.B1(n_2074),
.B2(n_2057),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2735),
.B(n_1951),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2714),
.B(n_1572),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2229),
.Y(n_3143)
);

NOR2xp33_ASAP7_75t_R g3144 ( 
.A(n_2712),
.B(n_2029),
.Y(n_3144)
);

OR2x6_ASAP7_75t_L g3145 ( 
.A(n_2224),
.B(n_1957),
.Y(n_3145)
);

NOR3xp33_ASAP7_75t_L g3146 ( 
.A(n_2505),
.B(n_1834),
.C(n_1840),
.Y(n_3146)
);

INVxp67_ASAP7_75t_L g3147 ( 
.A(n_2638),
.Y(n_3147)
);

INVx1_ASAP7_75t_L g3148 ( 
.A(n_2229),
.Y(n_3148)
);

OAI21xp5_ASAP7_75t_L g3149 ( 
.A1(n_2531),
.A2(n_2056),
.B(n_1979),
.Y(n_3149)
);

BUFx12f_ASAP7_75t_L g3150 ( 
.A(n_2512),
.Y(n_3150)
);

OAI21xp33_ASAP7_75t_SL g3151 ( 
.A1(n_2163),
.A2(n_2173),
.B(n_2172),
.Y(n_3151)
);

OAI22xp5_ASAP7_75t_L g3152 ( 
.A1(n_2179),
.A2(n_1854),
.B1(n_1847),
.B2(n_1841),
.Y(n_3152)
);

AOI21xp5_ASAP7_75t_L g3153 ( 
.A1(n_2618),
.A2(n_2623),
.B(n_2620),
.Y(n_3153)
);

NAND2xp5_ASAP7_75t_L g3154 ( 
.A(n_2714),
.B(n_2435),
.Y(n_3154)
);

NAND2x1p5_ASAP7_75t_L g3155 ( 
.A(n_2179),
.B(n_1957),
.Y(n_3155)
);

AND2x2_ASAP7_75t_L g3156 ( 
.A(n_2507),
.B(n_1783),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2618),
.A2(n_2623),
.B(n_2620),
.Y(n_3157)
);

AO21x1_ASAP7_75t_L g3158 ( 
.A1(n_2463),
.A2(n_2032),
.B(n_2047),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_SL g3159 ( 
.A(n_2759),
.B(n_1951),
.Y(n_3159)
);

AOI21xp5_ASAP7_75t_L g3160 ( 
.A1(n_2631),
.A2(n_2029),
.B(n_1951),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2435),
.B(n_1596),
.Y(n_3161)
);

INVx3_ASAP7_75t_L g3162 ( 
.A(n_2726),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2236),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2236),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2690),
.B(n_1836),
.Y(n_3165)
);

A2O1A1Ixp33_ASAP7_75t_L g3166 ( 
.A1(n_2463),
.A2(n_2459),
.B(n_2793),
.C(n_2722),
.Y(n_3166)
);

OAI22xp5_ASAP7_75t_L g3167 ( 
.A1(n_2783),
.A2(n_1854),
.B1(n_1847),
.B2(n_1840),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_2439),
.B(n_1596),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_2631),
.A2(n_2032),
.B(n_2047),
.Y(n_3169)
);

AOI21xp5_ASAP7_75t_L g3170 ( 
.A1(n_2633),
.A2(n_2032),
.B(n_2047),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2439),
.B(n_2440),
.Y(n_3171)
);

AND2x4_ASAP7_75t_L g3172 ( 
.A(n_2168),
.B(n_1984),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2440),
.B(n_1596),
.Y(n_3173)
);

OA22x2_ASAP7_75t_L g3174 ( 
.A1(n_2690),
.A2(n_2056),
.B1(n_2042),
.B2(n_2041),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2444),
.B(n_1618),
.Y(n_3175)
);

AND2x2_ASAP7_75t_L g3176 ( 
.A(n_2510),
.B(n_1765),
.Y(n_3176)
);

O2A1O1Ixp33_ASAP7_75t_L g3177 ( 
.A1(n_2267),
.A2(n_2042),
.B(n_2041),
.C(n_2016),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2510),
.B(n_1765),
.Y(n_3178)
);

AO21x1_ASAP7_75t_L g3179 ( 
.A1(n_2172),
.A2(n_2047),
.B(n_1928),
.Y(n_3179)
);

AOI33xp33_ASAP7_75t_L g3180 ( 
.A1(n_2524),
.A2(n_2042),
.A3(n_2041),
.B1(n_2016),
.B2(n_2004),
.B3(n_1984),
.Y(n_3180)
);

NOR2xp67_ASAP7_75t_L g3181 ( 
.A(n_2234),
.B(n_1984),
.Y(n_3181)
);

NAND2xp5_ASAP7_75t_L g3182 ( 
.A(n_2444),
.B(n_1618),
.Y(n_3182)
);

BUFx4f_ASAP7_75t_SL g3183 ( 
.A(n_2431),
.Y(n_3183)
);

O2A1O1Ixp33_ASAP7_75t_L g3184 ( 
.A1(n_2483),
.A2(n_2004),
.B(n_1632),
.C(n_1633),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2245),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2483),
.B(n_1618),
.Y(n_3186)
);

AOI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_2633),
.A2(n_1737),
.B(n_1794),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2634),
.A2(n_1695),
.B(n_1783),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2634),
.A2(n_1695),
.B(n_1783),
.Y(n_3189)
);

AOI221xp5_ASAP7_75t_L g3190 ( 
.A1(n_2249),
.A2(n_1632),
.B1(n_1633),
.B2(n_1636),
.C(n_1642),
.Y(n_3190)
);

INVx4_ASAP7_75t_L g3191 ( 
.A(n_2246),
.Y(n_3191)
);

INVxp67_ASAP7_75t_SL g3192 ( 
.A(n_2172),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2645),
.A2(n_1695),
.B(n_1782),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2245),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2654),
.B(n_1632),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2245),
.Y(n_3196)
);

AO22x1_ASAP7_75t_L g3197 ( 
.A1(n_2189),
.A2(n_1636),
.B1(n_1642),
.B2(n_2141),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2654),
.B(n_1636),
.Y(n_3198)
);

AO21x1_ASAP7_75t_L g3199 ( 
.A1(n_2173),
.A2(n_1642),
.B(n_2141),
.Y(n_3199)
);

NOR2xp33_ASAP7_75t_L g3200 ( 
.A(n_2670),
.B(n_2152),
.Y(n_3200)
);

AOI21xp5_ASAP7_75t_L g3201 ( 
.A1(n_2645),
.A2(n_1652),
.B(n_1656),
.Y(n_3201)
);

OR2x6_ASAP7_75t_SL g3202 ( 
.A(n_2581),
.B(n_2646),
.Y(n_3202)
);

O2A1O1Ixp5_ASAP7_75t_L g3203 ( 
.A1(n_2718),
.A2(n_2152),
.B(n_2141),
.C(n_2129),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_SL g3204 ( 
.A(n_2541),
.B(n_2799),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2737),
.Y(n_3205)
);

OR2x2_ASAP7_75t_L g3206 ( 
.A(n_2212),
.B(n_1652),
.Y(n_3206)
);

OA22x2_ASAP7_75t_L g3207 ( 
.A1(n_2799),
.A2(n_2152),
.B1(n_2129),
.B2(n_1660),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_L g3208 ( 
.A(n_2670),
.B(n_2129),
.Y(n_3208)
);

AOI22xp5_ASAP7_75t_L g3209 ( 
.A1(n_2524),
.A2(n_1656),
.B1(n_1658),
.B2(n_1660),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2661),
.A2(n_1656),
.B(n_1658),
.Y(n_3210)
);

NOR2xp33_ASAP7_75t_L g3211 ( 
.A(n_2732),
.B(n_1658),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2576),
.B(n_1660),
.Y(n_3212)
);

BUFx4f_ASAP7_75t_L g3213 ( 
.A(n_2227),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_2541),
.B(n_1665),
.Y(n_3214)
);

AOI21xp5_ASAP7_75t_L g3215 ( 
.A1(n_2661),
.A2(n_1665),
.B(n_1673),
.Y(n_3215)
);

CKINVDCx20_ASAP7_75t_R g3216 ( 
.A(n_2532),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_SL g3217 ( 
.A(n_2335),
.B(n_1673),
.Y(n_3217)
);

AND2x2_ASAP7_75t_L g3218 ( 
.A(n_2510),
.B(n_1676),
.Y(n_3218)
);

AOI21xp5_ASAP7_75t_L g3219 ( 
.A1(n_2662),
.A2(n_1676),
.B(n_1737),
.Y(n_3219)
);

INVx2_ASAP7_75t_L g3220 ( 
.A(n_2245),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2576),
.B(n_1744),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_2249),
.A2(n_1744),
.B1(n_1754),
.B2(n_1765),
.Y(n_3222)
);

INVxp67_ASAP7_75t_SL g3223 ( 
.A(n_2173),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2260),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_2335),
.B(n_1754),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_2589),
.B(n_1766),
.Y(n_3226)
);

AOI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_2666),
.A2(n_1766),
.B(n_1780),
.Y(n_3227)
);

AND2x2_ASAP7_75t_L g3228 ( 
.A(n_2163),
.B(n_1766),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_2589),
.B(n_1780),
.Y(n_3229)
);

A2O1A1Ixp33_ASAP7_75t_L g3230 ( 
.A1(n_2459),
.A2(n_1782),
.B(n_2163),
.C(n_2351),
.Y(n_3230)
);

OAI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_2249),
.A2(n_2178),
.B1(n_2175),
.B2(n_2731),
.Y(n_3231)
);

INVx2_ASAP7_75t_SL g3232 ( 
.A(n_2737),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_2249),
.B(n_2299),
.Y(n_3233)
);

AOI21xp5_ASAP7_75t_L g3234 ( 
.A1(n_2484),
.A2(n_2776),
.B(n_2806),
.Y(n_3234)
);

O2A1O1Ixp33_ASAP7_75t_L g3235 ( 
.A1(n_2806),
.A2(n_2638),
.B(n_2228),
.C(n_2732),
.Y(n_3235)
);

AND2x4_ASAP7_75t_L g3236 ( 
.A(n_2168),
.B(n_2239),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2639),
.B(n_2686),
.Y(n_3237)
);

INVx3_ASAP7_75t_SL g3238 ( 
.A(n_2646),
.Y(n_3238)
);

OAI22xp5_ASAP7_75t_L g3239 ( 
.A1(n_2249),
.A2(n_2178),
.B1(n_2175),
.B2(n_2731),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_SL g3240 ( 
.A(n_2335),
.B(n_2361),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2584),
.Y(n_3241)
);

OR2x6_ASAP7_75t_L g3242 ( 
.A(n_2224),
.B(n_2365),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2639),
.B(n_2686),
.Y(n_3243)
);

AND2x2_ASAP7_75t_L g3244 ( 
.A(n_2249),
.B(n_2299),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_L g3245 ( 
.A(n_2672),
.B(n_2659),
.Y(n_3245)
);

AOI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2484),
.A2(n_2776),
.B(n_2224),
.Y(n_3246)
);

AOI22xp5_ASAP7_75t_L g3247 ( 
.A1(n_2351),
.A2(n_2361),
.B1(n_2335),
.B2(n_2672),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_SL g3248 ( 
.A(n_2335),
.B(n_2361),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2776),
.A2(n_2365),
.B(n_2702),
.Y(n_3249)
);

O2A1O1Ixp33_ASAP7_75t_L g3250 ( 
.A1(n_2228),
.A2(n_2362),
.B(n_2188),
.C(n_2222),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2696),
.B(n_2659),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_SL g3252 ( 
.A(n_2361),
.B(n_2704),
.Y(n_3252)
);

OAI22xp5_ASAP7_75t_L g3253 ( 
.A1(n_2175),
.A2(n_2178),
.B1(n_2731),
.B2(n_2717),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_2776),
.A2(n_2365),
.B(n_2702),
.Y(n_3254)
);

NAND3xp33_ASAP7_75t_L g3255 ( 
.A(n_2773),
.B(n_2771),
.C(n_2351),
.Y(n_3255)
);

NOR2xp33_ASAP7_75t_L g3256 ( 
.A(n_2512),
.B(n_2281),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2260),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2696),
.B(n_2697),
.Y(n_3258)
);

AOI21xp5_ASAP7_75t_L g3259 ( 
.A1(n_2776),
.A2(n_2365),
.B(n_2343),
.Y(n_3259)
);

NOR3xp33_ASAP7_75t_L g3260 ( 
.A(n_2718),
.B(n_2660),
.C(n_2653),
.Y(n_3260)
);

AO21x1_ASAP7_75t_L g3261 ( 
.A1(n_2181),
.A2(n_2184),
.B(n_2182),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_2365),
.A2(n_2343),
.B(n_2246),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_2365),
.A2(n_2343),
.B(n_2246),
.Y(n_3263)
);

BUFx6f_ASAP7_75t_L g3264 ( 
.A(n_2584),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2697),
.B(n_2598),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_SL g3266 ( 
.A(n_2361),
.B(n_2704),
.Y(n_3266)
);

A2O1A1Ixp33_ASAP7_75t_L g3267 ( 
.A1(n_2516),
.A2(n_2622),
.B(n_2361),
.C(n_2509),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2598),
.B(n_2752),
.Y(n_3268)
);

AOI22xp5_ASAP7_75t_L g3269 ( 
.A1(n_2766),
.A2(n_2295),
.B1(n_2472),
.B2(n_2434),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_SL g3270 ( 
.A(n_2516),
.B(n_2430),
.Y(n_3270)
);

OA22x2_ASAP7_75t_L g3271 ( 
.A1(n_2602),
.A2(n_2177),
.B1(n_2660),
.B2(n_2653),
.Y(n_3271)
);

AOI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_2365),
.A2(n_2343),
.B(n_2246),
.Y(n_3272)
);

O2A1O1Ixp5_ASAP7_75t_SL g3273 ( 
.A1(n_2210),
.A2(n_2233),
.B(n_2164),
.C(n_2393),
.Y(n_3273)
);

HB1xp67_ASAP7_75t_L g3274 ( 
.A(n_2362),
.Y(n_3274)
);

AOI21xp5_ASAP7_75t_L g3275 ( 
.A1(n_2246),
.A2(n_2511),
.B(n_2343),
.Y(n_3275)
);

O2A1O1Ixp33_ASAP7_75t_SL g3276 ( 
.A1(n_2177),
.A2(n_2766),
.B(n_2809),
.C(n_2418),
.Y(n_3276)
);

BUFx3_ASAP7_75t_L g3277 ( 
.A(n_2251),
.Y(n_3277)
);

AOI21x1_ASAP7_75t_L g3278 ( 
.A1(n_2446),
.A2(n_2456),
.B(n_2718),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2265),
.Y(n_3279)
);

NOR3xp33_ASAP7_75t_L g3280 ( 
.A(n_2653),
.B(n_2660),
.C(n_2302),
.Y(n_3280)
);

O2A1O1Ixp33_ASAP7_75t_L g3281 ( 
.A1(n_2159),
.A2(n_2222),
.B(n_2188),
.C(n_2622),
.Y(n_3281)
);

INVx3_ASAP7_75t_L g3282 ( 
.A(n_2726),
.Y(n_3282)
);

CKINVDCx10_ASAP7_75t_R g3283 ( 
.A(n_2232),
.Y(n_3283)
);

NAND2xp5_ASAP7_75t_L g3284 ( 
.A(n_2752),
.B(n_2295),
.Y(n_3284)
);

INVx3_ASAP7_75t_L g3285 ( 
.A(n_2726),
.Y(n_3285)
);

AND2x4_ASAP7_75t_L g3286 ( 
.A(n_2168),
.B(n_2239),
.Y(n_3286)
);

AOI21xp5_ASAP7_75t_L g3287 ( 
.A1(n_2511),
.A2(n_2573),
.B(n_2555),
.Y(n_3287)
);

NAND3xp33_ASAP7_75t_L g3288 ( 
.A(n_2773),
.B(n_2771),
.C(n_2622),
.Y(n_3288)
);

OAI22xp5_ASAP7_75t_L g3289 ( 
.A1(n_2717),
.A2(n_2572),
.B1(n_2552),
.B2(n_2684),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_2604),
.B(n_2698),
.Y(n_3290)
);

HB1xp67_ASAP7_75t_L g3291 ( 
.A(n_2809),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_2703),
.A2(n_2658),
.B1(n_2637),
.B2(n_2472),
.Y(n_3292)
);

INVxp67_ASAP7_75t_L g3293 ( 
.A(n_2159),
.Y(n_3293)
);

NOR2xp33_ASAP7_75t_L g3294 ( 
.A(n_2281),
.B(n_2310),
.Y(n_3294)
);

NOR3xp33_ASAP7_75t_L g3295 ( 
.A(n_2302),
.B(n_2749),
.C(n_2744),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2265),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2265),
.Y(n_3297)
);

NOR2x1_ASAP7_75t_L g3298 ( 
.A(n_2648),
.B(n_2393),
.Y(n_3298)
);

INVx3_ASAP7_75t_L g3299 ( 
.A(n_2726),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_2604),
.B(n_2698),
.Y(n_3300)
);

OAI22xp33_ASAP7_75t_L g3301 ( 
.A1(n_2430),
.A2(n_2770),
.B1(n_2695),
.B2(n_2286),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2734),
.B(n_2755),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2511),
.A2(n_2573),
.B(n_2555),
.Y(n_3303)
);

A2O1A1Ixp33_ASAP7_75t_SL g3304 ( 
.A1(n_2234),
.A2(n_2379),
.B(n_2315),
.C(n_2393),
.Y(n_3304)
);

OAI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_2717),
.A2(n_2572),
.B1(n_2552),
.B2(n_2684),
.Y(n_3305)
);

INVx3_ASAP7_75t_L g3306 ( 
.A(n_2726),
.Y(n_3306)
);

NOR2xp33_ASAP7_75t_L g3307 ( 
.A(n_2310),
.B(n_2616),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_2511),
.A2(n_2573),
.B(n_2555),
.Y(n_3308)
);

BUFx2_ASAP7_75t_L g3309 ( 
.A(n_2426),
.Y(n_3309)
);

OAI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_2552),
.A2(n_2572),
.B1(n_2684),
.B2(n_2733),
.Y(n_3310)
);

O2A1O1Ixp33_ASAP7_75t_L g3311 ( 
.A1(n_2803),
.A2(n_2808),
.B(n_2181),
.C(n_2184),
.Y(n_3311)
);

O2A1O1Ixp33_ASAP7_75t_L g3312 ( 
.A1(n_2803),
.A2(n_2808),
.B(n_2181),
.C(n_2184),
.Y(n_3312)
);

BUFx2_ASAP7_75t_L g3313 ( 
.A(n_2426),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2734),
.B(n_2755),
.Y(n_3314)
);

NOR2xp33_ASAP7_75t_L g3315 ( 
.A(n_2616),
.B(n_2532),
.Y(n_3315)
);

INVx3_ASAP7_75t_L g3316 ( 
.A(n_2726),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_2506),
.B(n_2514),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_SL g3318 ( 
.A(n_2511),
.B(n_2555),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_2431),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_2271),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_2555),
.A2(n_2573),
.B(n_2725),
.Y(n_3321)
);

A2O1A1Ixp33_ASAP7_75t_L g3322 ( 
.A1(n_2516),
.A2(n_2509),
.B(n_2488),
.C(n_2733),
.Y(n_3322)
);

OAI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_2506),
.A2(n_2515),
.B1(n_2518),
.B2(n_2514),
.Y(n_3323)
);

BUFx3_ASAP7_75t_L g3324 ( 
.A(n_2251),
.Y(n_3324)
);

A2O1A1Ixp33_ASAP7_75t_L g3325 ( 
.A1(n_2516),
.A2(n_2509),
.B(n_2488),
.C(n_2609),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_2725),
.A2(n_2800),
.B(n_2396),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_SL g3327 ( 
.A(n_2516),
.B(n_2430),
.Y(n_3327)
);

BUFx6f_ASAP7_75t_L g3328 ( 
.A(n_2584),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2506),
.B(n_2514),
.Y(n_3329)
);

BUFx2_ASAP7_75t_L g3330 ( 
.A(n_2426),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2271),
.Y(n_3331)
);

INVx3_ASAP7_75t_L g3332 ( 
.A(n_2729),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_SL g3333 ( 
.A(n_2516),
.B(n_2770),
.Y(n_3333)
);

AOI21xp5_ASAP7_75t_L g3334 ( 
.A1(n_2725),
.A2(n_2800),
.B(n_2396),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_2725),
.A2(n_2800),
.B(n_2396),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_2271),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_2616),
.B(n_2255),
.Y(n_3337)
);

BUFx6f_ASAP7_75t_L g3338 ( 
.A(n_2599),
.Y(n_3338)
);

A2O1A1Ixp33_ASAP7_75t_L g3339 ( 
.A1(n_2488),
.A2(n_2609),
.B(n_2404),
.C(n_2386),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_2515),
.B(n_2518),
.Y(n_3340)
);

O2A1O1Ixp33_ASAP7_75t_SL g3341 ( 
.A1(n_2177),
.A2(n_2475),
.B(n_2565),
.C(n_2560),
.Y(n_3341)
);

AO32x1_ASAP7_75t_L g3342 ( 
.A1(n_2210),
.A2(n_2233),
.A3(n_2164),
.B1(n_2190),
.B2(n_2187),
.Y(n_3342)
);

AOI21x1_ASAP7_75t_L g3343 ( 
.A1(n_2456),
.A2(n_2210),
.B(n_2302),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_2515),
.B(n_2518),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2520),
.B(n_2521),
.Y(n_3345)
);

OA22x2_ASAP7_75t_L g3346 ( 
.A1(n_2602),
.A2(n_2404),
.B1(n_2386),
.B2(n_2574),
.Y(n_3346)
);

O2A1O1Ixp33_ASAP7_75t_L g3347 ( 
.A1(n_2182),
.A2(n_2190),
.B(n_2192),
.C(n_2187),
.Y(n_3347)
);

O2A1O1Ixp33_ASAP7_75t_L g3348 ( 
.A1(n_2182),
.A2(n_2190),
.B(n_2192),
.C(n_2187),
.Y(n_3348)
);

BUFx6f_ASAP7_75t_L g3349 ( 
.A(n_2599),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_2725),
.A2(n_2800),
.B(n_2437),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_SL g3351 ( 
.A(n_2770),
.B(n_2554),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_2520),
.B(n_2521),
.Y(n_3352)
);

OAI22x1_ASAP7_75t_L g3353 ( 
.A1(n_2386),
.A2(n_2404),
.B1(n_2191),
.B2(n_2215),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2276),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_2520),
.B(n_2521),
.Y(n_3355)
);

NOR2xp67_ASAP7_75t_L g3356 ( 
.A(n_2234),
.B(n_2315),
.Y(n_3356)
);

HB1xp67_ASAP7_75t_L g3357 ( 
.A(n_2560),
.Y(n_3357)
);

BUFx6f_ASAP7_75t_L g3358 ( 
.A(n_2599),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_2276),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_2525),
.B(n_2534),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_2800),
.A2(n_2437),
.B(n_2180),
.Y(n_3361)
);

OAI22xp5_ASAP7_75t_L g3362 ( 
.A1(n_2525),
.A2(n_2548),
.B1(n_2550),
.B2(n_2534),
.Y(n_3362)
);

A2O1A1Ixp33_ASAP7_75t_SL g3363 ( 
.A1(n_2234),
.A2(n_2379),
.B(n_2315),
.C(n_2198),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_SL g3364 ( 
.A(n_2554),
.B(n_2730),
.Y(n_3364)
);

NOR2xp33_ASAP7_75t_L g3365 ( 
.A(n_2255),
.B(n_2384),
.Y(n_3365)
);

NAND2x1p5_ASAP7_75t_L g3366 ( 
.A(n_2648),
.B(n_2208),
.Y(n_3366)
);

A2O1A1Ixp33_ASAP7_75t_L g3367 ( 
.A1(n_2574),
.A2(n_2198),
.B(n_2202),
.C(n_2192),
.Y(n_3367)
);

O2A1O1Ixp33_ASAP7_75t_L g3368 ( 
.A1(n_2198),
.A2(n_2491),
.B(n_2492),
.C(n_2202),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_2255),
.B(n_2384),
.Y(n_3369)
);

OAI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_2202),
.A2(n_2492),
.B(n_2491),
.Y(n_3370)
);

OAI22xp5_ASAP7_75t_L g3371 ( 
.A1(n_2525),
.A2(n_2534),
.B1(n_2550),
.B2(n_2548),
.Y(n_3371)
);

AOI21x1_ASAP7_75t_L g3372 ( 
.A1(n_2740),
.A2(n_2492),
.B(n_2491),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_2299),
.B(n_2314),
.Y(n_3373)
);

O2A1O1Ixp33_ASAP7_75t_L g3374 ( 
.A1(n_2744),
.A2(n_2749),
.B(n_2432),
.C(n_2410),
.Y(n_3374)
);

NAND2xp33_ASAP7_75t_L g3375 ( 
.A(n_2795),
.B(n_2479),
.Y(n_3375)
);

NOR3xp33_ASAP7_75t_L g3376 ( 
.A(n_2478),
.B(n_2472),
.C(n_2434),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_2168),
.B(n_2239),
.Y(n_3377)
);

NOR2xp33_ASAP7_75t_L g3378 ( 
.A(n_2384),
.B(n_2677),
.Y(n_3378)
);

O2A1O1Ixp33_ASAP7_75t_L g3379 ( 
.A1(n_2410),
.A2(n_2432),
.B(n_2434),
.C(n_2791),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_2284),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2284),
.Y(n_3381)
);

BUFx8_ASAP7_75t_L g3382 ( 
.A(n_2332),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_2284),
.Y(n_3383)
);

NOR2xp33_ASAP7_75t_L g3384 ( 
.A(n_2677),
.B(n_2692),
.Y(n_3384)
);

CKINVDCx16_ASAP7_75t_R g3385 ( 
.A(n_2332),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_2677),
.B(n_2692),
.Y(n_3386)
);

AOI21xp5_ASAP7_75t_L g3387 ( 
.A1(n_2558),
.A2(n_2656),
.B(n_2644),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_2548),
.B(n_2550),
.Y(n_3388)
);

AOI21xp5_ASAP7_75t_L g3389 ( 
.A1(n_2558),
.A2(n_2656),
.B(n_2644),
.Y(n_3389)
);

OAI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_2543),
.A2(n_2553),
.B(n_2478),
.Y(n_3390)
);

AOI21xp5_ASAP7_75t_L g3391 ( 
.A1(n_2558),
.A2(n_2656),
.B(n_2644),
.Y(n_3391)
);

INVx1_ASAP7_75t_SL g3392 ( 
.A(n_2817),
.Y(n_3392)
);

AND2x2_ASAP7_75t_L g3393 ( 
.A(n_2840),
.B(n_2191),
.Y(n_3393)
);

OAI22xp5_ASAP7_75t_L g3394 ( 
.A1(n_2911),
.A2(n_2574),
.B1(n_2602),
.B2(n_2730),
.Y(n_3394)
);

NAND2xp5_ASAP7_75t_SL g3395 ( 
.A(n_3135),
.B(n_2366),
.Y(n_3395)
);

INVxp67_ASAP7_75t_SL g3396 ( 
.A(n_3250),
.Y(n_3396)
);

OAI21xp5_ASAP7_75t_L g3397 ( 
.A1(n_2967),
.A2(n_2553),
.B(n_2543),
.Y(n_3397)
);

AO31x2_ASAP7_75t_L g3398 ( 
.A1(n_3179),
.A2(n_2191),
.A3(n_2215),
.B(n_2207),
.Y(n_3398)
);

NAND2x1p5_ASAP7_75t_L g3399 ( 
.A(n_2834),
.B(n_2196),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_3153),
.B(n_2212),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3157),
.B(n_2258),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_2917),
.B(n_2918),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2978),
.B(n_2258),
.Y(n_3403)
);

OAI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_3014),
.A2(n_2215),
.B1(n_2248),
.B2(n_2207),
.Y(n_3404)
);

AND2x6_ASAP7_75t_L g3405 ( 
.A(n_2896),
.B(n_2196),
.Y(n_3405)
);

INVx5_ASAP7_75t_L g3406 ( 
.A(n_3242),
.Y(n_3406)
);

AO31x2_ASAP7_75t_L g3407 ( 
.A1(n_3179),
.A2(n_2248),
.A3(n_2253),
.B(n_2207),
.Y(n_3407)
);

NAND3xp33_ASAP7_75t_SL g3408 ( 
.A(n_2978),
.B(n_2874),
.C(n_2872),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_2943),
.B(n_2258),
.Y(n_3409)
);

OAI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_3014),
.A2(n_2253),
.B1(n_2248),
.B2(n_2376),
.Y(n_3410)
);

AO31x2_ASAP7_75t_L g3411 ( 
.A1(n_2985),
.A2(n_3036),
.A3(n_3199),
.B(n_3158),
.Y(n_3411)
);

OAI21xp5_ASAP7_75t_L g3412 ( 
.A1(n_3166),
.A2(n_2553),
.B(n_2543),
.Y(n_3412)
);

INVx4_ASAP7_75t_L g3413 ( 
.A(n_2834),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_SL g3414 ( 
.A(n_3070),
.B(n_2366),
.Y(n_3414)
);

NOR2x1_ASAP7_75t_SL g3415 ( 
.A(n_3042),
.B(n_2196),
.Y(n_3415)
);

AO31x2_ASAP7_75t_L g3416 ( 
.A1(n_2985),
.A2(n_2253),
.A3(n_2237),
.B(n_2240),
.Y(n_3416)
);

OAI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_2964),
.A2(n_2478),
.B(n_2790),
.Y(n_3417)
);

BUFx3_ASAP7_75t_L g3418 ( 
.A(n_3382),
.Y(n_3418)
);

OAI22xp5_ASAP7_75t_L g3419 ( 
.A1(n_3322),
.A2(n_3339),
.B1(n_3325),
.B2(n_2882),
.Y(n_3419)
);

AOI21xp5_ASAP7_75t_L g3420 ( 
.A1(n_2982),
.A2(n_2823),
.B(n_2822),
.Y(n_3420)
);

AOI211x1_ASAP7_75t_L g3421 ( 
.A1(n_2964),
.A2(n_2314),
.B(n_2376),
.C(n_2261),
.Y(n_3421)
);

OA21x2_ASAP7_75t_L g3422 ( 
.A1(n_3203),
.A2(n_2240),
.B(n_2237),
.Y(n_3422)
);

AO31x2_ASAP7_75t_L g3423 ( 
.A1(n_3036),
.A2(n_2237),
.A3(n_2240),
.B(n_2292),
.Y(n_3423)
);

INVx3_ASAP7_75t_L g3424 ( 
.A(n_3236),
.Y(n_3424)
);

AND2x6_ASAP7_75t_L g3425 ( 
.A(n_2896),
.B(n_2196),
.Y(n_3425)
);

NAND2xp5_ASAP7_75t_L g3426 ( 
.A(n_2943),
.B(n_2383),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3258),
.B(n_2383),
.Y(n_3427)
);

BUFx6f_ASAP7_75t_L g3428 ( 
.A(n_2834),
.Y(n_3428)
);

O2A1O1Ixp5_ASAP7_75t_L g3429 ( 
.A1(n_3204),
.A2(n_2234),
.B(n_2379),
.C(n_2315),
.Y(n_3429)
);

OAI21x1_ASAP7_75t_L g3430 ( 
.A1(n_3350),
.A2(n_2693),
.B(n_2537),
.Y(n_3430)
);

OAI21x1_ASAP7_75t_L g3431 ( 
.A1(n_3055),
.A2(n_2693),
.B(n_2537),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3002),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_2836),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_3054),
.Y(n_3434)
);

AOI21xp5_ASAP7_75t_L g3435 ( 
.A1(n_2832),
.A2(n_2562),
.B(n_2519),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_2988),
.A2(n_2562),
.B(n_2519),
.Y(n_3436)
);

OAI21xp5_ASAP7_75t_L g3437 ( 
.A1(n_2882),
.A2(n_2792),
.B(n_2790),
.Y(n_3437)
);

INVx2_ASAP7_75t_SL g3438 ( 
.A(n_2829),
.Y(n_3438)
);

A2O1A1Ixp33_ASAP7_75t_L g3439 ( 
.A1(n_2839),
.A2(n_2376),
.B(n_2314),
.C(n_2168),
.Y(n_3439)
);

HB1xp67_ASAP7_75t_L g3440 ( 
.A(n_3291),
.Y(n_3440)
);

A2O1A1Ixp33_ASAP7_75t_L g3441 ( 
.A1(n_2839),
.A2(n_2376),
.B(n_2168),
.C(n_2247),
.Y(n_3441)
);

AO31x2_ASAP7_75t_L g3442 ( 
.A1(n_3199),
.A2(n_2356),
.A3(n_2373),
.B(n_2292),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_SL g3443 ( 
.A(n_2818),
.B(n_2366),
.Y(n_3443)
);

INVx4_ASAP7_75t_L g3444 ( 
.A(n_2834),
.Y(n_3444)
);

BUFx6f_ASAP7_75t_L g3445 ( 
.A(n_2834),
.Y(n_3445)
);

OAI21x1_ASAP7_75t_L g3446 ( 
.A1(n_3055),
.A2(n_2693),
.B(n_2537),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_L g3447 ( 
.A(n_2833),
.B(n_2286),
.Y(n_3447)
);

NAND2xp33_ASAP7_75t_L g3448 ( 
.A(n_2851),
.B(n_2795),
.Y(n_3448)
);

OAI21x1_ASAP7_75t_SL g3449 ( 
.A1(n_3261),
.A2(n_2266),
.B(n_2235),
.Y(n_3449)
);

OAI22xp5_ASAP7_75t_L g3450 ( 
.A1(n_2989),
.A2(n_2376),
.B1(n_2564),
.B2(n_2557),
.Y(n_3450)
);

OAI21x1_ASAP7_75t_L g3451 ( 
.A1(n_3343),
.A2(n_2387),
.B(n_2760),
.Y(n_3451)
);

OAI21x1_ASAP7_75t_L g3452 ( 
.A1(n_3343),
.A2(n_2387),
.B(n_2760),
.Y(n_3452)
);

OAI21xp5_ASAP7_75t_L g3453 ( 
.A1(n_2894),
.A2(n_2792),
.B(n_2791),
.Y(n_3453)
);

OAI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_2894),
.A2(n_2791),
.B(n_2703),
.Y(n_3454)
);

NAND3xp33_ASAP7_75t_L g3455 ( 
.A(n_2860),
.B(n_2565),
.C(n_2349),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3102),
.B(n_2402),
.Y(n_3456)
);

INVx2_ASAP7_75t_L g3457 ( 
.A(n_3002),
.Y(n_3457)
);

NAND2x1_ASAP7_75t_L g3458 ( 
.A(n_2828),
.B(n_2196),
.Y(n_3458)
);

AO21x2_ASAP7_75t_L g3459 ( 
.A1(n_3363),
.A2(n_2395),
.B(n_2394),
.Y(n_3459)
);

INVx5_ASAP7_75t_L g3460 ( 
.A(n_3242),
.Y(n_3460)
);

NAND3xp33_ASAP7_75t_L g3461 ( 
.A(n_2859),
.B(n_2842),
.C(n_2885),
.Y(n_3461)
);

AOI21x1_ASAP7_75t_SL g3462 ( 
.A1(n_2864),
.A2(n_2779),
.B(n_2772),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3002),
.Y(n_3463)
);

OAI21x1_ASAP7_75t_L g3464 ( 
.A1(n_3361),
.A2(n_2387),
.B(n_2760),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_L g3465 ( 
.A(n_3109),
.B(n_2402),
.Y(n_3465)
);

OAI21xp5_ASAP7_75t_L g3466 ( 
.A1(n_3288),
.A2(n_2703),
.B(n_2768),
.Y(n_3466)
);

AOI21x1_ASAP7_75t_L g3467 ( 
.A1(n_2828),
.A2(n_2782),
.B(n_2774),
.Y(n_3467)
);

OAI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_3288),
.A2(n_2703),
.B(n_2768),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_2836),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2856),
.Y(n_3470)
);

BUFx3_ASAP7_75t_L g3471 ( 
.A(n_3382),
.Y(n_3471)
);

AO32x2_ASAP7_75t_L g3472 ( 
.A1(n_3231),
.A2(n_2471),
.A3(n_2457),
.B1(n_2429),
.B2(n_2504),
.Y(n_3472)
);

OAI21xp5_ASAP7_75t_L g3473 ( 
.A1(n_2907),
.A2(n_2703),
.B(n_2774),
.Y(n_3473)
);

HB1xp67_ASAP7_75t_L g3474 ( 
.A(n_2817),
.Y(n_3474)
);

OAI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_2907),
.A2(n_2845),
.B(n_2879),
.Y(n_3475)
);

AOI21xp5_ASAP7_75t_L g3476 ( 
.A1(n_3063),
.A2(n_2991),
.B(n_2986),
.Y(n_3476)
);

AND3x2_ASAP7_75t_L g3477 ( 
.A(n_3294),
.B(n_2356),
.C(n_2292),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_2889),
.B(n_2338),
.Y(n_3478)
);

INVx3_ASAP7_75t_L g3479 ( 
.A(n_3236),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_2856),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_SL g3481 ( 
.A1(n_3267),
.A2(n_2517),
.B(n_2479),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3128),
.B(n_2403),
.Y(n_3482)
);

AO31x2_ASAP7_75t_L g3483 ( 
.A1(n_3158),
.A2(n_2373),
.A3(n_2356),
.B(n_2754),
.Y(n_3483)
);

A2O1A1Ixp33_ASAP7_75t_L g3484 ( 
.A1(n_3374),
.A2(n_2239),
.B(n_2273),
.C(n_2247),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3337),
.B(n_2403),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_SL g3486 ( 
.A1(n_3247),
.A2(n_2658),
.B(n_2637),
.Y(n_3486)
);

AOI21xp5_ASAP7_75t_L g3487 ( 
.A1(n_2984),
.A2(n_3031),
.B(n_2837),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3251),
.B(n_2557),
.Y(n_3488)
);

NAND2xp5_ASAP7_75t_L g3489 ( 
.A(n_2915),
.B(n_2557),
.Y(n_3489)
);

OAI21xp33_ASAP7_75t_L g3490 ( 
.A1(n_3255),
.A2(n_2746),
.B(n_2566),
.Y(n_3490)
);

INVx2_ASAP7_75t_SL g3491 ( 
.A(n_2829),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_2862),
.Y(n_3492)
);

OAI22xp5_ASAP7_75t_L g3493 ( 
.A1(n_2989),
.A2(n_2566),
.B1(n_2567),
.B2(n_2564),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_2862),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_2840),
.B(n_2426),
.Y(n_3495)
);

AND2x2_ASAP7_75t_L g3496 ( 
.A(n_3233),
.B(n_2426),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_SL g3497 ( 
.A(n_2818),
.B(n_2366),
.Y(n_3497)
);

INVx2_ASAP7_75t_SL g3498 ( 
.A(n_2829),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3233),
.B(n_2426),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_2915),
.B(n_2564),
.Y(n_3500)
);

INVx1_ASAP7_75t_L g3501 ( 
.A(n_2873),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3237),
.B(n_2566),
.Y(n_3502)
);

NAND2xp33_ASAP7_75t_L g3503 ( 
.A(n_3319),
.B(n_3144),
.Y(n_3503)
);

INVx5_ASAP7_75t_L g3504 ( 
.A(n_3242),
.Y(n_3504)
);

NAND2x1p5_ASAP7_75t_L g3505 ( 
.A(n_2834),
.B(n_2196),
.Y(n_3505)
);

AND2x4_ASAP7_75t_L g3506 ( 
.A(n_3242),
.B(n_2239),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3243),
.B(n_2567),
.Y(n_3507)
);

OAI21xp5_ASAP7_75t_L g3508 ( 
.A1(n_2883),
.A2(n_2703),
.B(n_2787),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_2873),
.Y(n_3509)
);

INVx2_ASAP7_75t_L g3510 ( 
.A(n_2852),
.Y(n_3510)
);

AOI21xp5_ASAP7_75t_SL g3511 ( 
.A1(n_3287),
.A2(n_2517),
.B(n_2479),
.Y(n_3511)
);

AOI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_2958),
.A2(n_2705),
.B(n_2656),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_2881),
.Y(n_3513)
);

A2O1A1Ixp33_ASAP7_75t_L g3514 ( 
.A1(n_2893),
.A2(n_2814),
.B(n_3379),
.C(n_3230),
.Y(n_3514)
);

AOI21xp5_ASAP7_75t_L g3515 ( 
.A1(n_2961),
.A2(n_2705),
.B(n_2656),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_2970),
.A2(n_2705),
.B(n_2656),
.Y(n_3516)
);

CKINVDCx11_ASAP7_75t_R g3517 ( 
.A(n_3216),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3244),
.B(n_2426),
.Y(n_3518)
);

OAI21x1_ASAP7_75t_L g3519 ( 
.A1(n_3387),
.A2(n_3391),
.B(n_3389),
.Y(n_3519)
);

INVx2_ASAP7_75t_L g3520 ( 
.A(n_2844),
.Y(n_3520)
);

OAI21xp5_ASAP7_75t_SL g3521 ( 
.A1(n_3247),
.A2(n_2658),
.B(n_2637),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_2844),
.Y(n_3522)
);

OA21x2_ASAP7_75t_L g3523 ( 
.A1(n_3073),
.A2(n_2395),
.B(n_2394),
.Y(n_3523)
);

OAI21xp5_ASAP7_75t_L g3524 ( 
.A1(n_2871),
.A2(n_2787),
.B(n_2746),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3311),
.B(n_3312),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_3295),
.B(n_2567),
.Y(n_3526)
);

OR2x2_ASAP7_75t_L g3527 ( 
.A(n_2827),
.B(n_2617),
.Y(n_3527)
);

OAI21xp5_ASAP7_75t_L g3528 ( 
.A1(n_3024),
.A2(n_2746),
.B(n_2475),
.Y(n_3528)
);

INVx1_ASAP7_75t_SL g3529 ( 
.A(n_2969),
.Y(n_3529)
);

INVx5_ASAP7_75t_L g3530 ( 
.A(n_3242),
.Y(n_3530)
);

OR2x6_ASAP7_75t_L g3531 ( 
.A(n_3259),
.B(n_3246),
.Y(n_3531)
);

OAI21x1_ASAP7_75t_L g3532 ( 
.A1(n_3273),
.A2(n_2176),
.B(n_2162),
.Y(n_3532)
);

AO21x1_ASAP7_75t_L g3533 ( 
.A1(n_3364),
.A2(n_2571),
.B(n_2568),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3370),
.B(n_2910),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_2881),
.Y(n_3535)
);

OAI22x1_ASAP7_75t_L g3536 ( 
.A1(n_3365),
.A2(n_2373),
.B1(n_2235),
.B2(n_2278),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3370),
.B(n_2568),
.Y(n_3537)
);

AO31x2_ASAP7_75t_L g3538 ( 
.A1(n_3261),
.A2(n_2761),
.A3(n_2804),
.B(n_2754),
.Y(n_3538)
);

BUFx2_ASAP7_75t_L g3539 ( 
.A(n_2936),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2910),
.B(n_2568),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3367),
.B(n_2571),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3265),
.B(n_2571),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_L g3543 ( 
.A1(n_2929),
.A2(n_3372),
.B(n_2878),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3154),
.B(n_2578),
.Y(n_3544)
);

AOI21xp5_ASAP7_75t_L g3545 ( 
.A1(n_3234),
.A2(n_2705),
.B(n_2656),
.Y(n_3545)
);

OAI21x1_ASAP7_75t_L g3546 ( 
.A1(n_2929),
.A2(n_3372),
.B(n_3326),
.Y(n_3546)
);

INVxp67_ASAP7_75t_L g3547 ( 
.A(n_3200),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3347),
.B(n_2578),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3348),
.B(n_2578),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3368),
.B(n_2580),
.Y(n_3550)
);

AO31x2_ASAP7_75t_L g3551 ( 
.A1(n_2932),
.A2(n_3222),
.A3(n_3082),
.B(n_3079),
.Y(n_3551)
);

BUFx12f_ASAP7_75t_L g3552 ( 
.A(n_3030),
.Y(n_3552)
);

OAI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3334),
.A2(n_3335),
.B(n_3090),
.Y(n_3553)
);

A2O1A1Ixp33_ASAP7_75t_L g3554 ( 
.A1(n_2893),
.A2(n_2239),
.B(n_2273),
.C(n_2247),
.Y(n_3554)
);

OAI21xp5_ASAP7_75t_L g3555 ( 
.A1(n_3024),
.A2(n_2746),
.B(n_2475),
.Y(n_3555)
);

NAND2x1_ASAP7_75t_L g3556 ( 
.A(n_2901),
.B(n_2196),
.Y(n_3556)
);

AOI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_2942),
.A2(n_2674),
.B(n_2668),
.Y(n_3557)
);

AO22x2_ASAP7_75t_L g3558 ( 
.A1(n_3103),
.A2(n_2327),
.B1(n_2247),
.B2(n_2273),
.Y(n_3558)
);

CKINVDCx5p33_ASAP7_75t_R g3559 ( 
.A(n_3283),
.Y(n_3559)
);

OAI21xp5_ASAP7_75t_L g3560 ( 
.A1(n_3117),
.A2(n_2746),
.B(n_2266),
.Y(n_3560)
);

AND2x2_ASAP7_75t_L g3561 ( 
.A(n_3244),
.B(n_2426),
.Y(n_3561)
);

OAI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_3096),
.A2(n_2746),
.B(n_2266),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3284),
.B(n_2580),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_2942),
.A2(n_2674),
.B(n_2668),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_2887),
.Y(n_3565)
);

BUFx4_ASAP7_75t_SL g3566 ( 
.A(n_3120),
.Y(n_3566)
);

NAND2xp5_ASAP7_75t_L g3567 ( 
.A(n_3071),
.B(n_2580),
.Y(n_3567)
);

OAI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_2816),
.A2(n_2278),
.B(n_2235),
.Y(n_3568)
);

A2O1A1Ixp33_ASAP7_75t_L g3569 ( 
.A1(n_3255),
.A2(n_2273),
.B(n_2247),
.C(n_2637),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3315),
.B(n_2366),
.Y(n_3570)
);

AOI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_2972),
.A2(n_2674),
.B(n_2668),
.Y(n_3571)
);

CKINVDCx20_ASAP7_75t_R g3572 ( 
.A(n_3052),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3302),
.B(n_2582),
.Y(n_3573)
);

AOI21x1_ASAP7_75t_L g3574 ( 
.A1(n_3278),
.A2(n_2782),
.B(n_2487),
.Y(n_3574)
);

INVx4_ASAP7_75t_L g3575 ( 
.A(n_2863),
.Y(n_3575)
);

O2A1O1Ixp5_ASAP7_75t_SL g3576 ( 
.A1(n_3103),
.A2(n_2487),
.B(n_2486),
.C(n_2395),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_L g3577 ( 
.A(n_3314),
.B(n_2582),
.Y(n_3577)
);

OAI22xp5_ASAP7_75t_L g3578 ( 
.A1(n_2819),
.A2(n_2583),
.B1(n_2585),
.B2(n_2582),
.Y(n_3578)
);

OAI21xp5_ASAP7_75t_L g3579 ( 
.A1(n_2816),
.A2(n_2307),
.B(n_2278),
.Y(n_3579)
);

INVx4_ASAP7_75t_L g3580 ( 
.A(n_2863),
.Y(n_3580)
);

NAND3xp33_ASAP7_75t_L g3581 ( 
.A(n_3034),
.B(n_2349),
.C(n_2486),
.Y(n_3581)
);

NOR2x1_ASAP7_75t_R g3582 ( 
.A(n_3150),
.B(n_2332),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_2887),
.Y(n_3583)
);

INVx1_ASAP7_75t_SL g3584 ( 
.A(n_2969),
.Y(n_3584)
);

NOR2xp33_ASAP7_75t_SL g3585 ( 
.A(n_3318),
.B(n_2349),
.Y(n_3585)
);

AND2x2_ASAP7_75t_L g3586 ( 
.A(n_3373),
.B(n_2426),
.Y(n_3586)
);

AOI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3069),
.A2(n_2875),
.B(n_2869),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_2935),
.B(n_2583),
.Y(n_3588)
);

INVx2_ASAP7_75t_SL g3589 ( 
.A(n_2829),
.Y(n_3589)
);

AOI21xp5_ASAP7_75t_L g3590 ( 
.A1(n_3069),
.A2(n_2674),
.B(n_2668),
.Y(n_3590)
);

O2A1O1Ixp5_ASAP7_75t_L g3591 ( 
.A1(n_3023),
.A2(n_2273),
.B(n_2247),
.C(n_2772),
.Y(n_3591)
);

AO21x1_ASAP7_75t_L g3592 ( 
.A1(n_3281),
.A2(n_2585),
.B(n_2583),
.Y(n_3592)
);

AOI21xp5_ASAP7_75t_L g3593 ( 
.A1(n_2876),
.A2(n_2674),
.B(n_2668),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_3321),
.A2(n_2674),
.B(n_2668),
.Y(n_3594)
);

OAI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_2904),
.A2(n_2307),
.B(n_2321),
.Y(n_3595)
);

OAI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_2815),
.A2(n_2307),
.B(n_2321),
.Y(n_3596)
);

INVx3_ASAP7_75t_SL g3597 ( 
.A(n_3319),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3373),
.B(n_2407),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3197),
.A2(n_3115),
.B(n_3249),
.Y(n_3599)
);

NOR3xp33_ASAP7_75t_L g3600 ( 
.A(n_2825),
.B(n_2339),
.C(n_2321),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_2935),
.B(n_2585),
.Y(n_3601)
);

BUFx2_ASAP7_75t_L g3602 ( 
.A(n_2936),
.Y(n_3602)
);

AO31x2_ASAP7_75t_L g3603 ( 
.A1(n_3222),
.A2(n_2761),
.A3(n_2804),
.B(n_2754),
.Y(n_3603)
);

INVx3_ASAP7_75t_L g3604 ( 
.A(n_3236),
.Y(n_3604)
);

OAI21x1_ASAP7_75t_SL g3605 ( 
.A1(n_3235),
.A2(n_3263),
.B(n_3262),
.Y(n_3605)
);

OAI21x1_ASAP7_75t_L g3606 ( 
.A1(n_2950),
.A2(n_2957),
.B(n_2953),
.Y(n_3606)
);

INVx4_ASAP7_75t_L g3607 ( 
.A(n_2863),
.Y(n_3607)
);

A2O1A1Ixp33_ASAP7_75t_L g3608 ( 
.A1(n_3260),
.A2(n_2273),
.B(n_2658),
.C(n_2637),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3171),
.B(n_2587),
.Y(n_3609)
);

AO31x2_ASAP7_75t_L g3610 ( 
.A1(n_3038),
.A2(n_2804),
.A3(n_2761),
.B(n_2285),
.Y(n_3610)
);

AO31x2_ASAP7_75t_L g3611 ( 
.A1(n_3038),
.A2(n_2285),
.A3(n_2287),
.B(n_2284),
.Y(n_3611)
);

AO21x1_ASAP7_75t_L g3612 ( 
.A1(n_3369),
.A2(n_2588),
.B(n_2587),
.Y(n_3612)
);

A2O1A1Ixp33_ASAP7_75t_L g3613 ( 
.A1(n_2919),
.A2(n_2658),
.B(n_2637),
.C(n_2341),
.Y(n_3613)
);

OAI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_2815),
.A2(n_2341),
.B(n_2339),
.Y(n_3614)
);

CKINVDCx5p33_ASAP7_75t_R g3615 ( 
.A(n_3283),
.Y(n_3615)
);

BUFx6f_ASAP7_75t_L g3616 ( 
.A(n_2863),
.Y(n_3616)
);

NOR2xp33_ASAP7_75t_L g3617 ( 
.A(n_2891),
.B(n_2895),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3301),
.B(n_2366),
.Y(n_3618)
);

AOI21xp5_ASAP7_75t_L g3619 ( 
.A1(n_2824),
.A2(n_2710),
.B(n_2705),
.Y(n_3619)
);

AND2x2_ASAP7_75t_L g3620 ( 
.A(n_2827),
.B(n_2407),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3268),
.B(n_2587),
.Y(n_3621)
);

AOI21xp5_ASAP7_75t_L g3622 ( 
.A1(n_2824),
.A2(n_2710),
.B(n_2705),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2909),
.Y(n_3623)
);

AO21x2_ASAP7_75t_L g3624 ( 
.A1(n_3304),
.A2(n_2405),
.B(n_2394),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_L g3625 ( 
.A(n_3310),
.B(n_3317),
.Y(n_3625)
);

A2O1A1Ixp33_ASAP7_75t_L g3626 ( 
.A1(n_2857),
.A2(n_2658),
.B(n_2341),
.C(n_2357),
.Y(n_3626)
);

AOI21xp5_ASAP7_75t_L g3627 ( 
.A1(n_2824),
.A2(n_2710),
.B(n_2705),
.Y(n_3627)
);

AOI21xp5_ASAP7_75t_L g3628 ( 
.A1(n_2824),
.A2(n_2710),
.B(n_2705),
.Y(n_3628)
);

OAI21xp5_ASAP7_75t_L g3629 ( 
.A1(n_2821),
.A2(n_2357),
.B(n_2339),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_2849),
.Y(n_3630)
);

NOR4xp25_ASAP7_75t_L g3631 ( 
.A(n_3058),
.B(n_2590),
.C(n_2591),
.D(n_2588),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_SL g3632 ( 
.A(n_2898),
.B(n_2877),
.Y(n_3632)
);

NAND2x1_ASAP7_75t_L g3633 ( 
.A(n_2901),
.B(n_2196),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3310),
.B(n_2588),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_2921),
.B(n_2407),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_2824),
.A2(n_2710),
.B(n_2591),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3254),
.A2(n_3115),
.B(n_2855),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_3329),
.B(n_2590),
.Y(n_3638)
);

OAI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_2821),
.A2(n_2357),
.B(n_2772),
.Y(n_3639)
);

OA21x2_ASAP7_75t_L g3640 ( 
.A1(n_2841),
.A2(n_2408),
.B(n_2405),
.Y(n_3640)
);

OAI21x1_ASAP7_75t_SL g3641 ( 
.A1(n_3272),
.A2(n_2287),
.B(n_2285),
.Y(n_3641)
);

OAI21x1_ASAP7_75t_L g3642 ( 
.A1(n_2938),
.A2(n_2641),
.B(n_2230),
.Y(n_3642)
);

OA21x2_ASAP7_75t_L g3643 ( 
.A1(n_2841),
.A2(n_2411),
.B(n_2408),
.Y(n_3643)
);

OAI21xp5_ASAP7_75t_L g3644 ( 
.A1(n_2983),
.A2(n_2779),
.B(n_2772),
.Y(n_3644)
);

AOI21xp5_ASAP7_75t_L g3645 ( 
.A1(n_2848),
.A2(n_2710),
.B(n_2591),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3340),
.B(n_2590),
.Y(n_3646)
);

OAI21x1_ASAP7_75t_L g3647 ( 
.A1(n_2941),
.A2(n_2259),
.B(n_2223),
.Y(n_3647)
);

OAI21x1_ASAP7_75t_L g3648 ( 
.A1(n_2948),
.A2(n_2903),
.B(n_2897),
.Y(n_3648)
);

AOI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3197),
.A2(n_2779),
.B(n_2772),
.Y(n_3649)
);

NAND2xp5_ASAP7_75t_SL g3650 ( 
.A(n_2898),
.B(n_3385),
.Y(n_3650)
);

NAND3xp33_ASAP7_75t_SL g3651 ( 
.A(n_3280),
.B(n_2655),
.C(n_2629),
.Y(n_3651)
);

BUFx3_ASAP7_75t_L g3652 ( 
.A(n_3382),
.Y(n_3652)
);

OAI21xp5_ASAP7_75t_L g3653 ( 
.A1(n_3066),
.A2(n_2781),
.B(n_2779),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_3385),
.B(n_2433),
.Y(n_3654)
);

OAI21x1_ASAP7_75t_L g3655 ( 
.A1(n_2906),
.A2(n_2259),
.B(n_2223),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_2974),
.B(n_2338),
.Y(n_3656)
);

AOI21xp5_ASAP7_75t_L g3657 ( 
.A1(n_2848),
.A2(n_2855),
.B(n_3160),
.Y(n_3657)
);

INVx2_ASAP7_75t_SL g3658 ( 
.A(n_2829),
.Y(n_3658)
);

OAI21xp5_ASAP7_75t_L g3659 ( 
.A1(n_3165),
.A2(n_2781),
.B(n_2779),
.Y(n_3659)
);

CKINVDCx5p33_ASAP7_75t_R g3660 ( 
.A(n_3150),
.Y(n_3660)
);

OAI21xp5_ASAP7_75t_L g3661 ( 
.A1(n_2962),
.A2(n_2781),
.B(n_2597),
.Y(n_3661)
);

BUFx6f_ASAP7_75t_L g3662 ( 
.A(n_2863),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_2909),
.Y(n_3663)
);

OAI21x1_ASAP7_75t_SL g3664 ( 
.A1(n_3275),
.A2(n_2287),
.B(n_2285),
.Y(n_3664)
);

NOR2x1_ASAP7_75t_L g3665 ( 
.A(n_3298),
.B(n_2675),
.Y(n_3665)
);

OAI21xp5_ASAP7_75t_L g3666 ( 
.A1(n_3298),
.A2(n_2781),
.B(n_2597),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3344),
.B(n_2596),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3345),
.B(n_2596),
.Y(n_3668)
);

NAND2x1_ASAP7_75t_L g3669 ( 
.A(n_2901),
.B(n_2196),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_2846),
.B(n_2433),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_3236),
.B(n_2200),
.Y(n_3671)
);

BUFx2_ASAP7_75t_R g3672 ( 
.A(n_3202),
.Y(n_3672)
);

BUFx12f_ASAP7_75t_L g3673 ( 
.A(n_2912),
.Y(n_3673)
);

NAND3xp33_ASAP7_75t_L g3674 ( 
.A(n_2892),
.B(n_3122),
.C(n_3095),
.Y(n_3674)
);

OAI22xp5_ASAP7_75t_L g3675 ( 
.A1(n_2819),
.A2(n_2597),
.B1(n_2610),
.B2(n_2596),
.Y(n_3675)
);

OAI21xp5_ASAP7_75t_L g3676 ( 
.A1(n_3050),
.A2(n_2781),
.B(n_2612),
.Y(n_3676)
);

OAI22x1_ASAP7_75t_L g3677 ( 
.A1(n_3269),
.A2(n_2457),
.B1(n_2471),
.B2(n_2429),
.Y(n_3677)
);

CKINVDCx5p33_ASAP7_75t_R g3678 ( 
.A(n_2912),
.Y(n_3678)
);

OA21x2_ASAP7_75t_L g3679 ( 
.A1(n_3067),
.A2(n_2412),
.B(n_2411),
.Y(n_3679)
);

NOR2x1_ASAP7_75t_L g3680 ( 
.A(n_3116),
.B(n_2675),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_2998),
.B(n_3245),
.Y(n_3681)
);

BUFx8_ASAP7_75t_L g3682 ( 
.A(n_2965),
.Y(n_3682)
);

OAI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3167),
.A2(n_2781),
.B(n_2612),
.Y(n_3683)
);

NAND2xp5_ASAP7_75t_L g3684 ( 
.A(n_3352),
.B(n_2610),
.Y(n_3684)
);

INVx2_ASAP7_75t_SL g3685 ( 
.A(n_2913),
.Y(n_3685)
);

BUFx3_ASAP7_75t_L g3686 ( 
.A(n_3382),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_2849),
.Y(n_3687)
);

OAI22xp5_ASAP7_75t_L g3688 ( 
.A1(n_3346),
.A2(n_2612),
.B1(n_2614),
.B2(n_2610),
.Y(n_3688)
);

BUFx10_ASAP7_75t_L g3689 ( 
.A(n_3208),
.Y(n_3689)
);

OAI21x1_ASAP7_75t_L g3690 ( 
.A1(n_2963),
.A2(n_3074),
.B(n_2843),
.Y(n_3690)
);

INVx4_ASAP7_75t_L g3691 ( 
.A(n_2863),
.Y(n_3691)
);

NOR2x1_ASAP7_75t_L g3692 ( 
.A(n_3184),
.B(n_2675),
.Y(n_3692)
);

NOR2xp33_ASAP7_75t_L g3693 ( 
.A(n_3307),
.B(n_2677),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3355),
.B(n_2614),
.Y(n_3694)
);

OAI22xp5_ASAP7_75t_L g3695 ( 
.A1(n_3346),
.A2(n_3269),
.B1(n_2867),
.B2(n_2838),
.Y(n_3695)
);

AO32x2_ASAP7_75t_L g3696 ( 
.A1(n_3231),
.A2(n_2504),
.A3(n_2570),
.B1(n_2801),
.B2(n_2617),
.Y(n_3696)
);

AOI22xp5_ASAP7_75t_L g3697 ( 
.A1(n_3351),
.A2(n_2695),
.B1(n_2493),
.B2(n_2655),
.Y(n_3697)
);

OAI21x1_ASAP7_75t_L g3698 ( 
.A1(n_3091),
.A2(n_2378),
.B(n_2325),
.Y(n_3698)
);

NOR2xp67_ASAP7_75t_SL g3699 ( 
.A(n_2965),
.B(n_2332),
.Y(n_3699)
);

BUFx6f_ASAP7_75t_L g3700 ( 
.A(n_3123),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_2921),
.B(n_2407),
.Y(n_3701)
);

A2O1A1Ixp33_ASAP7_75t_L g3702 ( 
.A1(n_2838),
.A2(n_2204),
.B(n_2225),
.C(n_2200),
.Y(n_3702)
);

CKINVDCx5p33_ASAP7_75t_R g3703 ( 
.A(n_3256),
.Y(n_3703)
);

AND2x2_ASAP7_75t_SL g3704 ( 
.A(n_3004),
.B(n_2200),
.Y(n_3704)
);

INVx1_ASAP7_75t_SL g3705 ( 
.A(n_2928),
.Y(n_3705)
);

AO31x2_ASAP7_75t_L g3706 ( 
.A1(n_3078),
.A2(n_2293),
.A3(n_2300),
.B(n_2287),
.Y(n_3706)
);

NOR2xp33_ASAP7_75t_L g3707 ( 
.A(n_2886),
.B(n_2677),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3360),
.B(n_2614),
.Y(n_3708)
);

AND2x4_ASAP7_75t_L g3709 ( 
.A(n_3286),
.B(n_3377),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_2849),
.Y(n_3710)
);

INVxp67_ASAP7_75t_SL g3711 ( 
.A(n_3357),
.Y(n_3711)
);

O2A1O1Ixp5_ASAP7_75t_L g3712 ( 
.A1(n_2899),
.A2(n_2784),
.B(n_2765),
.C(n_2442),
.Y(n_3712)
);

OR2x6_ASAP7_75t_L g3713 ( 
.A(n_2826),
.B(n_2200),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_2922),
.Y(n_3714)
);

OAI21xp33_ASAP7_75t_L g3715 ( 
.A1(n_3346),
.A2(n_2625),
.B(n_2624),
.Y(n_3715)
);

AOI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3088),
.A2(n_2625),
.B(n_2624),
.Y(n_3716)
);

AOI21xp33_ASAP7_75t_L g3717 ( 
.A1(n_3167),
.A2(n_2625),
.B(n_2624),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_2922),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_L g3719 ( 
.A(n_3388),
.B(n_2626),
.Y(n_3719)
);

A2O1A1Ixp33_ASAP7_75t_L g3720 ( 
.A1(n_3252),
.A2(n_2204),
.B(n_2225),
.C(n_2200),
.Y(n_3720)
);

AO21x2_ASAP7_75t_L g3721 ( 
.A1(n_3112),
.A2(n_2412),
.B(n_2411),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_2852),
.Y(n_3722)
);

BUFx3_ASAP7_75t_L g3723 ( 
.A(n_2853),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_3192),
.B(n_2626),
.Y(n_3724)
);

OAI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_3092),
.A2(n_2651),
.B(n_2626),
.Y(n_3725)
);

INVx3_ASAP7_75t_SL g3726 ( 
.A(n_3238),
.Y(n_3726)
);

AOI211x1_ASAP7_75t_L g3727 ( 
.A1(n_2861),
.A2(n_2261),
.B(n_2263),
.C(n_2256),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_2928),
.B(n_2617),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3375),
.A2(n_2652),
.B(n_2651),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3223),
.B(n_2651),
.Y(n_3730)
);

AOI21xp33_ASAP7_75t_L g3731 ( 
.A1(n_2830),
.A2(n_2664),
.B(n_2652),
.Y(n_3731)
);

OAI21x1_ASAP7_75t_L g3732 ( 
.A1(n_3037),
.A2(n_3155),
.B(n_2971),
.Y(n_3732)
);

BUFx6f_ASAP7_75t_L g3733 ( 
.A(n_3123),
.Y(n_3733)
);

OAI21x1_ASAP7_75t_L g3734 ( 
.A1(n_3037),
.A2(n_2462),
.B(n_2443),
.Y(n_3734)
);

OAI21x1_ASAP7_75t_L g3735 ( 
.A1(n_3155),
.A2(n_2971),
.B(n_3187),
.Y(n_3735)
);

NAND2xp33_ASAP7_75t_SL g3736 ( 
.A(n_3238),
.B(n_2517),
.Y(n_3736)
);

AO31x2_ASAP7_75t_L g3737 ( 
.A1(n_3078),
.A2(n_2300),
.A3(n_2306),
.B(n_2293),
.Y(n_3737)
);

AOI221xp5_ASAP7_75t_L g3738 ( 
.A1(n_3289),
.A2(n_2652),
.B1(n_2664),
.B2(n_2665),
.C(n_2667),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_2852),
.Y(n_3739)
);

BUFx3_ASAP7_75t_L g3740 ( 
.A(n_2853),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3290),
.B(n_2664),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_3300),
.B(n_2665),
.Y(n_3742)
);

AOI21xp5_ASAP7_75t_SL g3743 ( 
.A1(n_3303),
.A2(n_3308),
.B(n_3000),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3323),
.B(n_2665),
.Y(n_3744)
);

NOR2x1_ASAP7_75t_L g3745 ( 
.A(n_3323),
.B(n_2675),
.Y(n_3745)
);

OAI21x1_ASAP7_75t_L g3746 ( 
.A1(n_3188),
.A2(n_2462),
.B(n_2443),
.Y(n_3746)
);

AND2x2_ASAP7_75t_L g3747 ( 
.A(n_2939),
.B(n_2465),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_2939),
.B(n_2465),
.Y(n_3748)
);

OAI21x1_ASAP7_75t_L g3749 ( 
.A1(n_3189),
.A2(n_2502),
.B(n_2462),
.Y(n_3749)
);

OAI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_2880),
.A2(n_2671),
.B(n_2667),
.Y(n_3750)
);

OAI21x1_ASAP7_75t_L g3751 ( 
.A1(n_3193),
.A2(n_2523),
.B(n_2502),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_2848),
.A2(n_2710),
.B(n_2671),
.Y(n_3752)
);

NAND2xp5_ASAP7_75t_L g3753 ( 
.A(n_3362),
.B(n_2667),
.Y(n_3753)
);

AOI21x1_ASAP7_75t_L g3754 ( 
.A1(n_3084),
.A2(n_2415),
.B(n_2412),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_2848),
.A2(n_2710),
.B(n_2671),
.Y(n_3755)
);

A2O1A1Ixp33_ASAP7_75t_L g3756 ( 
.A1(n_3266),
.A2(n_2204),
.B(n_2225),
.C(n_2200),
.Y(n_3756)
);

OAI21x1_ASAP7_75t_L g3757 ( 
.A1(n_3201),
.A2(n_3215),
.B(n_3210),
.Y(n_3757)
);

AO32x2_ASAP7_75t_L g3758 ( 
.A1(n_3239),
.A2(n_2570),
.A3(n_2801),
.B1(n_2301),
.B2(n_2208),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_SL g3759 ( 
.A(n_2820),
.B(n_2433),
.Y(n_3759)
);

OAI22x1_ASAP7_75t_L g3760 ( 
.A1(n_3240),
.A2(n_3248),
.B1(n_2890),
.B2(n_2959),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3362),
.B(n_2452),
.Y(n_3761)
);

AOI21xp5_ASAP7_75t_L g3762 ( 
.A1(n_2848),
.A2(n_2710),
.B(n_2784),
.Y(n_3762)
);

BUFx2_ASAP7_75t_L g3763 ( 
.A(n_2936),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_L g3764 ( 
.A(n_3371),
.B(n_2452),
.Y(n_3764)
);

INVx1_ASAP7_75t_SL g3765 ( 
.A(n_2981),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_2855),
.A2(n_2784),
.B(n_2683),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_2855),
.A2(n_2784),
.B(n_2683),
.Y(n_3767)
);

OAI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_2979),
.A2(n_2683),
.B(n_2682),
.Y(n_3768)
);

OAI21x1_ASAP7_75t_L g3769 ( 
.A1(n_3219),
.A2(n_2523),
.B(n_2502),
.Y(n_3769)
);

AOI22xp5_ASAP7_75t_L g3770 ( 
.A1(n_2835),
.A2(n_2695),
.B1(n_2493),
.B2(n_2688),
.Y(n_3770)
);

INVx3_ASAP7_75t_SL g3771 ( 
.A(n_3238),
.Y(n_3771)
);

BUFx4_ASAP7_75t_SL g3772 ( 
.A(n_2896),
.Y(n_3772)
);

AOI21x1_ASAP7_75t_L g3773 ( 
.A1(n_3084),
.A2(n_2421),
.B(n_2415),
.Y(n_3773)
);

AO31x2_ASAP7_75t_L g3774 ( 
.A1(n_3152),
.A2(n_2300),
.A3(n_2306),
.B(n_2293),
.Y(n_3774)
);

HB1xp67_ASAP7_75t_L g3775 ( 
.A(n_2914),
.Y(n_3775)
);

INVx1_ASAP7_75t_L g3776 ( 
.A(n_2947),
.Y(n_3776)
);

AOI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_2847),
.A2(n_2695),
.B1(n_2688),
.B2(n_2629),
.Y(n_3777)
);

NAND2xp5_ASAP7_75t_L g3778 ( 
.A(n_3371),
.B(n_2682),
.Y(n_3778)
);

OAI21xp5_ASAP7_75t_L g3779 ( 
.A1(n_3105),
.A2(n_2687),
.B(n_2682),
.Y(n_3779)
);

AOI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_2855),
.A2(n_2784),
.B(n_2689),
.Y(n_3780)
);

OAI22x1_ASAP7_75t_L g3781 ( 
.A1(n_2992),
.A2(n_2256),
.B1(n_2263),
.B2(n_2261),
.Y(n_3781)
);

AO31x2_ASAP7_75t_L g3782 ( 
.A1(n_3152),
.A2(n_2300),
.A3(n_2306),
.B(n_2293),
.Y(n_3782)
);

AOI21xp5_ASAP7_75t_L g3783 ( 
.A1(n_3015),
.A2(n_2784),
.B(n_2689),
.Y(n_3783)
);

NOR2xp33_ASAP7_75t_L g3784 ( 
.A(n_2916),
.B(n_2677),
.Y(n_3784)
);

AND2x2_ASAP7_75t_L g3785 ( 
.A(n_2981),
.B(n_2465),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_2865),
.Y(n_3786)
);

AO31x2_ASAP7_75t_L g3787 ( 
.A1(n_3239),
.A2(n_2309),
.A3(n_2319),
.B(n_2306),
.Y(n_3787)
);

NAND2x1_ASAP7_75t_L g3788 ( 
.A(n_2901),
.B(n_2200),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_2947),
.Y(n_3789)
);

OAI21xp5_ASAP7_75t_L g3790 ( 
.A1(n_3022),
.A2(n_2689),
.B(n_2687),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3011),
.B(n_2687),
.Y(n_3791)
);

AOI21xp5_ASAP7_75t_L g3792 ( 
.A1(n_3169),
.A2(n_2700),
.B(n_2694),
.Y(n_3792)
);

NOR4xp25_ASAP7_75t_L g3793 ( 
.A(n_3061),
.B(n_2700),
.C(n_2701),
.D(n_2694),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_SL g3794 ( 
.A(n_3044),
.B(n_2433),
.Y(n_3794)
);

INVx4_ASAP7_75t_L g3795 ( 
.A(n_3191),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3044),
.B(n_2433),
.Y(n_3796)
);

INVx2_ASAP7_75t_L g3797 ( 
.A(n_2865),
.Y(n_3797)
);

NAND2xp5_ASAP7_75t_L g3798 ( 
.A(n_3051),
.B(n_2694),
.Y(n_3798)
);

OAI21x1_ASAP7_75t_L g3799 ( 
.A1(n_3227),
.A2(n_2579),
.B(n_2544),
.Y(n_3799)
);

NOR2xp33_ASAP7_75t_L g3800 ( 
.A(n_2934),
.B(n_2692),
.Y(n_3800)
);

AND2x4_ASAP7_75t_L g3801 ( 
.A(n_3286),
.B(n_2200),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_2952),
.Y(n_3802)
);

AOI21xp5_ASAP7_75t_L g3803 ( 
.A1(n_3170),
.A2(n_2701),
.B(n_2700),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3110),
.B(n_3274),
.Y(n_3804)
);

AND2x2_ASAP7_75t_L g3805 ( 
.A(n_2990),
.B(n_2465),
.Y(n_3805)
);

AO31x2_ASAP7_75t_L g3806 ( 
.A1(n_3087),
.A2(n_2370),
.A3(n_2367),
.B(n_2363),
.Y(n_3806)
);

AOI21xp5_ASAP7_75t_L g3807 ( 
.A1(n_3318),
.A2(n_2728),
.B(n_2701),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_SL g3808 ( 
.A(n_3044),
.B(n_2433),
.Y(n_3808)
);

AND2x2_ASAP7_75t_L g3809 ( 
.A(n_2990),
.B(n_2391),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_2826),
.A2(n_3004),
.B(n_3000),
.Y(n_3810)
);

NAND3x1_ASAP7_75t_L g3811 ( 
.A(n_3376),
.B(n_2263),
.C(n_2256),
.Y(n_3811)
);

A2O1A1Ixp33_ASAP7_75t_L g3812 ( 
.A1(n_3004),
.A2(n_2372),
.B(n_2316),
.C(n_2340),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_L g3813 ( 
.A(n_3137),
.B(n_2728),
.Y(n_3813)
);

OAI21x1_ASAP7_75t_L g3814 ( 
.A1(n_3012),
.A2(n_2579),
.B(n_2544),
.Y(n_3814)
);

AO31x2_ASAP7_75t_L g3815 ( 
.A1(n_3087),
.A2(n_2865),
.A3(n_2994),
.B(n_2925),
.Y(n_3815)
);

A2O1A1Ixp33_ASAP7_75t_L g3816 ( 
.A1(n_3270),
.A2(n_2372),
.B(n_2316),
.C(n_2340),
.Y(n_3816)
);

OAI21xp5_ASAP7_75t_SL g3817 ( 
.A1(n_3327),
.A2(n_2482),
.B(n_2454),
.Y(n_3817)
);

OA22x2_ASAP7_75t_L g3818 ( 
.A1(n_3056),
.A2(n_2391),
.B1(n_2765),
.B2(n_2324),
.Y(n_3818)
);

OAI21xp5_ASAP7_75t_L g3819 ( 
.A1(n_3214),
.A2(n_3043),
.B(n_3010),
.Y(n_3819)
);

OAI21x1_ASAP7_75t_L g3820 ( 
.A1(n_3012),
.A2(n_3366),
.B(n_3149),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_3138),
.B(n_2728),
.Y(n_3821)
);

OR2x2_ASAP7_75t_L g3822 ( 
.A(n_2993),
.B(n_2391),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3293),
.B(n_2741),
.Y(n_3823)
);

O2A1O1Ixp33_ASAP7_75t_L g3824 ( 
.A1(n_2905),
.A2(n_2757),
.B(n_2747),
.C(n_2742),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_2826),
.A2(n_2742),
.B(n_2741),
.Y(n_3825)
);

OAI21xp5_ASAP7_75t_L g3826 ( 
.A1(n_3043),
.A2(n_2742),
.B(n_2741),
.Y(n_3826)
);

INVx1_ASAP7_75t_L g3827 ( 
.A(n_2952),
.Y(n_3827)
);

OAI21x1_ASAP7_75t_SL g3828 ( 
.A1(n_3067),
.A2(n_2319),
.B(n_2309),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_2940),
.B(n_2747),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_2940),
.B(n_2747),
.Y(n_3830)
);

OAI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_3027),
.A2(n_2757),
.B(n_2801),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_2925),
.Y(n_3832)
);

HB1xp67_ASAP7_75t_L g3833 ( 
.A(n_3147),
.Y(n_3833)
);

AOI21xp5_ASAP7_75t_L g3834 ( 
.A1(n_2826),
.A2(n_2757),
.B(n_2789),
.Y(n_3834)
);

AND2x2_ASAP7_75t_L g3835 ( 
.A(n_2993),
.B(n_2391),
.Y(n_3835)
);

OA21x2_ASAP7_75t_L g3836 ( 
.A1(n_3390),
.A2(n_2421),
.B(n_2415),
.Y(n_3836)
);

OAI21x1_ASAP7_75t_L g3837 ( 
.A1(n_3366),
.A2(n_2579),
.B(n_2544),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3045),
.B(n_2454),
.Y(n_3838)
);

NOR2xp33_ASAP7_75t_L g3839 ( 
.A(n_2946),
.B(n_2692),
.Y(n_3839)
);

NAND2xp5_ASAP7_75t_L g3840 ( 
.A(n_2954),
.B(n_2309),
.Y(n_3840)
);

CKINVDCx11_ASAP7_75t_R g3841 ( 
.A(n_3202),
.Y(n_3841)
);

AOI21x1_ASAP7_75t_L g3842 ( 
.A1(n_3057),
.A2(n_2422),
.B(n_2421),
.Y(n_3842)
);

AOI21xp5_ASAP7_75t_L g3843 ( 
.A1(n_2826),
.A2(n_2798),
.B(n_2789),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3286),
.B(n_2204),
.Y(n_3844)
);

OAI21x1_ASAP7_75t_L g3845 ( 
.A1(n_3366),
.A2(n_2657),
.B(n_2579),
.Y(n_3845)
);

O2A1O1Ixp5_ASAP7_75t_L g3846 ( 
.A1(n_3072),
.A2(n_2765),
.B(n_2669),
.C(n_2679),
.Y(n_3846)
);

BUFx2_ASAP7_75t_SL g3847 ( 
.A(n_3181),
.Y(n_3847)
);

AOI21xp5_ASAP7_75t_L g3848 ( 
.A1(n_2966),
.A2(n_2798),
.B(n_2789),
.Y(n_3848)
);

NAND2x1p5_ASAP7_75t_L g3849 ( 
.A(n_2850),
.B(n_2204),
.Y(n_3849)
);

OAI21x1_ASAP7_75t_L g3850 ( 
.A1(n_3149),
.A2(n_3100),
.B(n_3007),
.Y(n_3850)
);

OAI21xp5_ASAP7_75t_L g3851 ( 
.A1(n_2973),
.A2(n_2764),
.B(n_2762),
.Y(n_3851)
);

INVx8_ASAP7_75t_L g3852 ( 
.A(n_2901),
.Y(n_3852)
);

OAI22xp5_ASAP7_75t_SL g3853 ( 
.A1(n_3353),
.A2(n_3183),
.B1(n_3305),
.B2(n_3289),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_2994),
.Y(n_3854)
);

INVx3_ASAP7_75t_L g3855 ( 
.A(n_3286),
.Y(n_3855)
);

OAI21xp33_ASAP7_75t_L g3856 ( 
.A1(n_2870),
.A2(n_2680),
.B(n_2673),
.Y(n_3856)
);

OAI22x1_ASAP7_75t_L g3857 ( 
.A1(n_3333),
.A2(n_2324),
.B1(n_2381),
.B2(n_2377),
.Y(n_3857)
);

AO21x2_ASAP7_75t_L g3858 ( 
.A1(n_3113),
.A2(n_2423),
.B(n_2422),
.Y(n_3858)
);

OAI21x1_ASAP7_75t_L g3859 ( 
.A1(n_3007),
.A2(n_2669),
.B(n_2657),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_2954),
.B(n_2309),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3003),
.B(n_2391),
.Y(n_3861)
);

NAND3xp33_ASAP7_75t_SL g3862 ( 
.A(n_2868),
.B(n_2269),
.C(n_2264),
.Y(n_3862)
);

NOR4xp25_ASAP7_75t_L g3863 ( 
.A(n_3151),
.B(n_2371),
.C(n_2374),
.D(n_2377),
.Y(n_3863)
);

AO221x2_ASAP7_75t_L g3864 ( 
.A1(n_3353),
.A2(n_2327),
.B1(n_2324),
.B2(n_2353),
.C(n_2371),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_2931),
.B(n_2319),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_2944),
.B(n_2692),
.Y(n_3866)
);

OAI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_3209),
.A2(n_2764),
.B(n_2762),
.Y(n_3867)
);

OAI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3209),
.A2(n_2785),
.B(n_2765),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3006),
.Y(n_3869)
);

NOR2xp33_ASAP7_75t_L g3870 ( 
.A(n_2884),
.B(n_2692),
.Y(n_3870)
);

OR2x2_ASAP7_75t_L g3871 ( 
.A(n_3003),
.B(n_2391),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3006),
.Y(n_3872)
);

INVx1_ASAP7_75t_L g3873 ( 
.A(n_2956),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3097),
.B(n_2391),
.Y(n_3874)
);

INVx5_ASAP7_75t_L g3875 ( 
.A(n_3041),
.Y(n_3875)
);

NAND2xp5_ASAP7_75t_L g3876 ( 
.A(n_2968),
.B(n_2319),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_L g3877 ( 
.A(n_2980),
.B(n_2348),
.Y(n_3877)
);

OAI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_3159),
.A2(n_2924),
.B(n_2933),
.Y(n_3878)
);

AO221x2_ASAP7_75t_L g3879 ( 
.A1(n_3151),
.A2(n_2327),
.B1(n_2371),
.B2(n_2374),
.C(n_2392),
.Y(n_3879)
);

NAND2x1p5_ASAP7_75t_L g3880 ( 
.A(n_2850),
.B(n_2204),
.Y(n_3880)
);

NOR2xp33_ASAP7_75t_L g3881 ( 
.A(n_2937),
.B(n_2454),
.Y(n_3881)
);

OAI22xp5_ASAP7_75t_L g3882 ( 
.A1(n_3056),
.A2(n_2161),
.B1(n_2185),
.B2(n_2195),
.Y(n_3882)
);

NAND2x1p5_ASAP7_75t_L g3883 ( 
.A(n_2850),
.B(n_2204),
.Y(n_3883)
);

NOR2xp67_ASAP7_75t_L g3884 ( 
.A(n_3356),
.B(n_2204),
.Y(n_3884)
);

AOI221xp5_ASAP7_75t_L g3885 ( 
.A1(n_3305),
.A2(n_2680),
.B1(n_2673),
.B2(n_2785),
.C(n_2374),
.Y(n_3885)
);

OAI21x1_ASAP7_75t_L g3886 ( 
.A1(n_2908),
.A2(n_2713),
.B(n_2679),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3177),
.A2(n_2798),
.B(n_2789),
.Y(n_3887)
);

OA21x2_ASAP7_75t_L g3888 ( 
.A1(n_3390),
.A2(n_2423),
.B(n_2422),
.Y(n_3888)
);

AOI21xp5_ASAP7_75t_L g3889 ( 
.A1(n_2996),
.A2(n_3225),
.B(n_3217),
.Y(n_3889)
);

OAI21xp5_ASAP7_75t_L g3890 ( 
.A1(n_2924),
.A2(n_2765),
.B(n_2753),
.Y(n_3890)
);

OAI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_2995),
.A2(n_3146),
.B(n_2996),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3020),
.Y(n_3892)
);

OAI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_2854),
.A2(n_2765),
.B(n_2753),
.Y(n_3893)
);

AND2x2_ASAP7_75t_L g3894 ( 
.A(n_3097),
.B(n_2805),
.Y(n_3894)
);

A2O1A1Ixp33_ASAP7_75t_L g3895 ( 
.A1(n_3045),
.A2(n_2372),
.B(n_2340),
.C(n_2316),
.Y(n_3895)
);

BUFx2_ASAP7_75t_L g3896 ( 
.A(n_2936),
.Y(n_3896)
);

A2O1A1Ixp33_ASAP7_75t_L g3897 ( 
.A1(n_3045),
.A2(n_2372),
.B(n_2340),
.C(n_2316),
.Y(n_3897)
);

NAND2x1p5_ASAP7_75t_L g3898 ( 
.A(n_3005),
.B(n_2204),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_2987),
.A2(n_2798),
.B(n_2789),
.Y(n_3899)
);

OAI21x1_ASAP7_75t_L g3900 ( 
.A1(n_2975),
.A2(n_2713),
.B(n_2679),
.Y(n_3900)
);

AOI221x1_ASAP7_75t_L g3901 ( 
.A1(n_3253),
.A2(n_2425),
.B1(n_2461),
.B2(n_2455),
.C(n_2470),
.Y(n_3901)
);

OAI21x1_ASAP7_75t_L g3902 ( 
.A1(n_2975),
.A2(n_2713),
.B(n_2679),
.Y(n_3902)
);

OAI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_3271),
.A2(n_2161),
.B1(n_2185),
.B2(n_2195),
.Y(n_3903)
);

AOI221xp5_ASAP7_75t_L g3904 ( 
.A1(n_3253),
.A2(n_2680),
.B1(n_2673),
.B2(n_2353),
.C(n_2352),
.Y(n_3904)
);

OAI21x1_ASAP7_75t_L g3905 ( 
.A1(n_2975),
.A2(n_2713),
.B(n_2467),
.Y(n_3905)
);

NOR2xp67_ASAP7_75t_L g3906 ( 
.A(n_3356),
.B(n_2225),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2999),
.B(n_2348),
.Y(n_3907)
);

INVx3_ASAP7_75t_L g3908 ( 
.A(n_3377),
.Y(n_3908)
);

INVx1_ASAP7_75t_L g3909 ( 
.A(n_2956),
.Y(n_3909)
);

BUFx2_ASAP7_75t_L g3910 ( 
.A(n_2936),
.Y(n_3910)
);

AOI21xp5_ASAP7_75t_L g3911 ( 
.A1(n_2987),
.A2(n_2798),
.B(n_2789),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_2976),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_3342),
.A2(n_2798),
.B(n_2635),
.Y(n_3913)
);

OAI21x1_ASAP7_75t_L g3914 ( 
.A1(n_3094),
.A2(n_2467),
.B(n_2458),
.Y(n_3914)
);

BUFx2_ASAP7_75t_L g3915 ( 
.A(n_3309),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3013),
.B(n_2385),
.Y(n_3916)
);

OAI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_2888),
.A2(n_2753),
.B(n_2635),
.Y(n_3917)
);

OR2x2_ASAP7_75t_L g3918 ( 
.A(n_3309),
.B(n_2225),
.Y(n_3918)
);

NOR2xp33_ASAP7_75t_L g3919 ( 
.A(n_2900),
.B(n_2454),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_SL g3920 ( 
.A(n_3124),
.B(n_2454),
.Y(n_3920)
);

OAI21x1_ASAP7_75t_L g3921 ( 
.A1(n_3094),
.A2(n_2458),
.B(n_2425),
.Y(n_3921)
);

AND2x2_ASAP7_75t_L g3922 ( 
.A(n_3313),
.B(n_2805),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_2976),
.Y(n_3923)
);

INVx5_ASAP7_75t_L g3924 ( 
.A(n_3041),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_2977),
.Y(n_3925)
);

OA22x2_ASAP7_75t_L g3926 ( 
.A1(n_3098),
.A2(n_2377),
.B1(n_2344),
.B2(n_2352),
.Y(n_3926)
);

AND2x4_ASAP7_75t_L g3927 ( 
.A(n_3377),
.B(n_2225),
.Y(n_3927)
);

NAND2xp5_ASAP7_75t_SL g3928 ( 
.A(n_3124),
.B(n_2454),
.Y(n_3928)
);

INVx2_ASAP7_75t_L g3929 ( 
.A(n_3076),
.Y(n_3929)
);

OA22x2_ASAP7_75t_L g3930 ( 
.A1(n_3098),
.A2(n_2304),
.B1(n_2392),
.B2(n_2353),
.Y(n_3930)
);

INVx3_ASAP7_75t_L g3931 ( 
.A(n_3377),
.Y(n_3931)
);

AOI21xp5_ASAP7_75t_L g3932 ( 
.A1(n_3342),
.A2(n_3207),
.B(n_2691),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_2977),
.Y(n_3933)
);

OAI21x1_ASAP7_75t_L g3934 ( 
.A1(n_3094),
.A2(n_2436),
.B(n_2428),
.Y(n_3934)
);

BUFx6f_ASAP7_75t_L g3935 ( 
.A(n_3123),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3106),
.B(n_2275),
.Y(n_3936)
);

OAI21x1_ASAP7_75t_L g3937 ( 
.A1(n_3162),
.A2(n_2436),
.B(n_2428),
.Y(n_3937)
);

INVx1_ASAP7_75t_SL g3938 ( 
.A(n_3313),
.Y(n_3938)
);

OAI22xp5_ASAP7_75t_L g3939 ( 
.A1(n_3271),
.A2(n_2870),
.B1(n_3132),
.B2(n_2951),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3330),
.Y(n_3940)
);

OAI21x1_ASAP7_75t_L g3941 ( 
.A1(n_3162),
.A2(n_2436),
.B(n_2428),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3106),
.B(n_2275),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3114),
.B(n_2275),
.Y(n_3943)
);

AOI221xp5_ASAP7_75t_SL g3944 ( 
.A1(n_2888),
.A2(n_2344),
.B1(n_2283),
.B2(n_2280),
.C(n_2296),
.Y(n_3944)
);

AOI21xp5_ASAP7_75t_L g3945 ( 
.A1(n_3402),
.A2(n_3487),
.B(n_3525),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3495),
.B(n_3330),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3495),
.B(n_3271),
.Y(n_3947)
);

OAI21xp5_ASAP7_75t_L g3948 ( 
.A1(n_3514),
.A2(n_2870),
.B(n_3140),
.Y(n_3948)
);

O2A1O1Ixp33_ASAP7_75t_L g3949 ( 
.A1(n_3419),
.A2(n_3276),
.B(n_3080),
.C(n_3099),
.Y(n_3949)
);

OAI21x1_ASAP7_75t_L g3950 ( 
.A1(n_3543),
.A2(n_3207),
.B(n_3162),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3433),
.Y(n_3951)
);

OAI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_3419),
.A2(n_3140),
.B(n_3132),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3510),
.Y(n_3953)
);

BUFx3_ASAP7_75t_L g3954 ( 
.A(n_3726),
.Y(n_3954)
);

AOI21xp5_ASAP7_75t_L g3955 ( 
.A1(n_3402),
.A2(n_3341),
.B(n_3085),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3433),
.Y(n_3956)
);

BUFx2_ASAP7_75t_L g3957 ( 
.A(n_3405),
.Y(n_3957)
);

INVx4_ASAP7_75t_L g3958 ( 
.A(n_3726),
.Y(n_3958)
);

A2O1A1Ixp33_ASAP7_75t_L g3959 ( 
.A1(n_3441),
.A2(n_3213),
.B(n_3124),
.C(n_3378),
.Y(n_3959)
);

INVx2_ASAP7_75t_SL g3960 ( 
.A(n_3709),
.Y(n_3960)
);

OAI21x1_ASAP7_75t_L g3961 ( 
.A1(n_3543),
.A2(n_3207),
.B(n_3282),
.Y(n_3961)
);

A2O1A1Ixp33_ASAP7_75t_L g3962 ( 
.A1(n_3591),
.A2(n_3213),
.B(n_3292),
.C(n_3180),
.Y(n_3962)
);

INVxp67_ASAP7_75t_L g3963 ( 
.A(n_3440),
.Y(n_3963)
);

AOI21xp5_ASAP7_75t_L g3964 ( 
.A1(n_3487),
.A2(n_3085),
.B(n_3041),
.Y(n_3964)
);

INVx3_ASAP7_75t_L g3965 ( 
.A(n_3709),
.Y(n_3965)
);

NAND3xp33_ASAP7_75t_L g3966 ( 
.A(n_3461),
.B(n_3525),
.C(n_3674),
.Y(n_3966)
);

BUFx6f_ASAP7_75t_L g3967 ( 
.A(n_3418),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_L g3968 ( 
.A(n_3392),
.B(n_2858),
.Y(n_3968)
);

AOI21xp5_ASAP7_75t_L g3969 ( 
.A1(n_3420),
.A2(n_3476),
.B(n_3702),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3392),
.B(n_2858),
.Y(n_3970)
);

INVx3_ASAP7_75t_L g3971 ( 
.A(n_3709),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_3420),
.A2(n_3085),
.B(n_3041),
.Y(n_3972)
);

OAI21x1_ASAP7_75t_L g3973 ( 
.A1(n_3546),
.A2(n_3285),
.B(n_3282),
.Y(n_3973)
);

A2O1A1Ixp33_ASAP7_75t_L g3974 ( 
.A1(n_3439),
.A2(n_3213),
.B(n_3008),
.C(n_3384),
.Y(n_3974)
);

BUFx2_ASAP7_75t_L g3975 ( 
.A(n_3405),
.Y(n_3975)
);

OAI22xp5_ASAP7_75t_L g3976 ( 
.A1(n_3697),
.A2(n_3140),
.B1(n_3139),
.B2(n_3085),
.Y(n_3976)
);

OA21x2_ASAP7_75t_L g3977 ( 
.A1(n_3657),
.A2(n_3141),
.B(n_3075),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3469),
.Y(n_3978)
);

AOI31xp67_ASAP7_75t_L g3979 ( 
.A1(n_3632),
.A2(n_3174),
.A3(n_3089),
.B(n_3133),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3469),
.Y(n_3980)
);

CKINVDCx9p33_ASAP7_75t_R g3981 ( 
.A(n_3656),
.Y(n_3981)
);

AOI22xp33_ASAP7_75t_L g3982 ( 
.A1(n_3408),
.A2(n_2503),
.B1(n_2482),
.B2(n_3041),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3510),
.Y(n_3983)
);

CKINVDCx5p33_ASAP7_75t_R g3984 ( 
.A(n_3517),
.Y(n_3984)
);

AOI22xp33_ASAP7_75t_L g3985 ( 
.A1(n_3461),
.A2(n_2503),
.B1(n_2482),
.B2(n_3085),
.Y(n_3985)
);

CKINVDCx11_ASAP7_75t_R g3986 ( 
.A(n_3552),
.Y(n_3986)
);

OAI22xp5_ASAP7_75t_L g3987 ( 
.A1(n_3697),
.A2(n_3191),
.B1(n_2195),
.B2(n_2161),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3586),
.B(n_2960),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_L g3989 ( 
.A(n_3529),
.B(n_3228),
.Y(n_3989)
);

A2O1A1Ixp33_ASAP7_75t_L g3990 ( 
.A1(n_3475),
.A2(n_3008),
.B(n_3386),
.C(n_3077),
.Y(n_3990)
);

OA21x2_ASAP7_75t_L g3991 ( 
.A1(n_3657),
.A2(n_3435),
.B(n_3436),
.Y(n_3991)
);

BUFx3_ASAP7_75t_L g3992 ( 
.A(n_3726),
.Y(n_3992)
);

BUFx6f_ASAP7_75t_L g3993 ( 
.A(n_3418),
.Y(n_3993)
);

OAI21x1_ASAP7_75t_L g3994 ( 
.A1(n_3546),
.A2(n_3476),
.B(n_3648),
.Y(n_3994)
);

INVx3_ASAP7_75t_L g3995 ( 
.A(n_3709),
.Y(n_3995)
);

OAI21x1_ASAP7_75t_L g3996 ( 
.A1(n_3648),
.A2(n_3285),
.B(n_3282),
.Y(n_3996)
);

INVx3_ASAP7_75t_L g3997 ( 
.A(n_3935),
.Y(n_3997)
);

BUFx4_ASAP7_75t_SL g3998 ( 
.A(n_3572),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3470),
.Y(n_3999)
);

AOI21xp5_ASAP7_75t_L g4000 ( 
.A1(n_3475),
.A2(n_3145),
.B(n_3123),
.Y(n_4000)
);

INVxp67_ASAP7_75t_L g4001 ( 
.A(n_3474),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_3529),
.B(n_3228),
.Y(n_4002)
);

OAI21xp5_ASAP7_75t_L g4003 ( 
.A1(n_3493),
.A2(n_3174),
.B(n_3181),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3584),
.B(n_3104),
.Y(n_4004)
);

AO32x2_ASAP7_75t_L g4005 ( 
.A1(n_3688),
.A2(n_3205),
.A3(n_3232),
.B1(n_3025),
.B2(n_2831),
.Y(n_4005)
);

INVx2_ASAP7_75t_L g4006 ( 
.A(n_3510),
.Y(n_4006)
);

INVx4_ASAP7_75t_L g4007 ( 
.A(n_3771),
.Y(n_4007)
);

AOI21xp5_ASAP7_75t_L g4008 ( 
.A1(n_3481),
.A2(n_3145),
.B(n_3123),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3584),
.B(n_3104),
.Y(n_4009)
);

HB1xp67_ASAP7_75t_L g4010 ( 
.A(n_3775),
.Y(n_4010)
);

AOI21xp33_ASAP7_75t_L g4011 ( 
.A1(n_3674),
.A2(n_3174),
.B(n_3211),
.Y(n_4011)
);

NOR4xp25_ASAP7_75t_L g4012 ( 
.A(n_3493),
.B(n_3186),
.C(n_2923),
.D(n_2926),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3400),
.B(n_2960),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3470),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_3481),
.A2(n_3145),
.B(n_2238),
.Y(n_4015)
);

OAI22x1_ASAP7_75t_L g4016 ( 
.A1(n_3745),
.A2(n_3285),
.B1(n_3299),
.B2(n_3282),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_3848),
.A2(n_3145),
.B(n_2238),
.Y(n_4017)
);

OA21x2_ASAP7_75t_L g4018 ( 
.A1(n_3435),
.A2(n_3190),
.B(n_3001),
.Y(n_4018)
);

NAND2xp5_ASAP7_75t_SL g4019 ( 
.A(n_3681),
.B(n_2913),
.Y(n_4019)
);

NAND2xp5_ASAP7_75t_L g4020 ( 
.A(n_3400),
.B(n_3033),
.Y(n_4020)
);

OAI22xp5_ASAP7_75t_L g4021 ( 
.A1(n_3770),
.A2(n_3191),
.B1(n_2195),
.B2(n_2161),
.Y(n_4021)
);

OAI21x1_ASAP7_75t_L g4022 ( 
.A1(n_3519),
.A2(n_3299),
.B(n_3285),
.Y(n_4022)
);

INVx1_ASAP7_75t_SL g4023 ( 
.A(n_3705),
.Y(n_4023)
);

OAI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_3450),
.A2(n_2920),
.B(n_3028),
.Y(n_4024)
);

A2O1A1Ixp33_ASAP7_75t_L g4025 ( 
.A1(n_3490),
.A2(n_3077),
.B(n_3119),
.C(n_3005),
.Y(n_4025)
);

OR2x2_ASAP7_75t_L g4026 ( 
.A(n_3456),
.B(n_3143),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_SL g4027 ( 
.A1(n_3895),
.A2(n_3077),
.B(n_3005),
.Y(n_4027)
);

INVx1_ASAP7_75t_SL g4028 ( 
.A(n_3705),
.Y(n_4028)
);

OAI21xp5_ASAP7_75t_L g4029 ( 
.A1(n_3450),
.A2(n_3021),
.B(n_3018),
.Y(n_4029)
);

BUFx3_ASAP7_75t_L g4030 ( 
.A(n_3771),
.Y(n_4030)
);

AOI22xp5_ASAP7_75t_L g4031 ( 
.A1(n_3695),
.A2(n_2482),
.B1(n_2503),
.B2(n_2327),
.Y(n_4031)
);

OAI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_3631),
.A2(n_3047),
.B(n_3046),
.Y(n_4032)
);

A2O1A1Ixp33_ASAP7_75t_L g4033 ( 
.A1(n_3490),
.A2(n_3119),
.B(n_3324),
.C(n_3277),
.Y(n_4033)
);

BUFx10_ASAP7_75t_L g4034 ( 
.A(n_3477),
.Y(n_4034)
);

NOR2xp33_ASAP7_75t_L g4035 ( 
.A(n_3447),
.B(n_2853),
.Y(n_4035)
);

BUFx10_ASAP7_75t_L g4036 ( 
.A(n_3428),
.Y(n_4036)
);

A2O1A1Ixp33_ASAP7_75t_L g4037 ( 
.A1(n_3878),
.A2(n_3119),
.B(n_3324),
.C(n_3277),
.Y(n_4037)
);

NAND2xp5_ASAP7_75t_L g4038 ( 
.A(n_3401),
.B(n_3033),
.Y(n_4038)
);

A2O1A1Ixp33_ASAP7_75t_L g4039 ( 
.A1(n_3878),
.A2(n_3277),
.B(n_3324),
.C(n_3042),
.Y(n_4039)
);

INVxp67_ASAP7_75t_SL g4040 ( 
.A(n_3692),
.Y(n_4040)
);

AOI21xp5_ASAP7_75t_L g4041 ( 
.A1(n_3848),
.A2(n_3145),
.B(n_2238),
.Y(n_4041)
);

OAI21x1_ASAP7_75t_L g4042 ( 
.A1(n_3519),
.A2(n_3306),
.B(n_3299),
.Y(n_4042)
);

O2A1O1Ixp33_ASAP7_75t_L g4043 ( 
.A1(n_3448),
.A2(n_2949),
.B(n_3198),
.C(n_3195),
.Y(n_4043)
);

AO32x1_ASAP7_75t_L g4044 ( 
.A1(n_3410),
.A2(n_3205),
.A3(n_3025),
.B1(n_3232),
.B2(n_2831),
.Y(n_4044)
);

NAND3xp33_ASAP7_75t_SL g4045 ( 
.A(n_3819),
.B(n_3017),
.C(n_3016),
.Y(n_4045)
);

HB1xp67_ASAP7_75t_L g4046 ( 
.A(n_3781),
.Y(n_4046)
);

INVxp67_ASAP7_75t_L g4047 ( 
.A(n_3833),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3401),
.B(n_3172),
.Y(n_4048)
);

AOI22xp5_ASAP7_75t_L g4049 ( 
.A1(n_3695),
.A2(n_2482),
.B1(n_2503),
.B2(n_2327),
.Y(n_4049)
);

OAI21x1_ASAP7_75t_L g4050 ( 
.A1(n_3732),
.A2(n_3306),
.B(n_3299),
.Y(n_4050)
);

NOR2xp33_ASAP7_75t_L g4051 ( 
.A(n_3617),
.B(n_2853),
.Y(n_4051)
);

OAI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_3631),
.A2(n_3048),
.B(n_3060),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3586),
.B(n_3306),
.Y(n_4053)
);

BUFx3_ASAP7_75t_L g4054 ( 
.A(n_3771),
.Y(n_4054)
);

AOI21xp5_ASAP7_75t_L g4055 ( 
.A1(n_3484),
.A2(n_2238),
.B(n_2225),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3485),
.B(n_3172),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3485),
.B(n_3172),
.Y(n_4057)
);

OAI21x1_ASAP7_75t_L g4058 ( 
.A1(n_3732),
.A2(n_3316),
.B(n_3306),
.Y(n_4058)
);

CKINVDCx5p33_ASAP7_75t_R g4059 ( 
.A(n_3566),
.Y(n_4059)
);

NOR2xp33_ASAP7_75t_L g4060 ( 
.A(n_3478),
.B(n_3009),
.Y(n_4060)
);

AND2x4_ASAP7_75t_L g4061 ( 
.A(n_3875),
.B(n_3316),
.Y(n_4061)
);

AOI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_3807),
.A2(n_2238),
.B(n_2225),
.Y(n_4062)
);

AO32x2_ASAP7_75t_L g4063 ( 
.A1(n_3688),
.A2(n_3342),
.A3(n_2301),
.B1(n_2208),
.B2(n_2313),
.Y(n_4063)
);

NOR2xp33_ASAP7_75t_L g4064 ( 
.A(n_3547),
.B(n_3009),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_L g4065 ( 
.A(n_3403),
.B(n_3172),
.Y(n_4065)
);

INVx2_ASAP7_75t_L g4066 ( 
.A(n_3520),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3403),
.B(n_3114),
.Y(n_4067)
);

OAI21xp5_ASAP7_75t_L g4068 ( 
.A1(n_3891),
.A2(n_3065),
.B(n_3142),
.Y(n_4068)
);

AOI21xp5_ASAP7_75t_L g4069 ( 
.A1(n_3807),
.A2(n_2241),
.B(n_2238),
.Y(n_4069)
);

AOI31xp67_ASAP7_75t_L g4070 ( 
.A1(n_3926),
.A2(n_3220),
.A3(n_3224),
.B(n_3185),
.Y(n_4070)
);

OR2x2_ASAP7_75t_L g4071 ( 
.A(n_3456),
.B(n_3297),
.Y(n_4071)
);

INVx2_ASAP7_75t_L g4072 ( 
.A(n_3520),
.Y(n_4072)
);

NOR2xp33_ASAP7_75t_L g4073 ( 
.A(n_3703),
.B(n_3009),
.Y(n_4073)
);

BUFx6f_ASAP7_75t_L g4074 ( 
.A(n_3418),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3520),
.Y(n_4075)
);

BUFx2_ASAP7_75t_L g4076 ( 
.A(n_3405),
.Y(n_4076)
);

AOI21xp5_ASAP7_75t_L g4077 ( 
.A1(n_3729),
.A2(n_2241),
.B(n_2238),
.Y(n_4077)
);

NAND3xp33_ASAP7_75t_L g4078 ( 
.A(n_3819),
.B(n_3009),
.C(n_2349),
.Y(n_4078)
);

HB1xp67_ASAP7_75t_L g4079 ( 
.A(n_3781),
.Y(n_4079)
);

NOR2x1_ASAP7_75t_L g4080 ( 
.A(n_3862),
.B(n_3332),
.Y(n_4080)
);

NOR2xp33_ASAP7_75t_SL g4081 ( 
.A(n_3672),
.B(n_2349),
.Y(n_4081)
);

INVx2_ASAP7_75t_L g4082 ( 
.A(n_3522),
.Y(n_4082)
);

BUFx2_ASAP7_75t_L g4083 ( 
.A(n_3405),
.Y(n_4083)
);

INVx3_ASAP7_75t_SL g4084 ( 
.A(n_3660),
.Y(n_4084)
);

BUFx6f_ASAP7_75t_L g4085 ( 
.A(n_3471),
.Y(n_4085)
);

O2A1O1Ixp33_ASAP7_75t_L g4086 ( 
.A1(n_3891),
.A2(n_3081),
.B(n_3130),
.C(n_3127),
.Y(n_4086)
);

INVx2_ASAP7_75t_L g4087 ( 
.A(n_3522),
.Y(n_4087)
);

OAI21xp5_ASAP7_75t_L g4088 ( 
.A1(n_3811),
.A2(n_3093),
.B(n_3161),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3480),
.Y(n_4089)
);

INVx1_ASAP7_75t_L g4090 ( 
.A(n_3480),
.Y(n_4090)
);

INVx4_ASAP7_75t_L g4091 ( 
.A(n_3471),
.Y(n_4091)
);

CKINVDCx11_ASAP7_75t_R g4092 ( 
.A(n_3552),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3791),
.B(n_3427),
.Y(n_4093)
);

O2A1O1Ixp33_ASAP7_75t_L g4094 ( 
.A1(n_3396),
.A2(n_3173),
.B(n_3175),
.C(n_3168),
.Y(n_4094)
);

INVx3_ASAP7_75t_L g4095 ( 
.A(n_3700),
.Y(n_4095)
);

AOI21xp5_ASAP7_75t_L g4096 ( 
.A1(n_3743),
.A2(n_2241),
.B(n_2238),
.Y(n_4096)
);

O2A1O1Ixp5_ASAP7_75t_SL g4097 ( 
.A1(n_3578),
.A2(n_3383),
.B(n_3001),
.C(n_3019),
.Y(n_4097)
);

INVx1_ASAP7_75t_L g4098 ( 
.A(n_3492),
.Y(n_4098)
);

AOI21x1_ASAP7_75t_L g4099 ( 
.A1(n_3699),
.A2(n_2450),
.B(n_2448),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_3743),
.A2(n_2241),
.B(n_2238),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3492),
.Y(n_4101)
);

OAI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_3811),
.A2(n_3182),
.B(n_3111),
.Y(n_4102)
);

OAI22xp5_ASAP7_75t_L g4103 ( 
.A1(n_3770),
.A2(n_3191),
.B1(n_2185),
.B2(n_2231),
.Y(n_4103)
);

OAI21x1_ASAP7_75t_L g4104 ( 
.A1(n_3467),
.A2(n_3359),
.B(n_2455),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3494),
.Y(n_4105)
);

INVx2_ASAP7_75t_L g4106 ( 
.A(n_3522),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3791),
.B(n_3156),
.Y(n_4107)
);

A2O1A1Ixp33_ASAP7_75t_L g4108 ( 
.A1(n_3554),
.A2(n_2250),
.B(n_2316),
.C(n_2241),
.Y(n_4108)
);

CKINVDCx11_ASAP7_75t_R g4109 ( 
.A(n_3552),
.Y(n_4109)
);

AOI21xp5_ASAP7_75t_L g4110 ( 
.A1(n_3792),
.A2(n_2250),
.B(n_2241),
.Y(n_4110)
);

AOI22xp5_ASAP7_75t_L g4111 ( 
.A1(n_3410),
.A2(n_2482),
.B1(n_2503),
.B2(n_2327),
.Y(n_4111)
);

AOI21xp33_ASAP7_75t_L g4112 ( 
.A1(n_3526),
.A2(n_3206),
.B(n_3118),
.Y(n_4112)
);

AOI21xp5_ASAP7_75t_L g4113 ( 
.A1(n_3792),
.A2(n_2250),
.B(n_2241),
.Y(n_4113)
);

INVx1_ASAP7_75t_L g4114 ( 
.A(n_3494),
.Y(n_4114)
);

NOR2x1_ASAP7_75t_R g4115 ( 
.A(n_3841),
.B(n_2738),
.Y(n_4115)
);

NOR2xp33_ASAP7_75t_L g4116 ( 
.A(n_3570),
.B(n_2503),
.Y(n_4116)
);

AND2x4_ASAP7_75t_L g4117 ( 
.A(n_3875),
.B(n_2241),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_L g4118 ( 
.A(n_3427),
.B(n_3409),
.Y(n_4118)
);

O2A1O1Ixp33_ASAP7_75t_L g4119 ( 
.A1(n_3394),
.A2(n_3108),
.B(n_3121),
.C(n_3226),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3409),
.B(n_3156),
.Y(n_4120)
);

AO31x2_ASAP7_75t_L g4121 ( 
.A1(n_3619),
.A2(n_3383),
.A3(n_3381),
.B(n_3196),
.Y(n_4121)
);

OAI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_3569),
.A2(n_3221),
.B(n_3212),
.Y(n_4122)
);

INVx3_ASAP7_75t_L g4123 ( 
.A(n_3935),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3711),
.B(n_3176),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_L g4125 ( 
.A(n_3488),
.B(n_3176),
.Y(n_4125)
);

AO21x1_ASAP7_75t_L g4126 ( 
.A1(n_3578),
.A2(n_2283),
.B(n_2280),
.Y(n_4126)
);

BUFx3_ASAP7_75t_L g4127 ( 
.A(n_3471),
.Y(n_4127)
);

O2A1O1Ixp33_ASAP7_75t_L g4128 ( 
.A1(n_3394),
.A2(n_3229),
.B(n_3206),
.C(n_2738),
.Y(n_4128)
);

BUFx6f_ASAP7_75t_L g4129 ( 
.A(n_3652),
.Y(n_4129)
);

AOI21x1_ASAP7_75t_L g4130 ( 
.A1(n_3699),
.A2(n_2477),
.B(n_2473),
.Y(n_4130)
);

AND2x4_ASAP7_75t_L g4131 ( 
.A(n_3875),
.B(n_2241),
.Y(n_4131)
);

O2A1O1Ixp5_ASAP7_75t_L g4132 ( 
.A1(n_3650),
.A2(n_3381),
.B(n_3039),
.C(n_3032),
.Y(n_4132)
);

AOI21xp5_ASAP7_75t_L g4133 ( 
.A1(n_3803),
.A2(n_2316),
.B(n_2250),
.Y(n_4133)
);

NAND3xp33_ASAP7_75t_SL g4134 ( 
.A(n_3533),
.B(n_2283),
.C(n_2280),
.Y(n_4134)
);

AO31x2_ASAP7_75t_L g4135 ( 
.A1(n_3622),
.A2(n_3083),
.A3(n_3354),
.B(n_2997),
.Y(n_4135)
);

CKINVDCx5p33_ASAP7_75t_R g4136 ( 
.A(n_3559),
.Y(n_4136)
);

OAI22xp5_ASAP7_75t_L g4137 ( 
.A1(n_3672),
.A2(n_2185),
.B1(n_2205),
.B2(n_2399),
.Y(n_4137)
);

AOI21xp5_ASAP7_75t_L g4138 ( 
.A1(n_3803),
.A2(n_2316),
.B(n_2250),
.Y(n_4138)
);

AOI21xp5_ASAP7_75t_L g4139 ( 
.A1(n_3557),
.A2(n_2316),
.B(n_2250),
.Y(n_4139)
);

OAI22x1_ASAP7_75t_L g4140 ( 
.A1(n_3745),
.A2(n_3257),
.B1(n_3129),
.B2(n_3126),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_L g4141 ( 
.A(n_3488),
.B(n_3178),
.Y(n_4141)
);

AOI22xp5_ASAP7_75t_L g4142 ( 
.A1(n_3853),
.A2(n_2327),
.B1(n_2368),
.B2(n_2805),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3563),
.B(n_3178),
.Y(n_4143)
);

CKINVDCx5p33_ASAP7_75t_R g4144 ( 
.A(n_3615),
.Y(n_4144)
);

AO22x2_ASAP7_75t_L g4145 ( 
.A1(n_3404),
.A2(n_3019),
.B1(n_3354),
.B2(n_3029),
.Y(n_4145)
);

HB1xp67_ASAP7_75t_L g4146 ( 
.A(n_3915),
.Y(n_4146)
);

AO22x1_ASAP7_75t_L g4147 ( 
.A1(n_3680),
.A2(n_2349),
.B1(n_2316),
.B2(n_2250),
.Y(n_4147)
);

AOI21xp5_ASAP7_75t_L g4148 ( 
.A1(n_3564),
.A2(n_2340),
.B(n_2250),
.Y(n_4148)
);

NOR2xp33_ASAP7_75t_L g4149 ( 
.A(n_3597),
.B(n_2913),
.Y(n_4149)
);

O2A1O1Ixp33_ASAP7_75t_L g4150 ( 
.A1(n_3534),
.A2(n_2738),
.B(n_2344),
.C(n_2381),
.Y(n_4150)
);

AO31x2_ASAP7_75t_L g4151 ( 
.A1(n_3622),
.A2(n_3196),
.A3(n_3126),
.B(n_3129),
.Y(n_4151)
);

OAI21xp5_ASAP7_75t_L g4152 ( 
.A1(n_3651),
.A2(n_2813),
.B(n_2812),
.Y(n_4152)
);

OAI22xp5_ASAP7_75t_L g4153 ( 
.A1(n_3777),
.A2(n_2205),
.B1(n_2399),
.B2(n_2231),
.Y(n_4153)
);

OAI22xp5_ASAP7_75t_L g4154 ( 
.A1(n_3777),
.A2(n_2205),
.B1(n_2399),
.B2(n_2231),
.Y(n_4154)
);

AOI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_3887),
.A2(n_2340),
.B(n_2250),
.Y(n_4155)
);

AO21x2_ASAP7_75t_L g4156 ( 
.A1(n_3627),
.A2(n_3039),
.B(n_3032),
.Y(n_4156)
);

NOR2xp33_ASAP7_75t_L g4157 ( 
.A(n_3597),
.B(n_2913),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3563),
.B(n_3218),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_3501),
.Y(n_4159)
);

AO31x2_ASAP7_75t_L g4160 ( 
.A1(n_3627),
.A2(n_3628),
.A3(n_3612),
.B(n_3533),
.Y(n_4160)
);

NAND2xp5_ASAP7_75t_L g4161 ( 
.A(n_3621),
.B(n_3218),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_3887),
.A2(n_2364),
.B(n_2340),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3621),
.B(n_2866),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3501),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_3593),
.A2(n_2364),
.B(n_2340),
.Y(n_4165)
);

AOI221x1_ASAP7_75t_L g4166 ( 
.A1(n_3675),
.A2(n_3164),
.B1(n_3062),
.B2(n_3257),
.C(n_3101),
.Y(n_4166)
);

AOI21xp5_ASAP7_75t_SL g4167 ( 
.A1(n_3897),
.A2(n_2364),
.B(n_2340),
.Y(n_4167)
);

A2O1A1Ixp33_ASAP7_75t_L g4168 ( 
.A1(n_3712),
.A2(n_2372),
.B(n_2364),
.C(n_2231),
.Y(n_4168)
);

AND2x4_ASAP7_75t_L g4169 ( 
.A(n_3875),
.B(n_2364),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3804),
.B(n_2866),
.Y(n_4170)
);

NOR2xp33_ASAP7_75t_L g4171 ( 
.A(n_3597),
.B(n_2913),
.Y(n_4171)
);

AOI21xp33_ASAP7_75t_L g4172 ( 
.A1(n_3526),
.A2(n_2372),
.B(n_2364),
.Y(n_4172)
);

O2A1O1Ixp33_ASAP7_75t_SL g4173 ( 
.A1(n_3816),
.A2(n_2304),
.B(n_2352),
.C(n_2392),
.Y(n_4173)
);

AOI21xp33_ASAP7_75t_L g4174 ( 
.A1(n_3760),
.A2(n_3605),
.B(n_3482),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_3509),
.Y(n_4175)
);

AO31x2_ASAP7_75t_L g4176 ( 
.A1(n_3628),
.A2(n_3136),
.A3(n_3148),
.B(n_3163),
.Y(n_4176)
);

NOR4xp25_ASAP7_75t_L g4177 ( 
.A(n_3715),
.B(n_2381),
.C(n_2304),
.D(n_2291),
.Y(n_4177)
);

AO21x1_ASAP7_75t_L g4178 ( 
.A1(n_3675),
.A2(n_3086),
.B(n_3059),
.Y(n_4178)
);

AOI21xp5_ASAP7_75t_L g4179 ( 
.A1(n_3587),
.A2(n_2372),
.B(n_2364),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_3804),
.B(n_2902),
.Y(n_4180)
);

OAI21x1_ASAP7_75t_L g4181 ( 
.A1(n_3735),
.A2(n_3026),
.B(n_2955),
.Y(n_4181)
);

NAND2xp5_ASAP7_75t_L g4182 ( 
.A(n_3542),
.B(n_2902),
.Y(n_4182)
);

NAND3xp33_ASAP7_75t_SL g4183 ( 
.A(n_3592),
.B(n_3101),
.C(n_3086),
.Y(n_4183)
);

NAND3xp33_ASAP7_75t_L g4184 ( 
.A(n_3576),
.B(n_2930),
.C(n_2927),
.Y(n_4184)
);

OAI21xp5_ASAP7_75t_L g4185 ( 
.A1(n_3639),
.A2(n_2813),
.B(n_2812),
.Y(n_4185)
);

OAI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3639),
.A2(n_2813),
.B(n_2812),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_3509),
.Y(n_4187)
);

BUFx12f_ASAP7_75t_L g4188 ( 
.A(n_3434),
.Y(n_4188)
);

AO31x2_ASAP7_75t_L g4189 ( 
.A1(n_3612),
.A2(n_3901),
.A3(n_3592),
.B(n_3636),
.Y(n_4189)
);

NOR2xp67_ASAP7_75t_L g4190 ( 
.A(n_3406),
.B(n_3136),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_3542),
.B(n_3035),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_3865),
.B(n_3035),
.Y(n_4192)
);

AOI21xp5_ASAP7_75t_L g4193 ( 
.A1(n_3590),
.A2(n_3541),
.B(n_3571),
.Y(n_4193)
);

INVx3_ASAP7_75t_SL g4194 ( 
.A(n_3678),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3865),
.B(n_3053),
.Y(n_4195)
);

BUFx4f_ASAP7_75t_SL g4196 ( 
.A(n_3673),
.Y(n_4196)
);

AND2x2_ASAP7_75t_L g4197 ( 
.A(n_3496),
.B(n_3148),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_3513),
.Y(n_4198)
);

NOR2xp33_ASAP7_75t_L g4199 ( 
.A(n_3707),
.B(n_2927),
.Y(n_4199)
);

OAI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_3421),
.A2(n_2205),
.B1(n_2399),
.B2(n_2254),
.Y(n_4200)
);

INVx1_ASAP7_75t_L g4201 ( 
.A(n_3513),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_3535),
.Y(n_4202)
);

OAI21x1_ASAP7_75t_L g4203 ( 
.A1(n_3757),
.A2(n_3515),
.B(n_3512),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3544),
.B(n_3567),
.Y(n_4204)
);

OAI21x1_ASAP7_75t_L g4205 ( 
.A1(n_3757),
.A2(n_3515),
.B(n_3512),
.Y(n_4205)
);

AOI21xp5_ASAP7_75t_L g4206 ( 
.A1(n_3541),
.A2(n_2372),
.B(n_2364),
.Y(n_4206)
);

OAI21xp5_ASAP7_75t_L g4207 ( 
.A1(n_3576),
.A2(n_2813),
.B(n_2812),
.Y(n_4207)
);

OAI22xp5_ASAP7_75t_L g4208 ( 
.A1(n_3421),
.A2(n_2369),
.B1(n_2254),
.B2(n_2274),
.Y(n_4208)
);

AOI21xp5_ASAP7_75t_L g4209 ( 
.A1(n_3594),
.A2(n_2372),
.B(n_2364),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_3496),
.B(n_3499),
.Y(n_4210)
);

AO21x1_ASAP7_75t_L g4211 ( 
.A1(n_3939),
.A2(n_3296),
.B(n_3279),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_3784),
.B(n_2927),
.Y(n_4212)
);

AO31x2_ASAP7_75t_L g4213 ( 
.A1(n_3636),
.A2(n_3279),
.A3(n_3296),
.B(n_3336),
.Y(n_4213)
);

AOI21xp5_ASAP7_75t_L g4214 ( 
.A1(n_3585),
.A2(n_2208),
.B(n_2313),
.Y(n_4214)
);

OAI21x1_ASAP7_75t_L g4215 ( 
.A1(n_3516),
.A2(n_3380),
.B(n_3026),
.Y(n_4215)
);

AOI21xp5_ASAP7_75t_L g4216 ( 
.A1(n_3585),
.A2(n_2208),
.B(n_2313),
.Y(n_4216)
);

AOI21xp5_ASAP7_75t_L g4217 ( 
.A1(n_3545),
.A2(n_3683),
.B(n_3511),
.Y(n_4217)
);

OAI22xp5_ASAP7_75t_SL g4218 ( 
.A1(n_3853),
.A2(n_3704),
.B1(n_3404),
.B2(n_3673),
.Y(n_4218)
);

OA21x2_ASAP7_75t_L g4219 ( 
.A1(n_3637),
.A2(n_3320),
.B(n_3331),
.Y(n_4219)
);

NOR2xp33_ASAP7_75t_L g4220 ( 
.A(n_3693),
.B(n_2927),
.Y(n_4220)
);

OR2x6_ASAP7_75t_L g4221 ( 
.A(n_3556),
.B(n_2748),
.Y(n_4221)
);

OAI22x1_ASAP7_75t_L g4222 ( 
.A1(n_3539),
.A2(n_3602),
.B1(n_3896),
.B2(n_3763),
.Y(n_4222)
);

A2O1A1Ixp33_ASAP7_75t_L g4223 ( 
.A1(n_3715),
.A2(n_2334),
.B(n_2254),
.C(n_2274),
.Y(n_4223)
);

AND2x2_ASAP7_75t_L g4224 ( 
.A(n_3499),
.B(n_3049),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_L g4225 ( 
.A(n_3866),
.B(n_2927),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_3535),
.Y(n_4226)
);

OR2x2_ASAP7_75t_L g4227 ( 
.A(n_3465),
.B(n_3049),
.Y(n_4227)
);

AOI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_3443),
.A2(n_2368),
.B1(n_2805),
.B2(n_2498),
.Y(n_4228)
);

INVx1_ASAP7_75t_L g4229 ( 
.A(n_3565),
.Y(n_4229)
);

O2A1O1Ixp33_ASAP7_75t_SL g4230 ( 
.A1(n_3395),
.A2(n_2632),
.B(n_2719),
.C(n_2727),
.Y(n_4230)
);

INVx3_ASAP7_75t_L g4231 ( 
.A(n_3700),
.Y(n_4231)
);

AOI21x1_ASAP7_75t_L g4232 ( 
.A1(n_3574),
.A2(n_3194),
.B(n_3107),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_3565),
.Y(n_4233)
);

AOI21xp5_ASAP7_75t_L g4234 ( 
.A1(n_3683),
.A2(n_2301),
.B(n_2313),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3518),
.B(n_3125),
.Y(n_4235)
);

OAI21x1_ASAP7_75t_L g4236 ( 
.A1(n_3532),
.A2(n_2427),
.B(n_2414),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3583),
.Y(n_4237)
);

INVx3_ASAP7_75t_L g4238 ( 
.A(n_3700),
.Y(n_4238)
);

OAI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_3596),
.A2(n_3629),
.B(n_3614),
.Y(n_4239)
);

AOI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_3511),
.A2(n_2301),
.B(n_2313),
.Y(n_4240)
);

OAI21xp5_ASAP7_75t_L g4241 ( 
.A1(n_3596),
.A2(n_3629),
.B(n_3614),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_3544),
.B(n_3053),
.Y(n_4242)
);

NAND2x1p5_ASAP7_75t_L g4243 ( 
.A(n_3679),
.B(n_2748),
.Y(n_4243)
);

OR2x2_ASAP7_75t_L g4244 ( 
.A(n_3465),
.B(n_3064),
.Y(n_4244)
);

INVxp67_ASAP7_75t_L g4245 ( 
.A(n_3800),
.Y(n_4245)
);

AOI22xp5_ASAP7_75t_L g4246 ( 
.A1(n_3497),
.A2(n_2368),
.B1(n_2594),
.B2(n_2413),
.Y(n_4246)
);

BUFx6f_ASAP7_75t_L g4247 ( 
.A(n_3652),
.Y(n_4247)
);

INVx1_ASAP7_75t_L g4248 ( 
.A(n_3583),
.Y(n_4248)
);

AO32x2_ASAP7_75t_L g4249 ( 
.A1(n_3903),
.A2(n_3342),
.A3(n_2301),
.B1(n_2727),
.B2(n_2707),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_3623),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_SL g4251 ( 
.A(n_3689),
.B(n_2930),
.Y(n_4251)
);

BUFx3_ASAP7_75t_L g4252 ( 
.A(n_3652),
.Y(n_4252)
);

AO22x2_ASAP7_75t_L g4253 ( 
.A1(n_3903),
.A2(n_3064),
.B1(n_2716),
.B2(n_2738),
.Y(n_4253)
);

NAND2xp5_ASAP7_75t_L g4254 ( 
.A(n_3567),
.B(n_2930),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_3518),
.B(n_2930),
.Y(n_4255)
);

NAND2xp5_ASAP7_75t_L g4256 ( 
.A(n_3609),
.B(n_2930),
.Y(n_4256)
);

NAND2xp5_ASAP7_75t_L g4257 ( 
.A(n_3609),
.B(n_2945),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_3502),
.B(n_2945),
.Y(n_4258)
);

AOI21xp5_ASAP7_75t_L g4259 ( 
.A1(n_3725),
.A2(n_2301),
.B(n_2719),
.Y(n_4259)
);

AO31x2_ASAP7_75t_L g4260 ( 
.A1(n_3645),
.A2(n_2427),
.A3(n_2414),
.B(n_2400),
.Y(n_4260)
);

AOI21xp5_ASAP7_75t_L g4261 ( 
.A1(n_3725),
.A2(n_2632),
.B(n_2691),
.Y(n_4261)
);

BUFx10_ASAP7_75t_L g4262 ( 
.A(n_3428),
.Y(n_4262)
);

NAND2xp33_ASAP7_75t_SL g4263 ( 
.A(n_3414),
.B(n_2945),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3502),
.B(n_2945),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_3783),
.A2(n_2719),
.B(n_2707),
.Y(n_4265)
);

AO31x2_ASAP7_75t_L g4266 ( 
.A1(n_3645),
.A2(n_2427),
.A3(n_2414),
.B(n_2400),
.Y(n_4266)
);

AOI21xp5_ASAP7_75t_L g4267 ( 
.A1(n_3783),
.A2(n_2707),
.B(n_2727),
.Y(n_4267)
);

AOI21xp5_ASAP7_75t_L g4268 ( 
.A1(n_3412),
.A2(n_2691),
.B(n_2767),
.Y(n_4268)
);

OAI21x1_ASAP7_75t_L g4269 ( 
.A1(n_3553),
.A2(n_2414),
.B(n_2400),
.Y(n_4269)
);

BUFx8_ASAP7_75t_L g4270 ( 
.A(n_3673),
.Y(n_4270)
);

AO31x2_ASAP7_75t_L g4271 ( 
.A1(n_3752),
.A2(n_3755),
.A3(n_3932),
.B(n_3637),
.Y(n_4271)
);

AO31x2_ASAP7_75t_L g4272 ( 
.A1(n_3752),
.A2(n_2400),
.A3(n_2811),
.B(n_2807),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_3507),
.B(n_2945),
.Y(n_4273)
);

BUFx2_ASAP7_75t_L g4274 ( 
.A(n_3405),
.Y(n_4274)
);

AO21x1_ASAP7_75t_L g4275 ( 
.A1(n_3939),
.A2(n_2758),
.B(n_2775),
.Y(n_4275)
);

NOR2xp33_ASAP7_75t_L g4276 ( 
.A(n_3839),
.B(n_3870),
.Y(n_4276)
);

BUFx3_ASAP7_75t_L g4277 ( 
.A(n_3686),
.Y(n_4277)
);

NAND2xp5_ASAP7_75t_L g4278 ( 
.A(n_3507),
.B(n_3040),
.Y(n_4278)
);

NAND3xp33_ASAP7_75t_SL g4279 ( 
.A(n_3599),
.B(n_2758),
.C(n_2775),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_3623),
.Y(n_4280)
);

AOI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_3412),
.A2(n_2767),
.B(n_2750),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_L g4282 ( 
.A(n_3689),
.B(n_3040),
.Y(n_4282)
);

AO31x2_ASAP7_75t_L g4283 ( 
.A1(n_3755),
.A2(n_2630),
.A3(n_2811),
.B(n_2807),
.Y(n_4283)
);

OAI21x1_ASAP7_75t_L g4284 ( 
.A1(n_3553),
.A2(n_2630),
.B(n_2811),
.Y(n_4284)
);

AOI21xp5_ASAP7_75t_L g4285 ( 
.A1(n_3779),
.A2(n_2767),
.B(n_2750),
.Y(n_4285)
);

OAI21x1_ASAP7_75t_L g4286 ( 
.A1(n_3690),
.A2(n_2630),
.B(n_2811),
.Y(n_4286)
);

O2A1O1Ixp33_ASAP7_75t_SL g4287 ( 
.A1(n_3812),
.A2(n_2758),
.B(n_2775),
.C(n_2778),
.Y(n_4287)
);

AND2x4_ASAP7_75t_L g4288 ( 
.A(n_3875),
.B(n_2748),
.Y(n_4288)
);

NOR2xp33_ASAP7_75t_L g4289 ( 
.A(n_3689),
.B(n_3040),
.Y(n_4289)
);

A2O1A1Ixp33_ASAP7_75t_L g4290 ( 
.A1(n_3608),
.A2(n_2254),
.B(n_2274),
.C(n_2277),
.Y(n_4290)
);

BUFx10_ASAP7_75t_L g4291 ( 
.A(n_3428),
.Y(n_4291)
);

NAND2xp5_ASAP7_75t_L g4292 ( 
.A(n_3573),
.B(n_3040),
.Y(n_4292)
);

AO31x2_ASAP7_75t_L g4293 ( 
.A1(n_3932),
.A2(n_2709),
.A3(n_2807),
.B(n_2796),
.Y(n_4293)
);

NOR2xp33_ASAP7_75t_L g4294 ( 
.A(n_3689),
.B(n_3040),
.Y(n_4294)
);

NAND2xp5_ASAP7_75t_L g4295 ( 
.A(n_3573),
.B(n_3068),
.Y(n_4295)
);

AO32x2_ASAP7_75t_L g4296 ( 
.A1(n_3438),
.A2(n_2528),
.A3(n_2542),
.B1(n_2595),
.B2(n_2628),
.Y(n_4296)
);

OAI21x1_ASAP7_75t_SL g4297 ( 
.A1(n_3415),
.A2(n_2627),
.B(n_2807),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_L g4298 ( 
.A(n_3577),
.B(n_3068),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_3577),
.B(n_3068),
.Y(n_4299)
);

AOI221x1_ASAP7_75t_L g4300 ( 
.A1(n_3760),
.A2(n_3358),
.B1(n_3349),
.B2(n_3338),
.C(n_3328),
.Y(n_4300)
);

AOI21xp5_ASAP7_75t_L g4301 ( 
.A1(n_3779),
.A2(n_2767),
.B(n_2750),
.Y(n_4301)
);

BUFx2_ASAP7_75t_L g4302 ( 
.A(n_3405),
.Y(n_4302)
);

OAI21xp5_ASAP7_75t_L g4303 ( 
.A1(n_3473),
.A2(n_2812),
.B(n_2813),
.Y(n_4303)
);

OAI21xp5_ASAP7_75t_L g4304 ( 
.A1(n_3473),
.A2(n_2812),
.B(n_2813),
.Y(n_4304)
);

INVx1_ASAP7_75t_L g4305 ( 
.A(n_3663),
.Y(n_4305)
);

HB1xp67_ASAP7_75t_L g4306 ( 
.A(n_3915),
.Y(n_4306)
);

AOI21xp5_ASAP7_75t_L g4307 ( 
.A1(n_3666),
.A2(n_2767),
.B(n_2748),
.Y(n_4307)
);

OAI21x1_ASAP7_75t_SL g4308 ( 
.A1(n_3415),
.A2(n_3605),
.B(n_3824),
.Y(n_4308)
);

AOI21xp5_ASAP7_75t_L g4309 ( 
.A1(n_3666),
.A2(n_2767),
.B(n_2748),
.Y(n_4309)
);

OAI21x1_ASAP7_75t_L g4310 ( 
.A1(n_3690),
.A2(n_2723),
.B(n_2650),
.Y(n_4310)
);

BUFx10_ASAP7_75t_L g4311 ( 
.A(n_3428),
.Y(n_4311)
);

A2O1A1Ixp33_ASAP7_75t_L g4312 ( 
.A1(n_3720),
.A2(n_2274),
.B(n_2277),
.C(n_2288),
.Y(n_4312)
);

A2O1A1Ixp33_ASAP7_75t_L g4313 ( 
.A1(n_3756),
.A2(n_2277),
.B(n_2288),
.C(n_2317),
.Y(n_4313)
);

OAI21x1_ASAP7_75t_L g4314 ( 
.A1(n_3606),
.A2(n_2663),
.B(n_2650),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3663),
.Y(n_4315)
);

O2A1O1Ixp33_ASAP7_75t_L g4316 ( 
.A1(n_3717),
.A2(n_2716),
.B(n_2640),
.C(n_2599),
.Y(n_4316)
);

BUFx6f_ASAP7_75t_L g4317 ( 
.A(n_3686),
.Y(n_4317)
);

A2O1A1Ixp33_ASAP7_75t_L g4318 ( 
.A1(n_3889),
.A2(n_2277),
.B(n_2288),
.C(n_2317),
.Y(n_4318)
);

OAI21xp5_ASAP7_75t_L g4319 ( 
.A1(n_3508),
.A2(n_2368),
.B(n_2716),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_3741),
.B(n_3742),
.Y(n_4320)
);

OAI21xp5_ASAP7_75t_L g4321 ( 
.A1(n_3508),
.A2(n_2368),
.B(n_2716),
.Y(n_4321)
);

OAI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_3890),
.A2(n_2368),
.B(n_2778),
.Y(n_4322)
);

INVxp67_ASAP7_75t_SL g4323 ( 
.A(n_3692),
.Y(n_4323)
);

AO31x2_ASAP7_75t_L g4324 ( 
.A1(n_3762),
.A2(n_2627),
.A3(n_2796),
.B(n_2709),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_3714),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_3714),
.Y(n_4326)
);

INVx3_ASAP7_75t_L g4327 ( 
.A(n_3700),
.Y(n_4327)
);

NAND2xp5_ASAP7_75t_L g4328 ( 
.A(n_3741),
.B(n_3068),
.Y(n_4328)
);

OAI22xp33_ASAP7_75t_L g4329 ( 
.A1(n_3817),
.A2(n_2288),
.B1(n_2317),
.B2(n_2322),
.Y(n_4329)
);

AO31x2_ASAP7_75t_L g4330 ( 
.A1(n_3762),
.A2(n_2627),
.A3(n_2796),
.B(n_2739),
.Y(n_4330)
);

AOI21xp5_ASAP7_75t_L g4331 ( 
.A1(n_3548),
.A2(n_2748),
.B(n_2767),
.Y(n_4331)
);

AND2x2_ASAP7_75t_L g4332 ( 
.A(n_3561),
.B(n_3068),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_3718),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_3548),
.A2(n_2767),
.B(n_2750),
.Y(n_4334)
);

AOI21xp5_ASAP7_75t_L g4335 ( 
.A1(n_3549),
.A2(n_3550),
.B(n_3759),
.Y(n_4335)
);

NAND2x1p5_ASAP7_75t_L g4336 ( 
.A(n_3679),
.B(n_2748),
.Y(n_4336)
);

AO31x2_ASAP7_75t_L g4337 ( 
.A1(n_3857),
.A2(n_2723),
.A3(n_2796),
.B(n_2621),
.Y(n_4337)
);

AOI22xp33_ASAP7_75t_SL g4338 ( 
.A1(n_3864),
.A2(n_2317),
.B1(n_2322),
.B2(n_2398),
.Y(n_4338)
);

BUFx2_ASAP7_75t_L g4339 ( 
.A(n_3405),
.Y(n_4339)
);

BUFx10_ASAP7_75t_L g4340 ( 
.A(n_3428),
.Y(n_4340)
);

NAND2xp5_ASAP7_75t_SL g4341 ( 
.A(n_3581),
.B(n_3131),
.Y(n_4341)
);

INVx3_ASAP7_75t_SL g4342 ( 
.A(n_3852),
.Y(n_4342)
);

NAND2xp5_ASAP7_75t_L g4343 ( 
.A(n_3742),
.B(n_3131),
.Y(n_4343)
);

INVx1_ASAP7_75t_L g4344 ( 
.A(n_3718),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3625),
.B(n_3131),
.Y(n_4345)
);

NOR2xp33_ASAP7_75t_L g4346 ( 
.A(n_3582),
.B(n_3131),
.Y(n_4346)
);

AOI21x1_ASAP7_75t_SL g4347 ( 
.A1(n_3482),
.A2(n_2797),
.B(n_2368),
.Y(n_4347)
);

BUFx3_ASAP7_75t_L g4348 ( 
.A(n_3686),
.Y(n_4348)
);

AOI21xp5_ASAP7_75t_L g4349 ( 
.A1(n_3549),
.A2(n_2748),
.B(n_2750),
.Y(n_4349)
);

NAND2xp33_ASAP7_75t_SL g4350 ( 
.A(n_3670),
.B(n_3131),
.Y(n_4350)
);

OAI21x1_ASAP7_75t_L g4351 ( 
.A1(n_3430),
.A2(n_2621),
.B(n_2663),
.Y(n_4351)
);

AOI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_3856),
.A2(n_2368),
.B1(n_2498),
.B2(n_2594),
.Y(n_4352)
);

OAI21x1_ASAP7_75t_L g4353 ( 
.A1(n_3430),
.A2(n_2621),
.B(n_2663),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_3776),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_3550),
.A2(n_2767),
.B(n_2750),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3776),
.Y(n_4356)
);

BUFx2_ASAP7_75t_R g4357 ( 
.A(n_3723),
.Y(n_4357)
);

INVx1_ASAP7_75t_L g4358 ( 
.A(n_3789),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_3789),
.Y(n_4359)
);

AOI21x1_ASAP7_75t_L g4360 ( 
.A1(n_3716),
.A2(n_2788),
.B(n_2490),
.Y(n_4360)
);

A2O1A1Ixp33_ASAP7_75t_L g4361 ( 
.A1(n_3889),
.A2(n_2322),
.B(n_2398),
.C(n_2334),
.Y(n_4361)
);

OAI22xp33_ASAP7_75t_L g4362 ( 
.A1(n_3817),
.A2(n_2322),
.B1(n_2398),
.B2(n_2334),
.Y(n_4362)
);

AOI21xp5_ASAP7_75t_L g4363 ( 
.A1(n_3613),
.A2(n_2750),
.B(n_2595),
.Y(n_4363)
);

BUFx10_ASAP7_75t_L g4364 ( 
.A(n_3428),
.Y(n_4364)
);

NOR2xp67_ASAP7_75t_L g4365 ( 
.A(n_3406),
.B(n_3134),
.Y(n_4365)
);

OAI21xp5_ASAP7_75t_L g4366 ( 
.A1(n_3890),
.A2(n_2368),
.B(n_2788),
.Y(n_4366)
);

AOI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_3750),
.A2(n_2750),
.B(n_2595),
.Y(n_4367)
);

AOI21xp5_ASAP7_75t_L g4368 ( 
.A1(n_3750),
.A2(n_2750),
.B(n_2595),
.Y(n_4368)
);

AOI221x1_ASAP7_75t_L g4369 ( 
.A1(n_3717),
.A2(n_3358),
.B1(n_3349),
.B2(n_3338),
.C(n_3328),
.Y(n_4369)
);

CKINVDCx5p33_ASAP7_75t_R g4370 ( 
.A(n_3682),
.Y(n_4370)
);

INVx1_ASAP7_75t_SL g4371 ( 
.A(n_3765),
.Y(n_4371)
);

BUFx3_ASAP7_75t_L g4372 ( 
.A(n_3405),
.Y(n_4372)
);

OAI22xp5_ASAP7_75t_L g4373 ( 
.A1(n_3581),
.A2(n_3455),
.B1(n_3626),
.B2(n_3856),
.Y(n_4373)
);

OAI21xp5_ASAP7_75t_L g4374 ( 
.A1(n_3397),
.A2(n_2368),
.B(n_2334),
.Y(n_4374)
);

A2O1A1Ixp33_ASAP7_75t_L g4375 ( 
.A1(n_3466),
.A2(n_2360),
.B(n_2345),
.C(n_2358),
.Y(n_4375)
);

A2O1A1Ixp33_ASAP7_75t_L g4376 ( 
.A1(n_3466),
.A2(n_2360),
.B(n_2345),
.C(n_2358),
.Y(n_4376)
);

O2A1O1Ixp33_ASAP7_75t_SL g4377 ( 
.A1(n_3618),
.A2(n_2797),
.B(n_2368),
.C(n_2786),
.Y(n_4377)
);

AOI21xp5_ASAP7_75t_L g4378 ( 
.A1(n_3768),
.A2(n_2333),
.B(n_2542),
.Y(n_4378)
);

OAI21xp5_ASAP7_75t_L g4379 ( 
.A1(n_3397),
.A2(n_2360),
.B(n_2345),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_SL g4380 ( 
.A(n_3600),
.B(n_3134),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_3625),
.B(n_3134),
.Y(n_4381)
);

NOR2xp33_ASAP7_75t_SL g4382 ( 
.A(n_3582),
.B(n_2797),
.Y(n_4382)
);

BUFx3_ASAP7_75t_L g4383 ( 
.A(n_3425),
.Y(n_4383)
);

NOR2xp33_ASAP7_75t_L g4384 ( 
.A(n_3919),
.B(n_3134),
.Y(n_4384)
);

INVx5_ASAP7_75t_L g4385 ( 
.A(n_3445),
.Y(n_4385)
);

OAI21xp5_ASAP7_75t_L g4386 ( 
.A1(n_3468),
.A2(n_2360),
.B(n_2345),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_SL g4387 ( 
.A(n_3659),
.B(n_3134),
.Y(n_4387)
);

BUFx4_ASAP7_75t_SL g4388 ( 
.A(n_3723),
.Y(n_4388)
);

BUFx10_ASAP7_75t_L g4389 ( 
.A(n_3445),
.Y(n_4389)
);

NAND3xp33_ASAP7_75t_L g4390 ( 
.A(n_3468),
.B(n_3437),
.C(n_3944),
.Y(n_4390)
);

NAND2xp5_ASAP7_75t_L g4391 ( 
.A(n_3829),
.B(n_3241),
.Y(n_4391)
);

O2A1O1Ixp33_ASAP7_75t_L g4392 ( 
.A1(n_3453),
.A2(n_2640),
.B(n_2358),
.C(n_2359),
.Y(n_4392)
);

OAI22x1_ASAP7_75t_L g4393 ( 
.A1(n_3539),
.A2(n_2621),
.B1(n_2786),
.B2(n_2780),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_3768),
.A2(n_2333),
.B(n_2542),
.Y(n_4394)
);

BUFx6f_ASAP7_75t_L g4395 ( 
.A(n_3723),
.Y(n_4395)
);

AOI21xp5_ASAP7_75t_L g4396 ( 
.A1(n_3653),
.A2(n_2333),
.B(n_2542),
.Y(n_4396)
);

AND2x4_ASAP7_75t_L g4397 ( 
.A(n_3875),
.B(n_3241),
.Y(n_4397)
);

AOI22xp33_ASAP7_75t_L g4398 ( 
.A1(n_3437),
.A2(n_2498),
.B1(n_2594),
.B2(n_2413),
.Y(n_4398)
);

O2A1O1Ixp33_ASAP7_75t_L g4399 ( 
.A1(n_3453),
.A2(n_2640),
.B(n_2358),
.C(n_2359),
.Y(n_4399)
);

AO31x2_ASAP7_75t_L g4400 ( 
.A1(n_3857),
.A2(n_2630),
.A3(n_2786),
.B(n_2780),
.Y(n_4400)
);

NOR2xp67_ASAP7_75t_L g4401 ( 
.A(n_3406),
.B(n_3358),
.Y(n_4401)
);

INVx4_ASAP7_75t_L g4402 ( 
.A(n_3740),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_3704),
.A2(n_2498),
.B1(n_2594),
.B2(n_2413),
.Y(n_4403)
);

NOR2xp33_ASAP7_75t_L g4404 ( 
.A(n_3682),
.B(n_3358),
.Y(n_4404)
);

INVx1_ASAP7_75t_SL g4405 ( 
.A(n_3765),
.Y(n_4405)
);

BUFx12f_ASAP7_75t_L g4406 ( 
.A(n_3682),
.Y(n_4406)
);

A2O1A1Ixp33_ASAP7_75t_L g4407 ( 
.A1(n_3810),
.A2(n_2398),
.B(n_2359),
.C(n_2369),
.Y(n_4407)
);

OAI22xp33_ASAP7_75t_L g4408 ( 
.A1(n_3486),
.A2(n_2369),
.B1(n_2359),
.B2(n_3358),
.Y(n_4408)
);

INVxp67_ASAP7_75t_SL g4409 ( 
.A(n_3665),
.Y(n_4409)
);

OAI21x1_ASAP7_75t_L g4410 ( 
.A1(n_3754),
.A2(n_3773),
.B(n_3446),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_SL g4411 ( 
.A(n_3659),
.B(n_3349),
.Y(n_4411)
);

AOI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_3653),
.A2(n_2333),
.B(n_2528),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_3829),
.B(n_3349),
.Y(n_4413)
);

OAI22x1_ASAP7_75t_L g4414 ( 
.A1(n_3602),
.A2(n_2619),
.B1(n_2786),
.B2(n_2613),
.Y(n_4414)
);

NOR2xp33_ASAP7_75t_SL g4415 ( 
.A(n_3680),
.B(n_2797),
.Y(n_4415)
);

INVx2_ASAP7_75t_SL g4416 ( 
.A(n_3700),
.Y(n_4416)
);

OAI21x1_ASAP7_75t_L g4417 ( 
.A1(n_3431),
.A2(n_2619),
.B(n_2706),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_3561),
.B(n_3349),
.Y(n_4418)
);

OAI21x1_ASAP7_75t_L g4419 ( 
.A1(n_3431),
.A2(n_2613),
.B(n_2706),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_3802),
.Y(n_4420)
);

BUFx2_ASAP7_75t_L g4421 ( 
.A(n_3425),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_3802),
.Y(n_4422)
);

AOI21xp5_ASAP7_75t_L g4423 ( 
.A1(n_3676),
.A2(n_2333),
.B(n_2542),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_L g4424 ( 
.A(n_3830),
.B(n_3338),
.Y(n_4424)
);

BUFx6f_ASAP7_75t_L g4425 ( 
.A(n_3740),
.Y(n_4425)
);

INVx2_ASAP7_75t_SL g4426 ( 
.A(n_3700),
.Y(n_4426)
);

AOI22xp33_ASAP7_75t_L g4427 ( 
.A1(n_3704),
.A2(n_2413),
.B1(n_2594),
.B2(n_2498),
.Y(n_4427)
);

AOI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_3885),
.A2(n_2413),
.B1(n_2594),
.B2(n_2498),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_3830),
.B(n_3338),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_3940),
.Y(n_4430)
);

INVx1_ASAP7_75t_L g4431 ( 
.A(n_3827),
.Y(n_4431)
);

O2A1O1Ixp33_ASAP7_75t_SL g4432 ( 
.A1(n_3794),
.A2(n_2513),
.B(n_2600),
.C(n_2611),
.Y(n_4432)
);

OAI21xp5_ASAP7_75t_L g4433 ( 
.A1(n_3595),
.A2(n_2369),
.B(n_2594),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_3393),
.B(n_3338),
.Y(n_4434)
);

OAI21x1_ASAP7_75t_L g4435 ( 
.A1(n_3446),
.A2(n_2743),
.B(n_2709),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_3426),
.B(n_3328),
.Y(n_4436)
);

AO31x2_ASAP7_75t_L g4437 ( 
.A1(n_3766),
.A2(n_2613),
.A3(n_2780),
.B(n_2777),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_SL g4438 ( 
.A(n_3736),
.B(n_3241),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_3426),
.B(n_3328),
.Y(n_4439)
);

AO31x2_ASAP7_75t_L g4440 ( 
.A1(n_3767),
.A2(n_2611),
.A3(n_2777),
.B(n_2769),
.Y(n_4440)
);

INVx1_ASAP7_75t_L g4441 ( 
.A(n_3827),
.Y(n_4441)
);

O2A1O1Ixp33_ASAP7_75t_SL g4442 ( 
.A1(n_3796),
.A2(n_2611),
.B(n_2777),
.C(n_2769),
.Y(n_4442)
);

OAI22xp5_ASAP7_75t_L g4443 ( 
.A1(n_3455),
.A2(n_2640),
.B1(n_2729),
.B2(n_2389),
.Y(n_4443)
);

AOI221x1_ASAP7_75t_L g4444 ( 
.A1(n_3677),
.A2(n_3328),
.B1(n_3241),
.B2(n_3264),
.C(n_2711),
.Y(n_4444)
);

AO31x2_ASAP7_75t_L g4445 ( 
.A1(n_3767),
.A2(n_2605),
.A3(n_2777),
.B(n_2769),
.Y(n_4445)
);

OAI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_3595),
.A2(n_2594),
.B(n_2498),
.Y(n_4446)
);

BUFx2_ASAP7_75t_L g4447 ( 
.A(n_3425),
.Y(n_4447)
);

CKINVDCx11_ASAP7_75t_R g4448 ( 
.A(n_3740),
.Y(n_4448)
);

AND2x2_ASAP7_75t_SL g4449 ( 
.A(n_3640),
.B(n_3264),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_3813),
.B(n_3264),
.Y(n_4450)
);

AO31x2_ASAP7_75t_L g4451 ( 
.A1(n_3780),
.A2(n_2605),
.A3(n_2769),
.B(n_2743),
.Y(n_4451)
);

AOI21xp5_ASAP7_75t_L g4452 ( 
.A1(n_3676),
.A2(n_2380),
.B(n_2528),
.Y(n_4452)
);

OAI21x1_ASAP7_75t_L g4453 ( 
.A1(n_3451),
.A2(n_2600),
.B(n_2575),
.Y(n_4453)
);

AO22x2_ASAP7_75t_L g4454 ( 
.A1(n_3834),
.A2(n_2600),
.B1(n_2743),
.B2(n_2739),
.Y(n_4454)
);

OAI21x1_ASAP7_75t_L g4455 ( 
.A1(n_3451),
.A2(n_2600),
.B(n_2575),
.Y(n_4455)
);

AOI221x1_ASAP7_75t_L g4456 ( 
.A1(n_3677),
.A2(n_3264),
.B1(n_3241),
.B2(n_2708),
.C(n_2501),
.Y(n_4456)
);

BUFx2_ASAP7_75t_R g4457 ( 
.A(n_3654),
.Y(n_4457)
);

O2A1O1Ixp5_ASAP7_75t_L g4458 ( 
.A1(n_3568),
.A2(n_2743),
.B(n_2739),
.C(n_2723),
.Y(n_4458)
);

OAI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_3417),
.A2(n_3524),
.B(n_3850),
.Y(n_4459)
);

AO31x2_ASAP7_75t_L g4460 ( 
.A1(n_3780),
.A2(n_2563),
.A3(n_2706),
.B(n_2739),
.Y(n_4460)
);

OAI21x1_ASAP7_75t_L g4461 ( 
.A1(n_3452),
.A2(n_2699),
.B(n_2563),
.Y(n_4461)
);

BUFx2_ASAP7_75t_L g4462 ( 
.A(n_3425),
.Y(n_4462)
);

NOR2xp67_ASAP7_75t_L g4463 ( 
.A(n_3406),
.B(n_3264),
.Y(n_4463)
);

O2A1O1Ixp5_ASAP7_75t_L g4464 ( 
.A1(n_3568),
.A2(n_2575),
.B(n_2706),
.C(n_2699),
.Y(n_4464)
);

AOI21xp5_ASAP7_75t_L g4465 ( 
.A1(n_3826),
.A2(n_2380),
.B(n_2628),
.Y(n_4465)
);

OAI22xp5_ASAP7_75t_L g4466 ( 
.A1(n_3904),
.A2(n_3486),
.B1(n_3521),
.B2(n_3885),
.Y(n_4466)
);

INVx1_ASAP7_75t_L g4467 ( 
.A(n_3873),
.Y(n_4467)
);

OAI21x1_ASAP7_75t_L g4468 ( 
.A1(n_3452),
.A2(n_2563),
.B(n_2636),
.Y(n_4468)
);

OA21x2_ASAP7_75t_L g4469 ( 
.A1(n_3944),
.A2(n_2575),
.B(n_2636),
.Y(n_4469)
);

AOI21xp5_ASAP7_75t_L g4470 ( 
.A1(n_3826),
.A2(n_2380),
.B(n_2628),
.Y(n_4470)
);

NAND2xp5_ASAP7_75t_L g4471 ( 
.A(n_3813),
.B(n_2642),
.Y(n_4471)
);

A2O1A1Ixp33_ASAP7_75t_L g4472 ( 
.A1(n_3810),
.A2(n_2389),
.B(n_2729),
.C(n_2536),
.Y(n_4472)
);

BUFx3_ASAP7_75t_L g4473 ( 
.A(n_3425),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_3821),
.B(n_2642),
.Y(n_4474)
);

CKINVDCx6p67_ASAP7_75t_R g4475 ( 
.A(n_3682),
.Y(n_4475)
);

OAI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_3417),
.A2(n_2594),
.B(n_2498),
.Y(n_4476)
);

NOR2xp33_ASAP7_75t_L g4477 ( 
.A(n_3881),
.B(n_2389),
.Y(n_4477)
);

AOI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_3644),
.A2(n_2380),
.B(n_2628),
.Y(n_4478)
);

CKINVDCx5p33_ASAP7_75t_R g4479 ( 
.A(n_3772),
.Y(n_4479)
);

A2O1A1Ixp33_ASAP7_75t_L g4480 ( 
.A1(n_3524),
.A2(n_2389),
.B(n_2729),
.C(n_2724),
.Y(n_4480)
);

INVx2_ASAP7_75t_SL g4481 ( 
.A(n_3733),
.Y(n_4481)
);

AOI22xp5_ASAP7_75t_L g4482 ( 
.A1(n_3882),
.A2(n_2594),
.B1(n_2413),
.B2(n_2498),
.Y(n_4482)
);

OAI21x1_ASAP7_75t_L g4483 ( 
.A1(n_3649),
.A2(n_2490),
.B(n_2513),
.Y(n_4483)
);

AOI21xp5_ASAP7_75t_L g4484 ( 
.A1(n_3644),
.A2(n_2628),
.B(n_2595),
.Y(n_4484)
);

INVx2_ASAP7_75t_SL g4485 ( 
.A(n_3733),
.Y(n_4485)
);

INVx2_ASAP7_75t_L g4486 ( 
.A(n_3630),
.Y(n_4486)
);

INVx4_ASAP7_75t_L g4487 ( 
.A(n_3795),
.Y(n_4487)
);

CKINVDCx5p33_ASAP7_75t_R g4488 ( 
.A(n_3491),
.Y(n_4488)
);

OAI22xp5_ASAP7_75t_L g4489 ( 
.A1(n_3904),
.A2(n_2729),
.B1(n_2389),
.B2(n_2551),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_3821),
.B(n_2642),
.Y(n_4490)
);

O2A1O1Ixp33_ASAP7_75t_L g4491 ( 
.A1(n_3489),
.A2(n_2490),
.B(n_2513),
.C(n_2605),
.Y(n_4491)
);

A2O1A1Ixp33_ASAP7_75t_L g4492 ( 
.A1(n_3521),
.A2(n_2389),
.B(n_2729),
.C(n_2551),
.Y(n_4492)
);

AO31x2_ASAP7_75t_L g4493 ( 
.A1(n_3913),
.A2(n_2490),
.A3(n_2526),
.B(n_2513),
.Y(n_4493)
);

OAI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_3850),
.A2(n_2594),
.B(n_2413),
.Y(n_4494)
);

OAI21xp5_ASAP7_75t_L g4495 ( 
.A1(n_3917),
.A2(n_2413),
.B(n_2498),
.Y(n_4495)
);

OAI22xp33_ASAP7_75t_L g4496 ( 
.A1(n_3818),
.A2(n_2389),
.B1(n_2729),
.B2(n_2549),
.Y(n_4496)
);

O2A1O1Ixp33_ASAP7_75t_L g4497 ( 
.A1(n_3489),
.A2(n_2526),
.B(n_2494),
.C(n_2636),
.Y(n_4497)
);

CKINVDCx11_ASAP7_75t_R g4498 ( 
.A(n_3733),
.Y(n_4498)
);

AOI221xp5_ASAP7_75t_L g4499 ( 
.A1(n_3793),
.A2(n_2389),
.B1(n_2729),
.B2(n_2650),
.C(n_2636),
.Y(n_4499)
);

INVx1_ASAP7_75t_L g4500 ( 
.A(n_3873),
.Y(n_4500)
);

AO31x2_ASAP7_75t_L g4501 ( 
.A1(n_3913),
.A2(n_2526),
.A3(n_2494),
.B(n_2650),
.Y(n_4501)
);

A2O1A1Ixp33_ASAP7_75t_L g4502 ( 
.A1(n_3738),
.A2(n_2389),
.B(n_2729),
.C(n_2540),
.Y(n_4502)
);

OAI21xp5_ASAP7_75t_L g4503 ( 
.A1(n_3917),
.A2(n_2413),
.B(n_2498),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3798),
.B(n_2642),
.Y(n_4504)
);

OAI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_3882),
.A2(n_2549),
.B1(n_2708),
.B2(n_2438),
.Y(n_4505)
);

AOI221xp5_ASAP7_75t_L g4506 ( 
.A1(n_3793),
.A2(n_2526),
.B1(n_2494),
.B2(n_2438),
.C(n_2464),
.Y(n_4506)
);

BUFx3_ASAP7_75t_L g4507 ( 
.A(n_3425),
.Y(n_4507)
);

OR2x2_ASAP7_75t_L g4508 ( 
.A(n_3940),
.B(n_2494),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_L g4509 ( 
.A(n_3798),
.B(n_2642),
.Y(n_4509)
);

OAI22x1_ASAP7_75t_L g4510 ( 
.A1(n_3763),
.A2(n_2419),
.B1(n_2528),
.B2(n_2642),
.Y(n_4510)
);

OAI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_3429),
.A2(n_2413),
.B(n_2810),
.Y(n_4511)
);

OAI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_3661),
.A2(n_2413),
.B(n_2810),
.Y(n_4512)
);

NAND2xp5_ASAP7_75t_L g4513 ( 
.A(n_3876),
.B(n_2642),
.Y(n_4513)
);

AOI21xp5_ASAP7_75t_L g4514 ( 
.A1(n_3661),
.A2(n_2419),
.B(n_2528),
.Y(n_4514)
);

AND2x4_ASAP7_75t_L g4515 ( 
.A(n_3875),
.B(n_2551),
.Y(n_4515)
);

AOI221x1_ASAP7_75t_L g4516 ( 
.A1(n_3731),
.A2(n_3500),
.B1(n_3558),
.B2(n_3449),
.C(n_3579),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_3876),
.B(n_2642),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_3877),
.B(n_2642),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_3877),
.B(n_2642),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_SL g4520 ( 
.A(n_3406),
.B(n_2721),
.Y(n_4520)
);

OAI21x1_ASAP7_75t_L g4521 ( 
.A1(n_4410),
.A2(n_3449),
.B(n_3825),
.Y(n_4521)
);

BUFx2_ASAP7_75t_L g4522 ( 
.A(n_4372),
.Y(n_4522)
);

OAI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_3966),
.A2(n_3579),
.B(n_3846),
.Y(n_4523)
);

INVx2_ASAP7_75t_L g4524 ( 
.A(n_3953),
.Y(n_4524)
);

INVx1_ASAP7_75t_L g4525 ( 
.A(n_3951),
.Y(n_4525)
);

OAI21xp5_ASAP7_75t_L g4526 ( 
.A1(n_3966),
.A2(n_3818),
.B(n_3555),
.Y(n_4526)
);

OAI22xp33_ASAP7_75t_L g4527 ( 
.A1(n_4031),
.A2(n_3818),
.B1(n_3713),
.B2(n_3899),
.Y(n_4527)
);

CKINVDCx16_ASAP7_75t_R g4528 ( 
.A(n_4081),
.Y(n_4528)
);

OA21x2_ASAP7_75t_L g4529 ( 
.A1(n_4410),
.A2(n_3910),
.B(n_3896),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_3945),
.B(n_3863),
.Y(n_4530)
);

INVx2_ASAP7_75t_SL g4531 ( 
.A(n_4385),
.Y(n_4531)
);

INVx3_ASAP7_75t_L g4532 ( 
.A(n_4372),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4335),
.B(n_4118),
.Y(n_4533)
);

INVx8_ASAP7_75t_L g4534 ( 
.A(n_4406),
.Y(n_4534)
);

INVx2_ASAP7_75t_R g4535 ( 
.A(n_4385),
.Y(n_4535)
);

AO31x2_ASAP7_75t_L g4536 ( 
.A1(n_4516),
.A2(n_3536),
.A3(n_3910),
.B(n_3843),
.Y(n_4536)
);

OAI21xp5_ASAP7_75t_L g4537 ( 
.A1(n_3969),
.A2(n_3555),
.B(n_3528),
.Y(n_4537)
);

BUFx3_ASAP7_75t_L g4538 ( 
.A(n_4406),
.Y(n_4538)
);

OAI22xp5_ASAP7_75t_L g4539 ( 
.A1(n_4466),
.A2(n_3738),
.B1(n_3930),
.B2(n_3926),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_3947),
.B(n_3558),
.Y(n_4540)
);

INVx5_ASAP7_75t_L g4541 ( 
.A(n_4221),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_3951),
.Y(n_4542)
);

AOI22xp5_ASAP7_75t_L g4543 ( 
.A1(n_4218),
.A2(n_3864),
.B1(n_3558),
.B2(n_3899),
.Y(n_4543)
);

AOI22xp33_ASAP7_75t_SL g4544 ( 
.A1(n_3952),
.A2(n_3864),
.B1(n_3879),
.B2(n_3558),
.Y(n_4544)
);

AO32x2_ASAP7_75t_L g4545 ( 
.A1(n_4416),
.A2(n_3589),
.A3(n_3658),
.B1(n_3498),
.B2(n_3491),
.Y(n_4545)
);

BUFx2_ASAP7_75t_SL g4546 ( 
.A(n_4385),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_L g4547 ( 
.A(n_4084),
.B(n_3424),
.Y(n_4547)
);

OA21x2_ASAP7_75t_L g4548 ( 
.A1(n_4516),
.A2(n_3921),
.B(n_3734),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_3956),
.Y(n_4549)
);

OAI22xp5_ASAP7_75t_L g4550 ( 
.A1(n_4390),
.A2(n_3926),
.B1(n_3930),
.B2(n_3558),
.Y(n_4550)
);

OAI21xp5_ASAP7_75t_L g4551 ( 
.A1(n_4390),
.A2(n_3528),
.B(n_3562),
.Y(n_4551)
);

AOI21xp33_ASAP7_75t_L g4552 ( 
.A1(n_4211),
.A2(n_3500),
.B(n_3930),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_3947),
.B(n_3424),
.Y(n_4553)
);

AOI22xp33_ASAP7_75t_L g4554 ( 
.A1(n_4218),
.A2(n_3852),
.B1(n_3713),
.B2(n_3506),
.Y(n_4554)
);

OR2x6_ASAP7_75t_L g4555 ( 
.A(n_4167),
.B(n_3556),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4084),
.B(n_3424),
.Y(n_4556)
);

CKINVDCx5p33_ASAP7_75t_R g4557 ( 
.A(n_3998),
.Y(n_4557)
);

AND2x4_ASAP7_75t_L g4558 ( 
.A(n_4473),
.B(n_3406),
.Y(n_4558)
);

OAI21x1_ASAP7_75t_L g4559 ( 
.A1(n_4203),
.A2(n_3464),
.B(n_3458),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4026),
.B(n_3863),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4026),
.B(n_3540),
.Y(n_4561)
);

OAI22xp5_ASAP7_75t_L g4562 ( 
.A1(n_3952),
.A2(n_3454),
.B1(n_3540),
.B2(n_3634),
.Y(n_4562)
);

AND2x4_ASAP7_75t_L g4563 ( 
.A(n_4383),
.B(n_3406),
.Y(n_4563)
);

OAI21x1_ASAP7_75t_L g4564 ( 
.A1(n_4203),
.A2(n_4205),
.B(n_3994),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_3956),
.Y(n_4565)
);

BUFx12f_ASAP7_75t_L g4566 ( 
.A(n_3986),
.Y(n_4566)
);

OAI22xp5_ASAP7_75t_L g4567 ( 
.A1(n_3948),
.A2(n_3454),
.B1(n_3634),
.B2(n_3893),
.Y(n_4567)
);

INVx6_ASAP7_75t_L g4568 ( 
.A(n_4270),
.Y(n_4568)
);

OAI21x1_ASAP7_75t_L g4569 ( 
.A1(n_4205),
.A2(n_3458),
.B(n_3820),
.Y(n_4569)
);

AND2x2_ASAP7_75t_L g4570 ( 
.A(n_4210),
.B(n_3758),
.Y(n_4570)
);

A2O1A1Ixp33_ASAP7_75t_L g4571 ( 
.A1(n_3949),
.A2(n_3669),
.B(n_3788),
.C(n_3633),
.Y(n_4571)
);

AOI221x1_ASAP7_75t_L g4572 ( 
.A1(n_3948),
.A2(n_4167),
.B1(n_4027),
.B2(n_4045),
.C(n_4174),
.Y(n_4572)
);

AOI22xp33_ASAP7_75t_L g4573 ( 
.A1(n_4078),
.A2(n_3852),
.B1(n_3713),
.B2(n_3506),
.Y(n_4573)
);

BUFx2_ASAP7_75t_R g4574 ( 
.A(n_3984),
.Y(n_4574)
);

OR2x2_ASAP7_75t_L g4575 ( 
.A(n_4244),
.B(n_4023),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_3978),
.Y(n_4576)
);

AOI22xp33_ASAP7_75t_L g4577 ( 
.A1(n_4078),
.A2(n_3852),
.B1(n_3713),
.B2(n_3506),
.Y(n_4577)
);

CKINVDCx20_ASAP7_75t_R g4578 ( 
.A(n_3984),
.Y(n_4578)
);

O2A1O1Ixp33_ASAP7_75t_L g4579 ( 
.A1(n_4373),
.A2(n_3562),
.B(n_3560),
.C(n_3731),
.Y(n_4579)
);

NOR2xp33_ASAP7_75t_L g4580 ( 
.A(n_4084),
.B(n_3424),
.Y(n_4580)
);

OR2x2_ASAP7_75t_L g4581 ( 
.A(n_4244),
.B(n_3398),
.Y(n_4581)
);

O2A1O1Ixp5_ASAP7_75t_L g4582 ( 
.A1(n_4211),
.A2(n_3669),
.B(n_3788),
.C(n_3633),
.Y(n_4582)
);

INVxp67_ASAP7_75t_L g4583 ( 
.A(n_4046),
.Y(n_4583)
);

AOI22xp33_ASAP7_75t_L g4584 ( 
.A1(n_4239),
.A2(n_3852),
.B1(n_3713),
.B2(n_3506),
.Y(n_4584)
);

INVx2_ASAP7_75t_L g4585 ( 
.A(n_3983),
.Y(n_4585)
);

AOI21xp5_ASAP7_75t_L g4586 ( 
.A1(n_4110),
.A2(n_3643),
.B(n_3640),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_3978),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_3980),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4210),
.B(n_3758),
.Y(n_4589)
);

OAI222xp33_ASAP7_75t_L g4590 ( 
.A1(n_4031),
.A2(n_3728),
.B1(n_3527),
.B2(n_3911),
.C1(n_3871),
.C2(n_3822),
.Y(n_4590)
);

CKINVDCx5p33_ASAP7_75t_R g4591 ( 
.A(n_4059),
.Y(n_4591)
);

INVx3_ASAP7_75t_SL g4592 ( 
.A(n_4475),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_3980),
.Y(n_4593)
);

OAI21x1_ASAP7_75t_L g4594 ( 
.A1(n_4232),
.A2(n_3842),
.B(n_3462),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_3999),
.Y(n_4595)
);

NOR3xp33_ASAP7_75t_L g4596 ( 
.A(n_4459),
.B(n_3560),
.C(n_3851),
.Y(n_4596)
);

OAI21x1_ASAP7_75t_SL g4597 ( 
.A1(n_4275),
.A2(n_4126),
.B(n_4178),
.Y(n_4597)
);

OAI22xp5_ASAP7_75t_L g4598 ( 
.A1(n_4502),
.A2(n_3893),
.B1(n_3868),
.B2(n_3643),
.Y(n_4598)
);

INVx1_ASAP7_75t_L g4599 ( 
.A(n_3999),
.Y(n_4599)
);

AND2x4_ASAP7_75t_L g4600 ( 
.A(n_4372),
.B(n_3460),
.Y(n_4600)
);

AO21x2_ASAP7_75t_L g4601 ( 
.A1(n_4183),
.A2(n_3664),
.B(n_3641),
.Y(n_4601)
);

OAI21x1_ASAP7_75t_L g4602 ( 
.A1(n_4050),
.A2(n_4058),
.B(n_3973),
.Y(n_4602)
);

NOR2xp33_ASAP7_75t_L g4603 ( 
.A(n_4194),
.B(n_3479),
.Y(n_4603)
);

AOI22xp33_ASAP7_75t_SL g4604 ( 
.A1(n_4081),
.A2(n_3864),
.B1(n_3879),
.B2(n_3640),
.Y(n_4604)
);

OA21x2_ASAP7_75t_L g4605 ( 
.A1(n_4166),
.A2(n_3914),
.B(n_3814),
.Y(n_4605)
);

NAND2x1_ASAP7_75t_L g4606 ( 
.A(n_4027),
.B(n_4080),
.Y(n_4606)
);

AO31x2_ASAP7_75t_L g4607 ( 
.A1(n_4275),
.A2(n_4178),
.A3(n_4456),
.B(n_4126),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4014),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4014),
.Y(n_4609)
);

INVx2_ASAP7_75t_L g4610 ( 
.A(n_4006),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4071),
.B(n_3836),
.Y(n_4611)
);

BUFx5_ASAP7_75t_L g4612 ( 
.A(n_4383),
.Y(n_4612)
);

INVx2_ASAP7_75t_L g4613 ( 
.A(n_4006),
.Y(n_4613)
);

AOI22xp33_ASAP7_75t_SL g4614 ( 
.A1(n_4415),
.A2(n_3879),
.B1(n_3640),
.B2(n_3643),
.Y(n_4614)
);

NOR2xp33_ASAP7_75t_L g4615 ( 
.A(n_4194),
.B(n_3479),
.Y(n_4615)
);

OR2x2_ASAP7_75t_L g4616 ( 
.A(n_4023),
.B(n_4028),
.Y(n_4616)
);

INVx1_ASAP7_75t_SL g4617 ( 
.A(n_4028),
.Y(n_4617)
);

INVx3_ASAP7_75t_L g4618 ( 
.A(n_4383),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4089),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4089),
.Y(n_4620)
);

INVx6_ASAP7_75t_L g4621 ( 
.A(n_4270),
.Y(n_4621)
);

NOR2xp33_ASAP7_75t_L g4622 ( 
.A(n_4194),
.B(n_3479),
.Y(n_4622)
);

AND2x4_ASAP7_75t_L g4623 ( 
.A(n_4473),
.B(n_3460),
.Y(n_4623)
);

BUFx6f_ASAP7_75t_L g4624 ( 
.A(n_4385),
.Y(n_4624)
);

OAI211xp5_ASAP7_75t_L g4625 ( 
.A1(n_4012),
.A2(n_3790),
.B(n_3868),
.C(n_3831),
.Y(n_4625)
);

CKINVDCx5p33_ASAP7_75t_R g4626 ( 
.A(n_4059),
.Y(n_4626)
);

AND2x2_ASAP7_75t_L g4627 ( 
.A(n_3965),
.B(n_3479),
.Y(n_4627)
);

AOI22xp33_ASAP7_75t_L g4628 ( 
.A1(n_4239),
.A2(n_3531),
.B1(n_3935),
.B2(n_3733),
.Y(n_4628)
);

INVx3_ASAP7_75t_L g4629 ( 
.A(n_4473),
.Y(n_4629)
);

INVx2_ASAP7_75t_L g4630 ( 
.A(n_4066),
.Y(n_4630)
);

O2A1O1Ixp33_ASAP7_75t_L g4631 ( 
.A1(n_4012),
.A2(n_3601),
.B(n_3588),
.C(n_3790),
.Y(n_4631)
);

INVx2_ASAP7_75t_L g4632 ( 
.A(n_4072),
.Y(n_4632)
);

BUFx12f_ASAP7_75t_L g4633 ( 
.A(n_4092),
.Y(n_4633)
);

INVx2_ASAP7_75t_L g4634 ( 
.A(n_4072),
.Y(n_4634)
);

OA21x2_ASAP7_75t_L g4635 ( 
.A1(n_4166),
.A2(n_3905),
.B(n_3934),
.Y(n_4635)
);

BUFx2_ASAP7_75t_SL g4636 ( 
.A(n_4385),
.Y(n_4636)
);

INVx2_ASAP7_75t_SL g4637 ( 
.A(n_4385),
.Y(n_4637)
);

BUFx6f_ASAP7_75t_L g4638 ( 
.A(n_4449),
.Y(n_4638)
);

BUFx3_ASAP7_75t_L g4639 ( 
.A(n_4270),
.Y(n_4639)
);

AND2x4_ASAP7_75t_L g4640 ( 
.A(n_4507),
.B(n_3460),
.Y(n_4640)
);

AND2x4_ASAP7_75t_L g4641 ( 
.A(n_4507),
.B(n_3460),
.Y(n_4641)
);

OAI22xp5_ASAP7_75t_L g4642 ( 
.A1(n_4049),
.A2(n_3643),
.B1(n_3753),
.B2(n_3744),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4090),
.Y(n_4643)
);

BUFx12f_ASAP7_75t_L g4644 ( 
.A(n_4109),
.Y(n_4644)
);

OAI21xp5_ASAP7_75t_L g4645 ( 
.A1(n_4049),
.A2(n_3911),
.B(n_3843),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_4071),
.B(n_3836),
.Y(n_4646)
);

AO21x2_ASAP7_75t_L g4647 ( 
.A1(n_4134),
.A2(n_3664),
.B(n_3641),
.Y(n_4647)
);

NAND3xp33_ASAP7_75t_L g4648 ( 
.A(n_4068),
.B(n_3879),
.C(n_3727),
.Y(n_4648)
);

INVx2_ASAP7_75t_L g4649 ( 
.A(n_4075),
.Y(n_4649)
);

AO32x2_ASAP7_75t_L g4650 ( 
.A1(n_4416),
.A2(n_3498),
.A3(n_3685),
.B1(n_3658),
.B2(n_3589),
.Y(n_4650)
);

OAI21x1_ASAP7_75t_L g4651 ( 
.A1(n_3950),
.A2(n_3859),
.B(n_3934),
.Y(n_4651)
);

OAI21x1_ASAP7_75t_L g4652 ( 
.A1(n_3961),
.A2(n_3941),
.B(n_3937),
.Y(n_4652)
);

AND2x4_ASAP7_75t_L g4653 ( 
.A(n_4507),
.B(n_3460),
.Y(n_4653)
);

AND2x2_ASAP7_75t_SL g4654 ( 
.A(n_4415),
.B(n_3836),
.Y(n_4654)
);

AOI21xp33_ASAP7_75t_SL g4655 ( 
.A1(n_4370),
.A2(n_3838),
.B(n_3808),
.Y(n_4655)
);

INVx4_ASAP7_75t_SL g4656 ( 
.A(n_4196),
.Y(n_4656)
);

AND2x2_ASAP7_75t_L g4657 ( 
.A(n_3965),
.B(n_3604),
.Y(n_4657)
);

AO31x2_ASAP7_75t_L g4658 ( 
.A1(n_4456),
.A2(n_3536),
.A3(n_3413),
.B(n_3444),
.Y(n_4658)
);

O2A1O1Ixp33_ASAP7_75t_SL g4659 ( 
.A1(n_4223),
.A2(n_3928),
.B(n_3920),
.C(n_3823),
.Y(n_4659)
);

AOI21x1_ASAP7_75t_L g4660 ( 
.A1(n_4147),
.A2(n_3906),
.B(n_3884),
.Y(n_4660)
);

INVx1_ASAP7_75t_L g4661 ( 
.A(n_4090),
.Y(n_4661)
);

OAI21x1_ASAP7_75t_L g4662 ( 
.A1(n_3961),
.A2(n_4042),
.B(n_4022),
.Y(n_4662)
);

OAI21x1_ASAP7_75t_SL g4663 ( 
.A1(n_4308),
.A2(n_3665),
.B(n_3828),
.Y(n_4663)
);

AND2x4_ASAP7_75t_L g4664 ( 
.A(n_4076),
.B(n_4462),
.Y(n_4664)
);

OR2x2_ASAP7_75t_L g4665 ( 
.A(n_4371),
.B(n_3398),
.Y(n_4665)
);

AOI22xp33_ASAP7_75t_L g4666 ( 
.A1(n_4241),
.A2(n_3531),
.B1(n_3935),
.B2(n_3733),
.Y(n_4666)
);

INVx2_ASAP7_75t_L g4667 ( 
.A(n_4075),
.Y(n_4667)
);

OAI21x1_ASAP7_75t_L g4668 ( 
.A1(n_4022),
.A2(n_4042),
.B(n_4483),
.Y(n_4668)
);

INVx8_ASAP7_75t_L g4669 ( 
.A(n_4479),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4227),
.B(n_3836),
.Y(n_4670)
);

AND2x2_ASAP7_75t_L g4671 ( 
.A(n_4249),
.B(n_3758),
.Y(n_4671)
);

NOR2xp33_ASAP7_75t_L g4672 ( 
.A(n_4051),
.B(n_3604),
.Y(n_4672)
);

INVx1_ASAP7_75t_L g4673 ( 
.A(n_4098),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4098),
.Y(n_4674)
);

INVx4_ASAP7_75t_SL g4675 ( 
.A(n_4342),
.Y(n_4675)
);

INVx3_ASAP7_75t_L g4676 ( 
.A(n_3997),
.Y(n_4676)
);

BUFx6f_ASAP7_75t_L g4677 ( 
.A(n_4449),
.Y(n_4677)
);

NOR2xp33_ASAP7_75t_L g4678 ( 
.A(n_4245),
.B(n_3604),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4111),
.A2(n_3744),
.B1(n_3778),
.B2(n_3753),
.Y(n_4679)
);

OA21x2_ASAP7_75t_L g4680 ( 
.A1(n_4444),
.A2(n_3941),
.B(n_3937),
.Y(n_4680)
);

AOI22xp33_ASAP7_75t_L g4681 ( 
.A1(n_4241),
.A2(n_3531),
.B1(n_3935),
.B2(n_3733),
.Y(n_4681)
);

OAI22xp33_ASAP7_75t_L g4682 ( 
.A1(n_4142),
.A2(n_3531),
.B1(n_3924),
.B2(n_3460),
.Y(n_4682)
);

AND2x2_ASAP7_75t_L g4683 ( 
.A(n_4249),
.B(n_3758),
.Y(n_4683)
);

INVx1_ASAP7_75t_SL g4684 ( 
.A(n_4371),
.Y(n_4684)
);

AO21x2_ASAP7_75t_L g4685 ( 
.A1(n_4308),
.A2(n_3624),
.B(n_3459),
.Y(n_4685)
);

AOI21xp5_ASAP7_75t_L g4686 ( 
.A1(n_4113),
.A2(n_3531),
.B(n_3523),
.Y(n_4686)
);

NAND2x1p5_ASAP7_75t_L g4687 ( 
.A(n_4080),
.B(n_3460),
.Y(n_4687)
);

CKINVDCx16_ASAP7_75t_R g4688 ( 
.A(n_4382),
.Y(n_4688)
);

A2O1A1Ixp33_ASAP7_75t_L g4689 ( 
.A1(n_4055),
.A2(n_3906),
.B(n_3884),
.C(n_3503),
.Y(n_4689)
);

OAI21x1_ASAP7_75t_L g4690 ( 
.A1(n_4360),
.A2(n_3996),
.B(n_4236),
.Y(n_4690)
);

OAI21x1_ASAP7_75t_L g4691 ( 
.A1(n_3996),
.A2(n_3505),
.B(n_3399),
.Y(n_4691)
);

OR2x2_ASAP7_75t_L g4692 ( 
.A(n_4405),
.B(n_3398),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4101),
.Y(n_4693)
);

OAI22xp33_ASAP7_75t_L g4694 ( 
.A1(n_4142),
.A2(n_3924),
.B1(n_3504),
.B2(n_3530),
.Y(n_4694)
);

A2O1A1Ixp33_ASAP7_75t_L g4695 ( 
.A1(n_4217),
.A2(n_3504),
.B(n_3530),
.C(n_3924),
.Y(n_4695)
);

BUFx2_ASAP7_75t_L g4696 ( 
.A(n_3957),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4101),
.Y(n_4697)
);

INVx1_ASAP7_75t_L g4698 ( 
.A(n_4105),
.Y(n_4698)
);

AO21x2_ASAP7_75t_L g4699 ( 
.A1(n_4459),
.A2(n_3624),
.B(n_3459),
.Y(n_4699)
);

INVx1_ASAP7_75t_L g4700 ( 
.A(n_4105),
.Y(n_4700)
);

INVx1_ASAP7_75t_L g4701 ( 
.A(n_4114),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4114),
.Y(n_4702)
);

INVx2_ASAP7_75t_L g4703 ( 
.A(n_4082),
.Y(n_4703)
);

AND2x2_ASAP7_75t_L g4704 ( 
.A(n_4249),
.B(n_3758),
.Y(n_4704)
);

OR2x2_ASAP7_75t_L g4705 ( 
.A(n_4405),
.B(n_3398),
.Y(n_4705)
);

OAI22xp5_ASAP7_75t_SL g4706 ( 
.A1(n_4338),
.A2(n_3888),
.B1(n_3898),
.B2(n_3727),
.Y(n_4706)
);

AOI21xp5_ASAP7_75t_L g4707 ( 
.A1(n_4133),
.A2(n_4138),
.B(n_4155),
.Y(n_4707)
);

OAI21xp5_ASAP7_75t_L g4708 ( 
.A1(n_4152),
.A2(n_3851),
.B(n_3601),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4227),
.B(n_3888),
.Y(n_4709)
);

OAI22xp5_ASAP7_75t_L g4710 ( 
.A1(n_4111),
.A2(n_3778),
.B1(n_3764),
.B2(n_3761),
.Y(n_4710)
);

NOR2xp67_ASAP7_75t_L g4711 ( 
.A(n_4016),
.B(n_3504),
.Y(n_4711)
);

NAND2x1p5_ASAP7_75t_L g4712 ( 
.A(n_4449),
.B(n_3504),
.Y(n_4712)
);

CKINVDCx20_ASAP7_75t_R g4713 ( 
.A(n_4136),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4087),
.Y(n_4714)
);

AOI21xp5_ASAP7_75t_L g4715 ( 
.A1(n_4162),
.A2(n_3523),
.B(n_3888),
.Y(n_4715)
);

BUFx3_ASAP7_75t_L g4716 ( 
.A(n_4270),
.Y(n_4716)
);

OAI22xp33_ASAP7_75t_L g4717 ( 
.A1(n_4352),
.A2(n_3924),
.B1(n_3504),
.B2(n_3530),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_3965),
.B(n_3604),
.Y(n_4718)
);

AOI22xp33_ASAP7_75t_L g4719 ( 
.A1(n_4476),
.A2(n_3935),
.B1(n_3530),
.B2(n_3504),
.Y(n_4719)
);

OAI211xp5_ASAP7_75t_L g4720 ( 
.A1(n_4011),
.A2(n_3831),
.B(n_3588),
.C(n_3888),
.Y(n_4720)
);

NOR2xp33_ASAP7_75t_L g4721 ( 
.A(n_4276),
.B(n_3855),
.Y(n_4721)
);

AND2x4_ASAP7_75t_L g4722 ( 
.A(n_3957),
.B(n_3504),
.Y(n_4722)
);

AND2x4_ASAP7_75t_L g4723 ( 
.A(n_3975),
.B(n_3530),
.Y(n_4723)
);

INVx2_ASAP7_75t_L g4724 ( 
.A(n_4106),
.Y(n_4724)
);

OAI221xp5_ASAP7_75t_L g4725 ( 
.A1(n_4152),
.A2(n_3867),
.B1(n_3898),
.B2(n_3728),
.C(n_3527),
.Y(n_4725)
);

AOI22xp33_ASAP7_75t_L g4726 ( 
.A1(n_4476),
.A2(n_3530),
.B1(n_3425),
.B2(n_3924),
.Y(n_4726)
);

OAI22xp5_ASAP7_75t_L g4727 ( 
.A1(n_4352),
.A2(n_3764),
.B1(n_3761),
.B2(n_3537),
.Y(n_4727)
);

AND2x2_ASAP7_75t_L g4728 ( 
.A(n_3971),
.B(n_3855),
.Y(n_4728)
);

NOR2xp33_ASAP7_75t_L g4729 ( 
.A(n_4064),
.B(n_3855),
.Y(n_4729)
);

BUFx3_ASAP7_75t_L g4730 ( 
.A(n_3954),
.Y(n_4730)
);

BUFx2_ASAP7_75t_L g4731 ( 
.A(n_3975),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4106),
.Y(n_4732)
);

AOI22xp33_ASAP7_75t_L g4733 ( 
.A1(n_4512),
.A2(n_3530),
.B1(n_3425),
.B2(n_3924),
.Y(n_4733)
);

NOR2xp67_ASAP7_75t_L g4734 ( 
.A(n_4016),
.B(n_4206),
.Y(n_4734)
);

BUFx2_ASAP7_75t_L g4735 ( 
.A(n_4076),
.Y(n_4735)
);

NOR2xp33_ASAP7_75t_L g4736 ( 
.A(n_4047),
.B(n_3855),
.Y(n_4736)
);

INVx1_ASAP7_75t_L g4737 ( 
.A(n_4159),
.Y(n_4737)
);

AO21x2_ASAP7_75t_L g4738 ( 
.A1(n_4279),
.A2(n_4193),
.B(n_4069),
.Y(n_4738)
);

OA21x2_ASAP7_75t_L g4739 ( 
.A1(n_4444),
.A2(n_4300),
.B(n_4168),
.Y(n_4739)
);

AO21x2_ASAP7_75t_L g4740 ( 
.A1(n_4062),
.A2(n_3624),
.B(n_3459),
.Y(n_4740)
);

AO21x2_ASAP7_75t_L g4741 ( 
.A1(n_4184),
.A2(n_3624),
.B(n_3459),
.Y(n_4741)
);

BUFx8_ASAP7_75t_SL g4742 ( 
.A(n_4188),
.Y(n_4742)
);

A2O1A1Ixp33_ASAP7_75t_L g4743 ( 
.A1(n_4179),
.A2(n_3924),
.B(n_3844),
.C(n_3927),
.Y(n_4743)
);

CKINVDCx5p33_ASAP7_75t_R g4744 ( 
.A(n_4188),
.Y(n_4744)
);

OAI21xp5_ASAP7_75t_L g4745 ( 
.A1(n_3962),
.A2(n_3698),
.B(n_3642),
.Y(n_4745)
);

NOR2xp67_ASAP7_75t_L g4746 ( 
.A(n_4331),
.B(n_3413),
.Y(n_4746)
);

INVx3_ASAP7_75t_L g4747 ( 
.A(n_3997),
.Y(n_4747)
);

AOI22xp33_ASAP7_75t_L g4748 ( 
.A1(n_4512),
.A2(n_3927),
.B1(n_3801),
.B2(n_3844),
.Y(n_4748)
);

NOR2xp33_ASAP7_75t_SL g4749 ( 
.A(n_4357),
.B(n_3795),
.Y(n_4749)
);

BUFx3_ASAP7_75t_L g4750 ( 
.A(n_3954),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4204),
.B(n_3416),
.Y(n_4751)
);

OAI21x1_ASAP7_75t_SL g4752 ( 
.A1(n_4003),
.A2(n_3828),
.B(n_3537),
.Y(n_4752)
);

NOR2xp67_ASAP7_75t_L g4753 ( 
.A(n_4334),
.B(n_3413),
.Y(n_4753)
);

NOR2x1_ASAP7_75t_SL g4754 ( 
.A(n_4221),
.B(n_3721),
.Y(n_4754)
);

AND2x4_ASAP7_75t_L g4755 ( 
.A(n_4083),
.B(n_3908),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4159),
.Y(n_4756)
);

BUFx3_ASAP7_75t_L g4757 ( 
.A(n_3954),
.Y(n_4757)
);

AO31x2_ASAP7_75t_L g4758 ( 
.A1(n_4510),
.A2(n_3575),
.A3(n_3580),
.B(n_3607),
.Y(n_4758)
);

BUFx6f_ASAP7_75t_L g4759 ( 
.A(n_4036),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4164),
.Y(n_4760)
);

BUFx12f_ASAP7_75t_L g4761 ( 
.A(n_4136),
.Y(n_4761)
);

OAI21xp5_ASAP7_75t_L g4762 ( 
.A1(n_4268),
.A2(n_3655),
.B(n_3647),
.Y(n_4762)
);

INVx1_ASAP7_75t_L g4763 ( 
.A(n_4164),
.Y(n_4763)
);

INVx2_ASAP7_75t_SL g4764 ( 
.A(n_4036),
.Y(n_4764)
);

A2O1A1Ixp33_ASAP7_75t_L g4765 ( 
.A1(n_4281),
.A2(n_3801),
.B(n_3844),
.C(n_3927),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_SL g4766 ( 
.A(n_4068),
.B(n_4094),
.Y(n_4766)
);

INVx1_ASAP7_75t_SL g4767 ( 
.A(n_4146),
.Y(n_4767)
);

OAI21x1_ASAP7_75t_SL g4768 ( 
.A1(n_4003),
.A2(n_3823),
.B(n_3730),
.Y(n_4768)
);

BUFx5_ASAP7_75t_L g4769 ( 
.A(n_4288),
.Y(n_4769)
);

INVx1_ASAP7_75t_L g4770 ( 
.A(n_4175),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4175),
.Y(n_4771)
);

AOI21xp5_ASAP7_75t_L g4772 ( 
.A1(n_4077),
.A2(n_3523),
.B(n_3721),
.Y(n_4772)
);

NAND2x1p5_ASAP7_75t_L g4773 ( 
.A(n_4365),
.B(n_3413),
.Y(n_4773)
);

OAI21xp33_ASAP7_75t_SL g4774 ( 
.A1(n_4040),
.A2(n_3393),
.B(n_3444),
.Y(n_4774)
);

AOI22x1_ASAP7_75t_L g4775 ( 
.A1(n_4323),
.A2(n_3691),
.B1(n_3607),
.B2(n_3580),
.Y(n_4775)
);

AOI21x1_ASAP7_75t_L g4776 ( 
.A1(n_4147),
.A2(n_3687),
.B(n_3630),
.Y(n_4776)
);

NAND3xp33_ASAP7_75t_L g4777 ( 
.A(n_4349),
.B(n_4355),
.C(n_4097),
.Y(n_4777)
);

OAI22xp33_ASAP7_75t_L g4778 ( 
.A1(n_4246),
.A2(n_3795),
.B1(n_3822),
.B2(n_3871),
.Y(n_4778)
);

AOI221xp5_ASAP7_75t_L g4779 ( 
.A1(n_4024),
.A2(n_3867),
.B1(n_3840),
.B2(n_3860),
.C(n_3907),
.Y(n_4779)
);

A2O1A1Ixp33_ASAP7_75t_L g4780 ( 
.A1(n_4492),
.A2(n_3844),
.B(n_3801),
.C(n_3671),
.Y(n_4780)
);

AOI221xp5_ASAP7_75t_L g4781 ( 
.A1(n_4024),
.A2(n_3840),
.B1(n_3860),
.B2(n_3907),
.C(n_3916),
.Y(n_4781)
);

BUFx3_ASAP7_75t_L g4782 ( 
.A(n_3992),
.Y(n_4782)
);

INVx1_ASAP7_75t_L g4783 ( 
.A(n_4187),
.Y(n_4783)
);

A2O1A1Ixp33_ASAP7_75t_L g4784 ( 
.A1(n_4108),
.A2(n_3801),
.B(n_3671),
.C(n_3927),
.Y(n_4784)
);

AOI222xp33_ASAP7_75t_L g4785 ( 
.A1(n_4029),
.A2(n_3724),
.B1(n_3730),
.B2(n_3916),
.C1(n_3708),
.C2(n_3684),
.Y(n_4785)
);

OAI21x1_ASAP7_75t_L g4786 ( 
.A1(n_4243),
.A2(n_3880),
.B(n_3849),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4187),
.Y(n_4787)
);

AOI21x1_ASAP7_75t_L g4788 ( 
.A1(n_4099),
.A2(n_3687),
.B(n_3630),
.Y(n_4788)
);

OAI22xp5_ASAP7_75t_L g4789 ( 
.A1(n_4428),
.A2(n_4290),
.B1(n_4457),
.B2(n_4499),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4198),
.Y(n_4790)
);

OAI21x1_ASAP7_75t_L g4791 ( 
.A1(n_4336),
.A2(n_3880),
.B(n_3849),
.Y(n_4791)
);

BUFx10_ASAP7_75t_L g4792 ( 
.A(n_4370),
.Y(n_4792)
);

INVx1_ASAP7_75t_L g4793 ( 
.A(n_4198),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4139),
.A2(n_3523),
.B(n_3721),
.Y(n_4794)
);

INVxp67_ASAP7_75t_L g4795 ( 
.A(n_4079),
.Y(n_4795)
);

OAI221xp5_ASAP7_75t_L g4796 ( 
.A1(n_4037),
.A2(n_3898),
.B1(n_3883),
.B2(n_3880),
.C(n_3795),
.Y(n_4796)
);

OAI21x1_ASAP7_75t_L g4797 ( 
.A1(n_4336),
.A2(n_4104),
.B(n_4130),
.Y(n_4797)
);

A2O1A1Ixp33_ASAP7_75t_L g4798 ( 
.A1(n_4096),
.A2(n_4100),
.B(n_3959),
.C(n_4392),
.Y(n_4798)
);

OAI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_4318),
.A2(n_3749),
.B(n_3746),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4201),
.Y(n_4800)
);

OR2x2_ASAP7_75t_L g4801 ( 
.A(n_4222),
.B(n_3398),
.Y(n_4801)
);

OAI22xp5_ASAP7_75t_L g4802 ( 
.A1(n_4428),
.A2(n_3724),
.B1(n_3598),
.B2(n_3668),
.Y(n_4802)
);

AOI22xp33_ASAP7_75t_L g4803 ( 
.A1(n_4319),
.A2(n_3671),
.B1(n_3931),
.B2(n_3908),
.Y(n_4803)
);

AO21x2_ASAP7_75t_L g4804 ( 
.A1(n_4184),
.A2(n_3721),
.B(n_3858),
.Y(n_4804)
);

AOI22xp33_ASAP7_75t_L g4805 ( 
.A1(n_4319),
.A2(n_3671),
.B1(n_3908),
.B2(n_3931),
.Y(n_4805)
);

AOI21x1_ASAP7_75t_L g4806 ( 
.A1(n_4130),
.A2(n_3710),
.B(n_3687),
.Y(n_4806)
);

AOI221xp5_ASAP7_75t_L g4807 ( 
.A1(n_4029),
.A2(n_3943),
.B1(n_3942),
.B2(n_3936),
.C(n_3638),
.Y(n_4807)
);

INVxp67_ASAP7_75t_SL g4808 ( 
.A(n_4393),
.Y(n_4808)
);

INVx2_ASAP7_75t_SL g4809 ( 
.A(n_4036),
.Y(n_4809)
);

INVx2_ASAP7_75t_SL g4810 ( 
.A(n_4036),
.Y(n_4810)
);

NAND2x1_ASAP7_75t_L g4811 ( 
.A(n_4297),
.B(n_3444),
.Y(n_4811)
);

INVx1_ASAP7_75t_L g4812 ( 
.A(n_4201),
.Y(n_4812)
);

NAND2x1p5_ASAP7_75t_L g4813 ( 
.A(n_4365),
.B(n_3444),
.Y(n_4813)
);

AND2x4_ASAP7_75t_L g4814 ( 
.A(n_4083),
.B(n_3908),
.Y(n_4814)
);

AND2x2_ASAP7_75t_L g4815 ( 
.A(n_4249),
.B(n_3758),
.Y(n_4815)
);

INVx1_ASAP7_75t_L g4816 ( 
.A(n_4202),
.Y(n_4816)
);

AO21x2_ASAP7_75t_L g4817 ( 
.A1(n_4209),
.A2(n_4165),
.B(n_4041),
.Y(n_4817)
);

AOI221xp5_ASAP7_75t_L g4818 ( 
.A1(n_4489),
.A2(n_3943),
.B1(n_3942),
.B2(n_3936),
.C(n_3638),
.Y(n_4818)
);

AOI221xp5_ASAP7_75t_L g4819 ( 
.A1(n_4177),
.A2(n_3708),
.B1(n_3646),
.B2(n_3667),
.C(n_3668),
.Y(n_4819)
);

NAND2xp5_ASAP7_75t_L g4820 ( 
.A(n_4320),
.B(n_3416),
.Y(n_4820)
);

INVx3_ASAP7_75t_L g4821 ( 
.A(n_3997),
.Y(n_4821)
);

AOI22xp33_ASAP7_75t_L g4822 ( 
.A1(n_4321),
.A2(n_3931),
.B1(n_3874),
.B2(n_3809),
.Y(n_4822)
);

AND2x2_ASAP7_75t_L g4823 ( 
.A(n_3971),
.B(n_3931),
.Y(n_4823)
);

BUFx6f_ASAP7_75t_L g4824 ( 
.A(n_4262),
.Y(n_4824)
);

AOI21x1_ASAP7_75t_L g4825 ( 
.A1(n_4190),
.A2(n_3710),
.B(n_3854),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4013),
.B(n_3416),
.Y(n_4826)
);

AO21x2_ASAP7_75t_L g4827 ( 
.A1(n_4017),
.A2(n_3858),
.B(n_3751),
.Y(n_4827)
);

NAND2x1p5_ASAP7_75t_L g4828 ( 
.A(n_4401),
.B(n_3607),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4202),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4249),
.B(n_3696),
.Y(n_4830)
);

AO21x2_ASAP7_75t_L g4831 ( 
.A1(n_4496),
.A2(n_3858),
.B(n_3769),
.Y(n_4831)
);

OAI21x1_ASAP7_75t_SL g4832 ( 
.A1(n_4015),
.A2(n_3684),
.B(n_3694),
.Y(n_4832)
);

O2A1O1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_3976),
.A2(n_3694),
.B(n_3667),
.C(n_3646),
.Y(n_4833)
);

A2O1A1Ixp33_ASAP7_75t_L g4834 ( 
.A1(n_4399),
.A2(n_3809),
.B(n_3835),
.C(n_3874),
.Y(n_4834)
);

AND2x4_ASAP7_75t_L g4835 ( 
.A(n_4274),
.B(n_3575),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4361),
.A2(n_3598),
.B1(n_3719),
.B2(n_3918),
.Y(n_4836)
);

NOR2xp33_ASAP7_75t_L g4837 ( 
.A(n_4073),
.B(n_3918),
.Y(n_4837)
);

BUFx3_ASAP7_75t_L g4838 ( 
.A(n_3992),
.Y(n_4838)
);

OAI21x1_ASAP7_75t_SL g4839 ( 
.A1(n_4008),
.A2(n_3719),
.B(n_3575),
.Y(n_4839)
);

BUFx3_ASAP7_75t_L g4840 ( 
.A(n_3992),
.Y(n_4840)
);

AND2x4_ASAP7_75t_L g4841 ( 
.A(n_4274),
.B(n_3580),
.Y(n_4841)
);

OR2x2_ASAP7_75t_L g4842 ( 
.A(n_4222),
.B(n_3398),
.Y(n_4842)
);

OA21x2_ASAP7_75t_L g4843 ( 
.A1(n_4369),
.A2(n_3799),
.B(n_3837),
.Y(n_4843)
);

INVx1_ASAP7_75t_L g4844 ( 
.A(n_4226),
.Y(n_4844)
);

AOI21xp33_ASAP7_75t_L g4845 ( 
.A1(n_4043),
.A2(n_3938),
.B(n_3422),
.Y(n_4845)
);

INVx1_ASAP7_75t_SL g4846 ( 
.A(n_4306),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4226),
.Y(n_4847)
);

NOR2xp33_ASAP7_75t_L g4848 ( 
.A(n_4448),
.B(n_3685),
.Y(n_4848)
);

O2A1O1Ixp33_ASAP7_75t_L g4849 ( 
.A1(n_4480),
.A2(n_3938),
.B(n_3933),
.C(n_3925),
.Y(n_4849)
);

INVx1_ASAP7_75t_L g4850 ( 
.A(n_4229),
.Y(n_4850)
);

OA21x2_ASAP7_75t_L g4851 ( 
.A1(n_4472),
.A2(n_3845),
.B(n_3837),
.Y(n_4851)
);

AO21x2_ASAP7_75t_L g4852 ( 
.A1(n_3955),
.A2(n_3933),
.B(n_3925),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4229),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_SL g4854 ( 
.A(n_3958),
.B(n_3445),
.Y(n_4854)
);

BUFx3_ASAP7_75t_L g4855 ( 
.A(n_4030),
.Y(n_4855)
);

AND2x4_ASAP7_75t_L g4856 ( 
.A(n_4302),
.B(n_3691),
.Y(n_4856)
);

BUFx8_ASAP7_75t_L g4857 ( 
.A(n_4296),
.Y(n_4857)
);

OAI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_4246),
.A2(n_3616),
.B1(n_3662),
.B2(n_3445),
.Y(n_4858)
);

INVx1_ASAP7_75t_SL g4859 ( 
.A(n_4430),
.Y(n_4859)
);

INVx1_ASAP7_75t_SL g4860 ( 
.A(n_4010),
.Y(n_4860)
);

OAI22xp5_ASAP7_75t_L g4861 ( 
.A1(n_4375),
.A2(n_3847),
.B1(n_3861),
.B2(n_3835),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4020),
.B(n_3416),
.Y(n_4862)
);

AOI22xp33_ASAP7_75t_L g4863 ( 
.A1(n_4321),
.A2(n_3861),
.B1(n_3894),
.B2(n_3922),
.Y(n_4863)
);

NOR2xp33_ASAP7_75t_L g4864 ( 
.A(n_4060),
.B(n_3894),
.Y(n_4864)
);

INVx4_ASAP7_75t_SL g4865 ( 
.A(n_4342),
.Y(n_4865)
);

AOI22xp33_ASAP7_75t_L g4866 ( 
.A1(n_3985),
.A2(n_3922),
.B1(n_3616),
.B2(n_3445),
.Y(n_4866)
);

INVx1_ASAP7_75t_L g4867 ( 
.A(n_4233),
.Y(n_4867)
);

OAI21x1_ASAP7_75t_SL g4868 ( 
.A1(n_4379),
.A2(n_3691),
.B(n_3923),
.Y(n_4868)
);

A2O1A1Ixp33_ASAP7_75t_L g4869 ( 
.A1(n_4312),
.A2(n_3445),
.B(n_3616),
.C(n_3662),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4233),
.Y(n_4870)
);

XNOR2xp5_ASAP7_75t_L g4871 ( 
.A(n_4144),
.B(n_3620),
.Y(n_4871)
);

AND2x4_ASAP7_75t_L g4872 ( 
.A(n_4302),
.B(n_4339),
.Y(n_4872)
);

AO21x2_ASAP7_75t_L g4873 ( 
.A1(n_4148),
.A2(n_3909),
.B(n_3923),
.Y(n_4873)
);

NOR2x1_ASAP7_75t_SL g4874 ( 
.A(n_4221),
.B(n_3847),
.Y(n_4874)
);

OAI22xp33_ASAP7_75t_L g4875 ( 
.A1(n_4228),
.A2(n_3616),
.B1(n_3662),
.B2(n_3691),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4038),
.B(n_3416),
.Y(n_4876)
);

AND2x4_ASAP7_75t_L g4877 ( 
.A(n_4339),
.B(n_3407),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4237),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4093),
.B(n_3416),
.Y(n_4879)
);

OR2x6_ASAP7_75t_L g4880 ( 
.A(n_3972),
.B(n_3616),
.Y(n_4880)
);

BUFx2_ASAP7_75t_L g4881 ( 
.A(n_4421),
.Y(n_4881)
);

AO21x1_ASAP7_75t_L g4882 ( 
.A1(n_4350),
.A2(n_3912),
.B(n_3909),
.Y(n_4882)
);

OAI21x1_ASAP7_75t_L g4883 ( 
.A1(n_4097),
.A2(n_3902),
.B(n_3900),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4237),
.Y(n_4884)
);

AND2x4_ASAP7_75t_SL g4885 ( 
.A(n_4034),
.B(n_3616),
.Y(n_4885)
);

AOI21xp5_ASAP7_75t_L g4886 ( 
.A1(n_4173),
.A2(n_3422),
.B(n_3662),
.Y(n_4886)
);

INVx1_ASAP7_75t_L g4887 ( 
.A(n_4248),
.Y(n_4887)
);

AOI21xp33_ASAP7_75t_SL g4888 ( 
.A1(n_4479),
.A2(n_3422),
.B(n_3912),
.Y(n_4888)
);

BUFx8_ASAP7_75t_L g4889 ( 
.A(n_4296),
.Y(n_4889)
);

A2O1A1Ixp33_ASAP7_75t_SL g4890 ( 
.A1(n_4032),
.A2(n_3432),
.B(n_3457),
.C(n_3463),
.Y(n_4890)
);

O2A1O1Ixp5_ASAP7_75t_L g4891 ( 
.A1(n_4341),
.A2(n_3432),
.B(n_3457),
.C(n_3463),
.Y(n_4891)
);

CKINVDCx11_ASAP7_75t_R g4892 ( 
.A(n_4475),
.Y(n_4892)
);

OA21x2_ASAP7_75t_L g4893 ( 
.A1(n_4506),
.A2(n_3902),
.B(n_3886),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4248),
.Y(n_4894)
);

OAI22xp5_ASAP7_75t_L g4895 ( 
.A1(n_4376),
.A2(n_3620),
.B1(n_3701),
.B2(n_3747),
.Y(n_4895)
);

INVx4_ASAP7_75t_L g4896 ( 
.A(n_3958),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_L g4897 ( 
.A(n_4345),
.B(n_3407),
.Y(n_4897)
);

AOI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4495),
.A2(n_3662),
.B1(n_3635),
.B2(n_3701),
.Y(n_4898)
);

O2A1O1Ixp33_ASAP7_75t_SL g4899 ( 
.A1(n_4137),
.A2(n_3929),
.B(n_3892),
.C(n_3872),
.Y(n_4899)
);

OAI21xp5_ASAP7_75t_L g4900 ( 
.A1(n_4025),
.A2(n_3422),
.B(n_3785),
.Y(n_4900)
);

AOI22xp33_ASAP7_75t_L g4901 ( 
.A1(n_4495),
.A2(n_3662),
.B1(n_3635),
.B2(n_3747),
.Y(n_4901)
);

NAND3xp33_ASAP7_75t_L g4902 ( 
.A(n_4128),
.B(n_3748),
.C(n_3785),
.Y(n_4902)
);

NOR2xp33_ASAP7_75t_SL g4903 ( 
.A(n_4115),
.B(n_2419),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4250),
.Y(n_4904)
);

AOI22xp5_ASAP7_75t_L g4905 ( 
.A1(n_4153),
.A2(n_3805),
.B1(n_3748),
.B2(n_2642),
.Y(n_4905)
);

AOI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4154),
.A2(n_3805),
.B1(n_2642),
.B2(n_2810),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4250),
.Y(n_4907)
);

OR2x6_ASAP7_75t_L g4908 ( 
.A(n_3964),
.B(n_3872),
.Y(n_4908)
);

AO21x2_ASAP7_75t_L g4909 ( 
.A1(n_4000),
.A2(n_3722),
.B(n_3872),
.Y(n_4909)
);

INVx1_ASAP7_75t_L g4910 ( 
.A(n_4280),
.Y(n_4910)
);

AOI21x1_ASAP7_75t_L g4911 ( 
.A1(n_4190),
.A2(n_3722),
.B(n_3869),
.Y(n_4911)
);

NAND2xp5_ASAP7_75t_SL g4912 ( 
.A(n_3958),
.B(n_3786),
.Y(n_4912)
);

OAI21xp5_ASAP7_75t_L g4913 ( 
.A1(n_4033),
.A2(n_3786),
.B(n_3869),
.Y(n_4913)
);

AO21x2_ASAP7_75t_L g4914 ( 
.A1(n_4156),
.A2(n_4267),
.B(n_4265),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4280),
.Y(n_4915)
);

AO22x2_ASAP7_75t_L g4916 ( 
.A1(n_4307),
.A2(n_3739),
.B1(n_3854),
.B2(n_3832),
.Y(n_4916)
);

OAI221xp5_ASAP7_75t_L g4917 ( 
.A1(n_4039),
.A2(n_4386),
.B1(n_4366),
.B2(n_4322),
.C(n_4379),
.Y(n_4917)
);

AOI21xp33_ASAP7_75t_L g4918 ( 
.A1(n_4086),
.A2(n_3786),
.B(n_3739),
.Y(n_4918)
);

NAND2xp5_ASAP7_75t_L g4919 ( 
.A(n_4381),
.B(n_3407),
.Y(n_4919)
);

CKINVDCx8_ASAP7_75t_R g4920 ( 
.A(n_3967),
.Y(n_4920)
);

BUFx4f_ASAP7_75t_SL g4921 ( 
.A(n_4030),
.Y(n_4921)
);

AO22x2_ASAP7_75t_L g4922 ( 
.A1(n_4309),
.A2(n_3797),
.B1(n_3696),
.B2(n_3472),
.Y(n_4922)
);

BUFx2_ASAP7_75t_L g4923 ( 
.A(n_4421),
.Y(n_4923)
);

OR2x6_ASAP7_75t_L g4924 ( 
.A(n_4240),
.B(n_2643),
.Y(n_4924)
);

OA21x2_ASAP7_75t_L g4925 ( 
.A1(n_4215),
.A2(n_3411),
.B(n_3696),
.Y(n_4925)
);

OAI21x1_ASAP7_75t_L g4926 ( 
.A1(n_4215),
.A2(n_4494),
.B(n_4181),
.Y(n_4926)
);

NOR2x1_ASAP7_75t_L g4927 ( 
.A(n_4030),
.B(n_3696),
.Y(n_4927)
);

OAI22xp33_ASAP7_75t_L g4928 ( 
.A1(n_4228),
.A2(n_2724),
.B1(n_2438),
.B2(n_2464),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4447),
.B(n_3696),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4409),
.B(n_3407),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4305),
.Y(n_4931)
);

INVx3_ASAP7_75t_L g4932 ( 
.A(n_4095),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4305),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4315),
.Y(n_4934)
);

INVx3_ASAP7_75t_L g4935 ( 
.A(n_4095),
.Y(n_4935)
);

CKINVDCx20_ASAP7_75t_R g4936 ( 
.A(n_4144),
.Y(n_4936)
);

AOI21x1_ASAP7_75t_L g4937 ( 
.A1(n_4380),
.A2(n_3472),
.B(n_3411),
.Y(n_4937)
);

OAI21x1_ASAP7_75t_L g4938 ( 
.A1(n_4494),
.A2(n_3411),
.B(n_3483),
.Y(n_4938)
);

OAI21x1_ASAP7_75t_L g4939 ( 
.A1(n_4181),
.A2(n_3411),
.B(n_3483),
.Y(n_4939)
);

O2A1O1Ixp33_ASAP7_75t_SL g4940 ( 
.A1(n_4137),
.A2(n_3472),
.B(n_3407),
.C(n_3411),
.Y(n_4940)
);

AND2x2_ASAP7_75t_L g4941 ( 
.A(n_4447),
.B(n_3472),
.Y(n_4941)
);

O2A1O1Ixp33_ASAP7_75t_L g4942 ( 
.A1(n_4313),
.A2(n_3551),
.B(n_3407),
.C(n_3472),
.Y(n_4942)
);

NOR2xp33_ASAP7_75t_SL g4943 ( 
.A(n_4115),
.B(n_2419),
.Y(n_4943)
);

OAI21x1_ASAP7_75t_L g4944 ( 
.A1(n_4347),
.A2(n_3483),
.B(n_3442),
.Y(n_4944)
);

OAI21xp5_ASAP7_75t_L g4945 ( 
.A1(n_4261),
.A2(n_2810),
.B(n_3551),
.Y(n_4945)
);

BUFx6f_ASAP7_75t_L g4946 ( 
.A(n_4262),
.Y(n_4946)
);

OAI21x1_ASAP7_75t_L g4947 ( 
.A1(n_4286),
.A2(n_3483),
.B(n_3442),
.Y(n_4947)
);

NAND2xp5_ASAP7_75t_L g4948 ( 
.A(n_4067),
.B(n_3538),
.Y(n_4948)
);

OAI21x1_ASAP7_75t_L g4949 ( 
.A1(n_4286),
.A2(n_3483),
.B(n_3442),
.Y(n_4949)
);

OAI21xp5_ASAP7_75t_L g4950 ( 
.A1(n_4150),
.A2(n_2810),
.B(n_3551),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4315),
.Y(n_4951)
);

AOI22xp33_ASAP7_75t_L g4952 ( 
.A1(n_4503),
.A2(n_2721),
.B1(n_2810),
.B2(n_2464),
.Y(n_4952)
);

INVxp67_ASAP7_75t_SL g4953 ( 
.A(n_4414),
.Y(n_4953)
);

BUFx3_ASAP7_75t_L g4954 ( 
.A(n_4054),
.Y(n_4954)
);

AND2x4_ASAP7_75t_L g4955 ( 
.A(n_4462),
.B(n_3442),
.Y(n_4955)
);

OAI22xp5_ASAP7_75t_L g4956 ( 
.A1(n_4386),
.A2(n_2549),
.B1(n_2438),
.B2(n_2464),
.Y(n_4956)
);

CKINVDCx5p33_ASAP7_75t_R g4957 ( 
.A(n_4388),
.Y(n_4957)
);

OAI21x1_ASAP7_75t_L g4958 ( 
.A1(n_4310),
.A2(n_3483),
.B(n_3442),
.Y(n_4958)
);

AOI21x1_ASAP7_75t_L g4959 ( 
.A1(n_4401),
.A2(n_3472),
.B(n_3442),
.Y(n_4959)
);

NAND3xp33_ASAP7_75t_L g4960 ( 
.A(n_3991),
.B(n_2721),
.C(n_2438),
.Y(n_4960)
);

INVx1_ASAP7_75t_SL g4961 ( 
.A(n_4488),
.Y(n_4961)
);

AND2x4_ASAP7_75t_L g4962 ( 
.A(n_4463),
.B(n_3815),
.Y(n_4962)
);

OA21x2_ASAP7_75t_L g4963 ( 
.A1(n_4458),
.A2(n_3423),
.B(n_3538),
.Y(n_4963)
);

OAI21x1_ASAP7_75t_L g4964 ( 
.A1(n_4310),
.A2(n_3423),
.B(n_3538),
.Y(n_4964)
);

OA21x2_ASAP7_75t_L g4965 ( 
.A1(n_4464),
.A2(n_4207),
.B(n_4285),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4325),
.Y(n_4966)
);

NAND2x1p5_ASAP7_75t_L g4967 ( 
.A(n_4463),
.B(n_2551),
.Y(n_4967)
);

OAI21x1_ASAP7_75t_L g4968 ( 
.A1(n_4259),
.A2(n_3423),
.B(n_3538),
.Y(n_4968)
);

AND2x2_ASAP7_75t_L g4969 ( 
.A(n_4253),
.B(n_3551),
.Y(n_4969)
);

AOI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4287),
.A2(n_2551),
.B(n_2438),
.Y(n_4970)
);

OR2x2_ASAP7_75t_L g4971 ( 
.A(n_4391),
.B(n_3603),
.Y(n_4971)
);

OAI21x1_ASAP7_75t_SL g4972 ( 
.A1(n_4374),
.A2(n_2419),
.B(n_2528),
.Y(n_4972)
);

OAI21x1_ASAP7_75t_L g4973 ( 
.A1(n_4269),
.A2(n_3423),
.B(n_3538),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4325),
.Y(n_4974)
);

INVx1_ASAP7_75t_SL g4975 ( 
.A(n_4488),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4326),
.Y(n_4976)
);

OA21x2_ASAP7_75t_L g4977 ( 
.A1(n_4207),
.A2(n_3423),
.B(n_3610),
.Y(n_4977)
);

INVx1_ASAP7_75t_L g4978 ( 
.A(n_4326),
.Y(n_4978)
);

BUFx2_ASAP7_75t_L g4979 ( 
.A(n_4054),
.Y(n_4979)
);

AO21x2_ASAP7_75t_L g4980 ( 
.A1(n_4156),
.A2(n_4301),
.B(n_4172),
.Y(n_4980)
);

OAI21x1_ASAP7_75t_L g4981 ( 
.A1(n_4269),
.A2(n_3774),
.B(n_3611),
.Y(n_4981)
);

NAND3xp33_ASAP7_75t_L g4982 ( 
.A(n_3991),
.B(n_2721),
.C(n_2438),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4001),
.B(n_3774),
.Y(n_4983)
);

OAI21x1_ASAP7_75t_L g4984 ( 
.A1(n_4219),
.A2(n_3774),
.B(n_3611),
.Y(n_4984)
);

OAI21x1_ASAP7_75t_L g4985 ( 
.A1(n_4219),
.A2(n_4284),
.B(n_4314),
.Y(n_4985)
);

NAND2x1p5_ASAP7_75t_L g4986 ( 
.A(n_4018),
.B(n_2643),
.Y(n_4986)
);

AO21x2_ASAP7_75t_L g4987 ( 
.A1(n_4032),
.A2(n_3774),
.B(n_3611),
.Y(n_4987)
);

OAI21x1_ASAP7_75t_L g4988 ( 
.A1(n_4219),
.A2(n_3737),
.B(n_3782),
.Y(n_4988)
);

AOI21xp5_ASAP7_75t_L g4989 ( 
.A1(n_4363),
.A2(n_2643),
.B(n_2438),
.Y(n_4989)
);

OAI21x1_ASAP7_75t_L g4990 ( 
.A1(n_4219),
.A2(n_3782),
.B(n_3611),
.Y(n_4990)
);

BUFx3_ASAP7_75t_L g4991 ( 
.A(n_4054),
.Y(n_4991)
);

AO21x2_ASAP7_75t_L g4992 ( 
.A1(n_4052),
.A2(n_3782),
.B(n_3611),
.Y(n_4992)
);

INVx8_ASAP7_75t_L g4993 ( 
.A(n_3967),
.Y(n_4993)
);

BUFx10_ASAP7_75t_L g4994 ( 
.A(n_3967),
.Y(n_4994)
);

AND2x4_ASAP7_75t_L g4995 ( 
.A(n_4117),
.B(n_3815),
.Y(n_4995)
);

OA21x2_ASAP7_75t_L g4996 ( 
.A1(n_4511),
.A2(n_3610),
.B(n_3603),
.Y(n_4996)
);

OAI21x1_ASAP7_75t_L g4997 ( 
.A1(n_4284),
.A2(n_3737),
.B(n_3782),
.Y(n_4997)
);

A2O1A1Ixp33_ASAP7_75t_L g4998 ( 
.A1(n_4263),
.A2(n_3610),
.B(n_2464),
.C(n_2466),
.Y(n_4998)
);

HB1xp67_ASAP7_75t_L g4999 ( 
.A(n_4486),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4333),
.Y(n_5000)
);

OAI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_3974),
.A2(n_2810),
.B(n_3610),
.Y(n_5001)
);

INVx4_ASAP7_75t_L g5002 ( 
.A(n_3958),
.Y(n_5002)
);

AND2x4_ASAP7_75t_L g5003 ( 
.A(n_4117),
.B(n_3815),
.Y(n_5003)
);

AND2x4_ASAP7_75t_SL g5004 ( 
.A(n_4034),
.B(n_4007),
.Y(n_5004)
);

OA21x2_ASAP7_75t_L g5005 ( 
.A1(n_4511),
.A2(n_3610),
.B(n_3603),
.Y(n_5005)
);

OA21x2_ASAP7_75t_L g5006 ( 
.A1(n_4132),
.A2(n_3603),
.B(n_3782),
.Y(n_5006)
);

AOI21xp5_ASAP7_75t_L g5007 ( 
.A1(n_4367),
.A2(n_2643),
.B(n_2464),
.Y(n_5007)
);

OAI21x1_ASAP7_75t_L g5008 ( 
.A1(n_4351),
.A2(n_3782),
.B(n_3737),
.Y(n_5008)
);

BUFx3_ASAP7_75t_L g5009 ( 
.A(n_3967),
.Y(n_5009)
);

NOR2x1_ASAP7_75t_SL g5010 ( 
.A(n_4221),
.B(n_3603),
.Y(n_5010)
);

OAI21x1_ASAP7_75t_L g5011 ( 
.A1(n_4353),
.A2(n_3706),
.B(n_3737),
.Y(n_5011)
);

INVx3_ASAP7_75t_L g5012 ( 
.A(n_4095),
.Y(n_5012)
);

AND2x2_ASAP7_75t_L g5013 ( 
.A(n_3971),
.B(n_3603),
.Y(n_5013)
);

INVxp67_ASAP7_75t_SL g5014 ( 
.A(n_4140),
.Y(n_5014)
);

AOI21xp5_ASAP7_75t_L g5015 ( 
.A1(n_4766),
.A2(n_4377),
.B(n_4230),
.Y(n_5015)
);

BUFx2_ASAP7_75t_L g5016 ( 
.A(n_4857),
.Y(n_5016)
);

AOI21xp5_ASAP7_75t_L g5017 ( 
.A1(n_4537),
.A2(n_4520),
.B(n_4044),
.Y(n_5017)
);

OAI22xp5_ASAP7_75t_L g5018 ( 
.A1(n_4544),
.A2(n_4403),
.B1(n_4427),
.B2(n_4407),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4533),
.B(n_3963),
.Y(n_5019)
);

BUFx3_ASAP7_75t_L g5020 ( 
.A(n_4566),
.Y(n_5020)
);

AND2x2_ASAP7_75t_L g5021 ( 
.A(n_4570),
.B(n_3995),
.Y(n_5021)
);

O2A1O1Ixp5_ASAP7_75t_L g5022 ( 
.A1(n_4530),
.A2(n_4411),
.B(n_4387),
.C(n_4438),
.Y(n_5022)
);

INVx1_ASAP7_75t_L g5023 ( 
.A(n_4525),
.Y(n_5023)
);

CKINVDCx5p33_ASAP7_75t_R g5024 ( 
.A(n_4742),
.Y(n_5024)
);

AOI21xp5_ASAP7_75t_L g5025 ( 
.A1(n_4537),
.A2(n_4044),
.B(n_4185),
.Y(n_5025)
);

OA21x2_ASAP7_75t_L g5026 ( 
.A1(n_4586),
.A2(n_4052),
.B(n_4088),
.Y(n_5026)
);

NAND2xp5_ASAP7_75t_L g5027 ( 
.A(n_4533),
.B(n_4170),
.Y(n_5027)
);

NAND2xp5_ASAP7_75t_L g5028 ( 
.A(n_4860),
.B(n_4785),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4525),
.Y(n_5029)
);

OA21x2_ASAP7_75t_L g5030 ( 
.A1(n_4586),
.A2(n_4715),
.B(n_4988),
.Y(n_5030)
);

AOI21xp33_ASAP7_75t_SL g5031 ( 
.A1(n_4592),
.A2(n_4035),
.B(n_4404),
.Y(n_5031)
);

OAI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_4530),
.A2(n_3990),
.B(n_4019),
.Y(n_5032)
);

NOR2xp33_ASAP7_75t_L g5033 ( 
.A(n_4592),
.B(n_4007),
.Y(n_5033)
);

OA21x2_ASAP7_75t_L g5034 ( 
.A1(n_4715),
.A2(n_4088),
.B(n_4102),
.Y(n_5034)
);

NAND2xp5_ASAP7_75t_L g5035 ( 
.A(n_4860),
.B(n_4180),
.Y(n_5035)
);

BUFx10_ASAP7_75t_L g5036 ( 
.A(n_4568),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_L g5037 ( 
.A(n_4785),
.B(n_3988),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4542),
.Y(n_5038)
);

BUFx2_ASAP7_75t_L g5039 ( 
.A(n_4857),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4781),
.B(n_3988),
.Y(n_5040)
);

OAI22xp5_ASAP7_75t_L g5041 ( 
.A1(n_4544),
.A2(n_4482),
.B1(n_3982),
.B2(n_4362),
.Y(n_5041)
);

INVx1_ASAP7_75t_L g5042 ( 
.A(n_4542),
.Y(n_5042)
);

OAI21x1_ASAP7_75t_L g5043 ( 
.A1(n_4776),
.A2(n_3991),
.B(n_4123),
.Y(n_5043)
);

NAND2x1p5_ASAP7_75t_L g5044 ( 
.A(n_4606),
.B(n_4487),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4549),
.Y(n_5045)
);

OAI21x1_ASAP7_75t_L g5046 ( 
.A1(n_4776),
.A2(n_3991),
.B(n_4123),
.Y(n_5046)
);

AO21x2_ASAP7_75t_L g5047 ( 
.A1(n_4597),
.A2(n_4251),
.B(n_4333),
.Y(n_5047)
);

OR2x6_ASAP7_75t_L g5048 ( 
.A(n_4606),
.B(n_4214),
.Y(n_5048)
);

AO31x2_ASAP7_75t_L g5049 ( 
.A1(n_4572),
.A2(n_4443),
.A3(n_4007),
.B(n_4487),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4549),
.Y(n_5050)
);

OAI22xp33_ASAP7_75t_L g5051 ( 
.A1(n_4572),
.A2(n_4382),
.B1(n_4482),
.B2(n_4103),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_4781),
.B(n_4163),
.Y(n_5052)
);

NAND3xp33_ASAP7_75t_L g5053 ( 
.A(n_4596),
.B(n_4112),
.C(n_4102),
.Y(n_5053)
);

BUFx6f_ASAP7_75t_L g5054 ( 
.A(n_4566),
.Y(n_5054)
);

BUFx12f_ASAP7_75t_L g5055 ( 
.A(n_4566),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_4807),
.B(n_4182),
.Y(n_5056)
);

INVxp67_ASAP7_75t_SL g5057 ( 
.A(n_4734),
.Y(n_5057)
);

INVx2_ASAP7_75t_SL g5058 ( 
.A(n_4792),
.Y(n_5058)
);

AOI22xp33_ASAP7_75t_L g5059 ( 
.A1(n_4596),
.A2(n_4446),
.B1(n_4503),
.B2(n_4186),
.Y(n_5059)
);

NOR2xp33_ASAP7_75t_SL g5060 ( 
.A(n_4574),
.B(n_4007),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4565),
.Y(n_5061)
);

A2O1A1Ixp33_ASAP7_75t_L g5062 ( 
.A1(n_4526),
.A2(n_4433),
.B(n_4446),
.C(n_4366),
.Y(n_5062)
);

OR2x6_ASAP7_75t_L g5063 ( 
.A(n_4546),
.B(n_4216),
.Y(n_5063)
);

HB1xp67_ASAP7_75t_L g5064 ( 
.A(n_4583),
.Y(n_5064)
);

OAI21x1_ASAP7_75t_L g5065 ( 
.A1(n_4597),
.A2(n_4985),
.B(n_4687),
.Y(n_5065)
);

INVx2_ASAP7_75t_L g5066 ( 
.A(n_4545),
.Y(n_5066)
);

AOI21xp33_ASAP7_75t_SL g5067 ( 
.A1(n_4592),
.A2(n_4346),
.B(n_4342),
.Y(n_5067)
);

AO31x2_ASAP7_75t_L g5068 ( 
.A1(n_4539),
.A2(n_4487),
.A3(n_4505),
.B(n_4402),
.Y(n_5068)
);

OAI21x1_ASAP7_75t_L g5069 ( 
.A1(n_4985),
.A2(n_4231),
.B(n_4123),
.Y(n_5069)
);

INVx2_ASAP7_75t_L g5070 ( 
.A(n_4545),
.Y(n_5070)
);

OAI22xp5_ASAP7_75t_L g5071 ( 
.A1(n_4543),
.A2(n_4329),
.B1(n_4398),
.B2(n_4374),
.Y(n_5071)
);

INVx2_ASAP7_75t_SL g5072 ( 
.A(n_4792),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4565),
.Y(n_5073)
);

INVx1_ASAP7_75t_L g5074 ( 
.A(n_4576),
.Y(n_5074)
);

AOI22xp33_ASAP7_75t_L g5075 ( 
.A1(n_4917),
.A2(n_4789),
.B1(n_4567),
.B2(n_4526),
.Y(n_5075)
);

AOI21xp5_ASAP7_75t_L g5076 ( 
.A1(n_4798),
.A2(n_4044),
.B(n_4185),
.Y(n_5076)
);

AOI22xp33_ASAP7_75t_L g5077 ( 
.A1(n_4917),
.A2(n_4186),
.B1(n_4322),
.B2(n_4433),
.Y(n_5077)
);

AOI21xp5_ASAP7_75t_L g5078 ( 
.A1(n_4659),
.A2(n_4044),
.B(n_4303),
.Y(n_5078)
);

OA21x2_ASAP7_75t_L g5079 ( 
.A1(n_4988),
.A2(n_4354),
.B(n_4344),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4807),
.B(n_4436),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_4570),
.B(n_3995),
.Y(n_5081)
);

INVx1_ASAP7_75t_L g5082 ( 
.A(n_4576),
.Y(n_5082)
);

BUFx2_ASAP7_75t_L g5083 ( 
.A(n_4857),
.Y(n_5083)
);

OAI21x1_ASAP7_75t_L g5084 ( 
.A1(n_4985),
.A2(n_4238),
.B(n_4231),
.Y(n_5084)
);

INVx2_ASAP7_75t_L g5085 ( 
.A(n_4545),
.Y(n_5085)
);

BUFx2_ASAP7_75t_L g5086 ( 
.A(n_4857),
.Y(n_5086)
);

HB1xp67_ASAP7_75t_L g5087 ( 
.A(n_4583),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_L g5088 ( 
.A(n_4779),
.B(n_4439),
.Y(n_5088)
);

NOR2xp33_ASAP7_75t_L g5089 ( 
.A(n_4538),
.B(n_3967),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_4587),
.Y(n_5090)
);

BUFx2_ASAP7_75t_L g5091 ( 
.A(n_4889),
.Y(n_5091)
);

OAI21xp5_ASAP7_75t_L g5092 ( 
.A1(n_4539),
.A2(n_4551),
.B(n_4523),
.Y(n_5092)
);

NAND2xp5_ASAP7_75t_L g5093 ( 
.A(n_4779),
.B(n_4224),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4587),
.Y(n_5094)
);

INVx3_ASAP7_75t_L g5095 ( 
.A(n_4624),
.Y(n_5095)
);

NOR2xp33_ASAP7_75t_L g5096 ( 
.A(n_4538),
.B(n_3993),
.Y(n_5096)
);

AOI21x1_ASAP7_75t_L g5097 ( 
.A1(n_4979),
.A2(n_4061),
.B(n_4344),
.Y(n_5097)
);

OA21x2_ASAP7_75t_L g5098 ( 
.A1(n_4988),
.A2(n_4356),
.B(n_4354),
.Y(n_5098)
);

BUFx2_ASAP7_75t_R g5099 ( 
.A(n_4957),
.Y(n_5099)
);

AOI21x1_ASAP7_75t_L g5100 ( 
.A1(n_4979),
.A2(n_4061),
.B(n_4356),
.Y(n_5100)
);

INVx2_ASAP7_75t_L g5101 ( 
.A(n_4545),
.Y(n_5101)
);

AO21x2_ASAP7_75t_L g5102 ( 
.A1(n_4707),
.A2(n_4359),
.B(n_4358),
.Y(n_5102)
);

OAI21x1_ASAP7_75t_L g5103 ( 
.A1(n_4687),
.A2(n_4238),
.B(n_4231),
.Y(n_5103)
);

OA21x2_ASAP7_75t_L g5104 ( 
.A1(n_4990),
.A2(n_4359),
.B(n_4358),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_4588),
.Y(n_5105)
);

INVx2_ASAP7_75t_L g5106 ( 
.A(n_4545),
.Y(n_5106)
);

HB1xp67_ASAP7_75t_L g5107 ( 
.A(n_4795),
.Y(n_5107)
);

BUFx3_ASAP7_75t_L g5108 ( 
.A(n_4633),
.Y(n_5108)
);

INVx1_ASAP7_75t_L g5109 ( 
.A(n_4588),
.Y(n_5109)
);

AND2x4_ASAP7_75t_L g5110 ( 
.A(n_4558),
.B(n_3995),
.Y(n_5110)
);

AND2x2_ASAP7_75t_L g5111 ( 
.A(n_4570),
.B(n_3960),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4593),
.Y(n_5112)
);

HB1xp67_ASAP7_75t_L g5113 ( 
.A(n_4795),
.Y(n_5113)
);

BUFx4_ASAP7_75t_R g5114 ( 
.A(n_4792),
.Y(n_5114)
);

AOI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_4523),
.A2(n_4044),
.B(n_4303),
.Y(n_5115)
);

OR2x2_ASAP7_75t_L g5116 ( 
.A(n_4581),
.B(n_4560),
.Y(n_5116)
);

OAI22xp5_ASAP7_75t_L g5117 ( 
.A1(n_4543),
.A2(n_4021),
.B1(n_4408),
.B2(n_3987),
.Y(n_5117)
);

OAI21x1_ASAP7_75t_L g5118 ( 
.A1(n_4687),
.A2(n_4327),
.B(n_4238),
.Y(n_5118)
);

OAI21x1_ASAP7_75t_L g5119 ( 
.A1(n_4687),
.A2(n_4327),
.B(n_4417),
.Y(n_5119)
);

AO31x2_ASAP7_75t_L g5120 ( 
.A1(n_4550),
.A2(n_4487),
.A3(n_4091),
.B(n_4402),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_4561),
.B(n_4224),
.Y(n_5121)
);

OAI21xp5_ASAP7_75t_L g5122 ( 
.A1(n_4551),
.A2(n_4316),
.B(n_4368),
.Y(n_5122)
);

AOI22xp5_ASAP7_75t_L g5123 ( 
.A1(n_4789),
.A2(n_4131),
.B1(n_4169),
.B2(n_4117),
.Y(n_5123)
);

AND2x4_ASAP7_75t_L g5124 ( 
.A(n_4558),
.B(n_4221),
.Y(n_5124)
);

OA21x2_ASAP7_75t_L g5125 ( 
.A1(n_4984),
.A2(n_4422),
.B(n_4420),
.Y(n_5125)
);

NAND2x1p5_ASAP7_75t_L g5126 ( 
.A(n_4624),
.B(n_4117),
.Y(n_5126)
);

OAI21x1_ASAP7_75t_L g5127 ( 
.A1(n_4662),
.A2(n_4327),
.B(n_4417),
.Y(n_5127)
);

A2O1A1Ixp33_ASAP7_75t_L g5128 ( 
.A1(n_4833),
.A2(n_4304),
.B(n_4412),
.C(n_4396),
.Y(n_5128)
);

CKINVDCx20_ASAP7_75t_R g5129 ( 
.A(n_4578),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_L g5130 ( 
.A(n_4561),
.B(n_4235),
.Y(n_5130)
);

HB1xp67_ASAP7_75t_L g5131 ( 
.A(n_4767),
.Y(n_5131)
);

NAND2x1p5_ASAP7_75t_L g5132 ( 
.A(n_4624),
.B(n_4131),
.Y(n_5132)
);

OA21x2_ASAP7_75t_L g5133 ( 
.A1(n_4984),
.A2(n_4422),
.B(n_4420),
.Y(n_5133)
);

INVx1_ASAP7_75t_L g5134 ( 
.A(n_4593),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_4595),
.Y(n_5135)
);

OAI21x1_ASAP7_75t_L g5136 ( 
.A1(n_4662),
.A2(n_4435),
.B(n_4419),
.Y(n_5136)
);

OAI21x1_ASAP7_75t_L g5137 ( 
.A1(n_4662),
.A2(n_4435),
.B(n_4419),
.Y(n_5137)
);

NOR2xp33_ASAP7_75t_L g5138 ( 
.A(n_4538),
.B(n_4633),
.Y(n_5138)
);

INVx2_ASAP7_75t_L g5139 ( 
.A(n_4545),
.Y(n_5139)
);

AO31x2_ASAP7_75t_L g5140 ( 
.A1(n_4550),
.A2(n_4091),
.A3(n_4402),
.B(n_4431),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_4625),
.A2(n_4304),
.B(n_4478),
.Y(n_5141)
);

AOI21xp5_ASAP7_75t_L g5142 ( 
.A1(n_4625),
.A2(n_4484),
.B(n_4514),
.Y(n_5142)
);

OA21x2_ASAP7_75t_L g5143 ( 
.A1(n_4984),
.A2(n_4441),
.B(n_4431),
.Y(n_5143)
);

AOI21xp5_ASAP7_75t_L g5144 ( 
.A1(n_4579),
.A2(n_4234),
.B(n_4423),
.Y(n_5144)
);

INVx2_ASAP7_75t_L g5145 ( 
.A(n_4545),
.Y(n_5145)
);

AND2x2_ASAP7_75t_L g5146 ( 
.A(n_4589),
.B(n_3960),
.Y(n_5146)
);

OR2x2_ASAP7_75t_L g5147 ( 
.A(n_4581),
.B(n_4413),
.Y(n_5147)
);

INVx1_ASAP7_75t_L g5148 ( 
.A(n_4595),
.Y(n_5148)
);

AOI21x1_ASAP7_75t_L g5149 ( 
.A1(n_4734),
.A2(n_4061),
.B(n_4441),
.Y(n_5149)
);

AOI21x1_ASAP7_75t_L g5150 ( 
.A1(n_4811),
.A2(n_4911),
.B(n_4825),
.Y(n_5150)
);

AOI21xp5_ASAP7_75t_L g5151 ( 
.A1(n_4579),
.A2(n_4452),
.B(n_4394),
.Y(n_5151)
);

AO21x1_ASAP7_75t_L g5152 ( 
.A1(n_4552),
.A2(n_4500),
.B(n_4467),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4617),
.B(n_4684),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_4599),
.Y(n_5154)
);

AOI21x1_ASAP7_75t_L g5155 ( 
.A1(n_4811),
.A2(n_4061),
.B(n_4467),
.Y(n_5155)
);

OR2x2_ASAP7_75t_L g5156 ( 
.A(n_4560),
.B(n_4897),
.Y(n_5156)
);

BUFx12f_ASAP7_75t_L g5157 ( 
.A(n_4633),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_4617),
.B(n_4235),
.Y(n_5158)
);

AND2x2_ASAP7_75t_L g5159 ( 
.A(n_4589),
.B(n_4253),
.Y(n_5159)
);

NAND2xp5_ASAP7_75t_L g5160 ( 
.A(n_4684),
.B(n_4048),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_4599),
.Y(n_5161)
);

OA21x2_ASAP7_75t_L g5162 ( 
.A1(n_4772),
.A2(n_4794),
.B(n_4964),
.Y(n_5162)
);

INVx1_ASAP7_75t_L g5163 ( 
.A(n_4608),
.Y(n_5163)
);

AO31x2_ASAP7_75t_L g5164 ( 
.A1(n_4874),
.A2(n_4091),
.A3(n_4402),
.B(n_4500),
.Y(n_5164)
);

INVx2_ASAP7_75t_L g5165 ( 
.A(n_4650),
.Y(n_5165)
);

AND2x2_ASAP7_75t_L g5166 ( 
.A(n_4589),
.B(n_4253),
.Y(n_5166)
);

BUFx2_ASAP7_75t_L g5167 ( 
.A(n_4889),
.Y(n_5167)
);

AOI22xp5_ASAP7_75t_L g5168 ( 
.A1(n_4567),
.A2(n_4200),
.B1(n_4208),
.B2(n_4116),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_4608),
.Y(n_5169)
);

NAND2xp5_ASAP7_75t_L g5170 ( 
.A(n_4562),
.B(n_4107),
.Y(n_5170)
);

OAI21x1_ASAP7_75t_L g5171 ( 
.A1(n_4521),
.A2(n_4455),
.B(n_4453),
.Y(n_5171)
);

OAI21x1_ASAP7_75t_SL g5172 ( 
.A1(n_4882),
.A2(n_4091),
.B(n_4426),
.Y(n_5172)
);

INVx1_ASAP7_75t_L g5173 ( 
.A(n_4609),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_L g5174 ( 
.A(n_4562),
.B(n_4616),
.Y(n_5174)
);

HB1xp67_ASAP7_75t_L g5175 ( 
.A(n_4767),
.Y(n_5175)
);

AOI21xp5_ASAP7_75t_L g5176 ( 
.A1(n_4707),
.A2(n_4378),
.B(n_4122),
.Y(n_5176)
);

INVx2_ASAP7_75t_L g5177 ( 
.A(n_4650),
.Y(n_5177)
);

A2O1A1Ixp33_ASAP7_75t_L g5178 ( 
.A1(n_4833),
.A2(n_4477),
.B(n_4122),
.C(n_4119),
.Y(n_5178)
);

AO21x2_ASAP7_75t_L g5179 ( 
.A1(n_4888),
.A2(n_4177),
.B(n_4453),
.Y(n_5179)
);

AND2x4_ASAP7_75t_L g5180 ( 
.A(n_4558),
.B(n_4131),
.Y(n_5180)
);

AND2x4_ASAP7_75t_L g5181 ( 
.A(n_4558),
.B(n_4131),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_4609),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_4598),
.A2(n_4470),
.B(n_4465),
.Y(n_5183)
);

INVx2_ASAP7_75t_L g5184 ( 
.A(n_4650),
.Y(n_5184)
);

AOI22xp33_ASAP7_75t_L g5185 ( 
.A1(n_4725),
.A2(n_4169),
.B1(n_4498),
.B2(n_4034),
.Y(n_5185)
);

OAI21xp5_ASAP7_75t_L g5186 ( 
.A1(n_4902),
.A2(n_4720),
.B(n_4648),
.Y(n_5186)
);

AO31x2_ASAP7_75t_L g5187 ( 
.A1(n_4874),
.A2(n_4289),
.A3(n_4282),
.B(n_4294),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_4598),
.A2(n_4145),
.B(n_4018),
.Y(n_5188)
);

NAND2x1p5_ASAP7_75t_L g5189 ( 
.A(n_4624),
.B(n_4169),
.Y(n_5189)
);

OA21x2_ASAP7_75t_L g5190 ( 
.A1(n_4772),
.A2(n_4461),
.B(n_4455),
.Y(n_5190)
);

HB1xp67_ASAP7_75t_L g5191 ( 
.A(n_4846),
.Y(n_5191)
);

OR2x2_ASAP7_75t_L g5192 ( 
.A(n_4897),
.B(n_4424),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_4540),
.B(n_4253),
.Y(n_5193)
);

NAND2x1p5_ASAP7_75t_L g5194 ( 
.A(n_4624),
.B(n_4169),
.Y(n_5194)
);

INVx2_ASAP7_75t_SL g5195 ( 
.A(n_4792),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_4619),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4619),
.Y(n_5197)
);

A2O1A1Ixp33_ASAP7_75t_L g5198 ( 
.A1(n_4902),
.A2(n_4648),
.B(n_5001),
.C(n_4631),
.Y(n_5198)
);

INVx2_ASAP7_75t_L g5199 ( 
.A(n_4650),
.Y(n_5199)
);

NOR2xp67_ASAP7_75t_L g5200 ( 
.A(n_4541),
.B(n_4426),
.Y(n_5200)
);

AOI22xp33_ASAP7_75t_L g5201 ( 
.A1(n_4725),
.A2(n_4034),
.B1(n_4065),
.B2(n_4348),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_4620),
.Y(n_5202)
);

AOI22xp33_ASAP7_75t_L g5203 ( 
.A1(n_5001),
.A2(n_4127),
.B1(n_4277),
.B2(n_4348),
.Y(n_5203)
);

OAI21x1_ASAP7_75t_L g5204 ( 
.A1(n_4521),
.A2(n_4468),
.B(n_4461),
.Y(n_5204)
);

AND2x2_ASAP7_75t_L g5205 ( 
.A(n_4540),
.B(n_4053),
.Y(n_5205)
);

AO21x2_ASAP7_75t_L g5206 ( 
.A1(n_4888),
.A2(n_4468),
.B(n_4288),
.Y(n_5206)
);

OR2x2_ASAP7_75t_L g5207 ( 
.A(n_4919),
.B(n_4429),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_4620),
.Y(n_5208)
);

HB1xp67_ASAP7_75t_L g5209 ( 
.A(n_4846),
.Y(n_5209)
);

OR2x2_ASAP7_75t_L g5210 ( 
.A(n_4919),
.B(n_4258),
.Y(n_5210)
);

AND2x4_ASAP7_75t_L g5211 ( 
.A(n_4563),
.B(n_4397),
.Y(n_5211)
);

OAI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4720),
.A2(n_4485),
.B(n_4481),
.Y(n_5212)
);

AND2x4_ASAP7_75t_L g5213 ( 
.A(n_4563),
.B(n_4397),
.Y(n_5213)
);

A2O1A1Ixp33_ASAP7_75t_L g5214 ( 
.A1(n_4631),
.A2(n_4149),
.B(n_4157),
.C(n_4171),
.Y(n_5214)
);

AO21x2_ASAP7_75t_L g5215 ( 
.A1(n_4794),
.A2(n_4288),
.B(n_4515),
.Y(n_5215)
);

OR2x2_ASAP7_75t_L g5216 ( 
.A(n_4971),
.B(n_4264),
.Y(n_5216)
);

INVx1_ASAP7_75t_L g5217 ( 
.A(n_4643),
.Y(n_5217)
);

INVx2_ASAP7_75t_L g5218 ( 
.A(n_4650),
.Y(n_5218)
);

AND2x2_ASAP7_75t_L g5219 ( 
.A(n_4664),
.B(n_4053),
.Y(n_5219)
);

OR2x6_ASAP7_75t_L g5220 ( 
.A(n_4546),
.B(n_3993),
.Y(n_5220)
);

OAI21x1_ASAP7_75t_L g5221 ( 
.A1(n_4521),
.A2(n_3977),
.B(n_4491),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4643),
.Y(n_5222)
);

AOI21xp5_ASAP7_75t_L g5223 ( 
.A1(n_4645),
.A2(n_4145),
.B(n_4018),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_4616),
.B(n_4004),
.Y(n_5224)
);

INVx1_ASAP7_75t_L g5225 ( 
.A(n_4661),
.Y(n_5225)
);

INVx1_ASAP7_75t_L g5226 ( 
.A(n_4661),
.Y(n_5226)
);

INVx2_ASAP7_75t_L g5227 ( 
.A(n_4650),
.Y(n_5227)
);

OA21x2_ASAP7_75t_L g5228 ( 
.A1(n_4964),
.A2(n_4288),
.B(n_4504),
.Y(n_5228)
);

AND2x2_ASAP7_75t_L g5229 ( 
.A(n_4664),
.B(n_4255),
.Y(n_5229)
);

INVx4_ASAP7_75t_L g5230 ( 
.A(n_4644),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4575),
.B(n_4009),
.Y(n_5231)
);

OAI21x1_ASAP7_75t_L g5232 ( 
.A1(n_4883),
.A2(n_3977),
.B(n_4497),
.Y(n_5232)
);

HB1xp67_ASAP7_75t_L g5233 ( 
.A(n_4859),
.Y(n_5233)
);

OA21x2_ASAP7_75t_L g5234 ( 
.A1(n_4964),
.A2(n_4509),
.B(n_4474),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_4673),
.Y(n_5235)
);

OA21x2_ASAP7_75t_L g5236 ( 
.A1(n_4973),
.A2(n_4490),
.B(n_4471),
.Y(n_5236)
);

AOI21xp5_ASAP7_75t_L g5237 ( 
.A1(n_4645),
.A2(n_4145),
.B(n_4018),
.Y(n_5237)
);

AND2x2_ASAP7_75t_L g5238 ( 
.A(n_4664),
.B(n_4255),
.Y(n_5238)
);

NAND2xp5_ASAP7_75t_L g5239 ( 
.A(n_4575),
.B(n_4197),
.Y(n_5239)
);

OAI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_4571),
.A2(n_4485),
.B(n_4481),
.Y(n_5240)
);

OAI21x1_ASAP7_75t_L g5241 ( 
.A1(n_4883),
.A2(n_3977),
.B(n_4469),
.Y(n_5241)
);

OAI21x1_ASAP7_75t_SL g5242 ( 
.A1(n_4882),
.A2(n_4057),
.B(n_4056),
.Y(n_5242)
);

CKINVDCx5p33_ASAP7_75t_R g5243 ( 
.A(n_4644),
.Y(n_5243)
);

AOI211xp5_ASAP7_75t_L g5244 ( 
.A1(n_4527),
.A2(n_4225),
.B(n_4384),
.C(n_4220),
.Y(n_5244)
);

AOI21xp5_ASAP7_75t_L g5245 ( 
.A1(n_4695),
.A2(n_4145),
.B(n_4432),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_4708),
.B(n_4197),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_4673),
.Y(n_5247)
);

INVx2_ASAP7_75t_L g5248 ( 
.A(n_4650),
.Y(n_5248)
);

CKINVDCx11_ASAP7_75t_R g5249 ( 
.A(n_4644),
.Y(n_5249)
);

AND2x2_ASAP7_75t_L g5250 ( 
.A(n_4664),
.B(n_4332),
.Y(n_5250)
);

OAI21x1_ASAP7_75t_L g5251 ( 
.A1(n_4883),
.A2(n_3977),
.B(n_4469),
.Y(n_5251)
);

NOR2xp33_ASAP7_75t_L g5252 ( 
.A(n_4574),
.B(n_3993),
.Y(n_5252)
);

OAI21x1_ASAP7_75t_L g5253 ( 
.A1(n_4886),
.A2(n_4469),
.B(n_4513),
.Y(n_5253)
);

INVx2_ASAP7_75t_L g5254 ( 
.A(n_4524),
.Y(n_5254)
);

AO31x2_ASAP7_75t_L g5255 ( 
.A1(n_4998),
.A2(n_4519),
.A3(n_4518),
.B(n_4517),
.Y(n_5255)
);

INVx1_ASAP7_75t_L g5256 ( 
.A(n_4674),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_4886),
.A2(n_4469),
.B(n_4508),
.Y(n_5257)
);

AOI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_4861),
.A2(n_4397),
.B1(n_4212),
.B2(n_4199),
.Y(n_5258)
);

AOI22xp5_ASAP7_75t_L g5259 ( 
.A1(n_4861),
.A2(n_4397),
.B1(n_4085),
.B2(n_4074),
.Y(n_5259)
);

BUFx12f_ASAP7_75t_L g5260 ( 
.A(n_4892),
.Y(n_5260)
);

OAI21x1_ASAP7_75t_L g5261 ( 
.A1(n_4797),
.A2(n_4508),
.B(n_4343),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_4524),
.Y(n_5262)
);

AOI21xp5_ASAP7_75t_L g5263 ( 
.A1(n_4708),
.A2(n_4442),
.B(n_4120),
.Y(n_5263)
);

INVx2_ASAP7_75t_L g5264 ( 
.A(n_4524),
.Y(n_5264)
);

OAI21xp5_ASAP7_75t_L g5265 ( 
.A1(n_4777),
.A2(n_3968),
.B(n_3970),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_4674),
.Y(n_5266)
);

BUFx2_ASAP7_75t_L g5267 ( 
.A(n_4889),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_4693),
.Y(n_5268)
);

BUFx6f_ASAP7_75t_L g5269 ( 
.A(n_4624),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_4693),
.Y(n_5270)
);

AOI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_4940),
.A2(n_4454),
.B(n_4299),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_4859),
.B(n_4328),
.Y(n_5272)
);

INVx2_ASAP7_75t_SL g5273 ( 
.A(n_4669),
.Y(n_5273)
);

OA21x2_ASAP7_75t_L g5274 ( 
.A1(n_4973),
.A2(n_4515),
.B(n_4271),
.Y(n_5274)
);

INVx2_ASAP7_75t_L g5275 ( 
.A(n_4585),
.Y(n_5275)
);

OAI21x1_ASAP7_75t_L g5276 ( 
.A1(n_4797),
.A2(n_4450),
.B(n_4298),
.Y(n_5276)
);

OAI21xp5_ASAP7_75t_L g5277 ( 
.A1(n_4777),
.A2(n_4273),
.B(n_4278),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_4950),
.A2(n_4454),
.B(n_4295),
.Y(n_5278)
);

AND2x4_ASAP7_75t_L g5279 ( 
.A(n_4563),
.B(n_4127),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4697),
.Y(n_5280)
);

INVx6_ASAP7_75t_L g5281 ( 
.A(n_4656),
.Y(n_5281)
);

OAI21x1_ASAP7_75t_L g5282 ( 
.A1(n_4797),
.A2(n_4292),
.B(n_4257),
.Y(n_5282)
);

AOI21xp5_ASAP7_75t_L g5283 ( 
.A1(n_4950),
.A2(n_4454),
.B(n_4515),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4697),
.Y(n_5284)
);

OR2x6_ASAP7_75t_L g5285 ( 
.A(n_4636),
.B(n_3993),
.Y(n_5285)
);

O2A1O1Ixp33_ASAP7_75t_L g5286 ( 
.A1(n_4768),
.A2(n_4256),
.B(n_4254),
.C(n_4002),
.Y(n_5286)
);

HB1xp67_ASAP7_75t_L g5287 ( 
.A(n_4665),
.Y(n_5287)
);

NOR2xp33_ASAP7_75t_L g5288 ( 
.A(n_4557),
.B(n_3993),
.Y(n_5288)
);

AOI21xp5_ASAP7_75t_L g5289 ( 
.A1(n_4706),
.A2(n_4454),
.B(n_4515),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_4721),
.B(n_4191),
.Y(n_5290)
);

CKINVDCx6p67_ASAP7_75t_R g5291 ( 
.A(n_4761),
.Y(n_5291)
);

HB1xp67_ASAP7_75t_L g5292 ( 
.A(n_4665),
.Y(n_5292)
);

OA21x2_ASAP7_75t_L g5293 ( 
.A1(n_4973),
.A2(n_4271),
.B(n_3989),
.Y(n_5293)
);

OAI21x1_ASAP7_75t_L g5294 ( 
.A1(n_4652),
.A2(n_4124),
.B(n_4141),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_4698),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_4698),
.Y(n_5296)
);

AND2x4_ASAP7_75t_L g5297 ( 
.A(n_4563),
.B(n_4127),
.Y(n_5297)
);

NAND2xp5_ASAP7_75t_L g5298 ( 
.A(n_4710),
.B(n_4242),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_4700),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4706),
.A2(n_4125),
.B(n_4161),
.Y(n_5300)
);

BUFx6f_ASAP7_75t_L g5301 ( 
.A(n_4624),
.Y(n_5301)
);

INVx2_ASAP7_75t_L g5302 ( 
.A(n_4585),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_4710),
.B(n_3946),
.Y(n_5303)
);

BUFx8_ASAP7_75t_L g5304 ( 
.A(n_4761),
.Y(n_5304)
);

INVx3_ASAP7_75t_L g5305 ( 
.A(n_4920),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_4682),
.A2(n_4143),
.B(n_4158),
.Y(n_5306)
);

AO31x2_ASAP7_75t_L g5307 ( 
.A1(n_5010),
.A2(n_4189),
.A3(n_4160),
.B(n_4063),
.Y(n_5307)
);

OAI21x1_ASAP7_75t_L g5308 ( 
.A1(n_4652),
.A2(n_4195),
.B(n_4192),
.Y(n_5308)
);

AO21x2_ASAP7_75t_L g5309 ( 
.A1(n_4754),
.A2(n_4686),
.B(n_4745),
.Y(n_5309)
);

INVx3_ASAP7_75t_L g5310 ( 
.A(n_4920),
.Y(n_5310)
);

BUFx12f_ASAP7_75t_L g5311 ( 
.A(n_4744),
.Y(n_5311)
);

NAND2x1p5_ASAP7_75t_L g5312 ( 
.A(n_4739),
.B(n_4252),
.Y(n_5312)
);

OAI21x1_ASAP7_75t_L g5313 ( 
.A1(n_4652),
.A2(n_4332),
.B(n_4418),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_4700),
.Y(n_5314)
);

OA21x2_ASAP7_75t_L g5315 ( 
.A1(n_4947),
.A2(n_4271),
.B(n_4160),
.Y(n_5315)
);

OA21x2_ASAP7_75t_L g5316 ( 
.A1(n_4947),
.A2(n_4271),
.B(n_4160),
.Y(n_5316)
);

INVx1_ASAP7_75t_L g5317 ( 
.A(n_4701),
.Y(n_5317)
);

NAND2xp5_ASAP7_75t_SL g5318 ( 
.A(n_4528),
.B(n_4074),
.Y(n_5318)
);

BUFx4f_ASAP7_75t_SL g5319 ( 
.A(n_4713),
.Y(n_5319)
);

INVx2_ASAP7_75t_L g5320 ( 
.A(n_4585),
.Y(n_5320)
);

INVx4_ASAP7_75t_L g5321 ( 
.A(n_4656),
.Y(n_5321)
);

AO21x2_ASAP7_75t_L g5322 ( 
.A1(n_4754),
.A2(n_4271),
.B(n_4189),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_4701),
.Y(n_5323)
);

AND2x2_ASAP7_75t_L g5324 ( 
.A(n_4872),
.B(n_4418),
.Y(n_5324)
);

OAI21x1_ASAP7_75t_L g5325 ( 
.A1(n_4651),
.A2(n_4063),
.B(n_4434),
.Y(n_5325)
);

OAI21x1_ASAP7_75t_L g5326 ( 
.A1(n_4651),
.A2(n_4063),
.B(n_4434),
.Y(n_5326)
);

INVx2_ASAP7_75t_SL g5327 ( 
.A(n_4669),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_4826),
.B(n_4862),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_4826),
.B(n_3946),
.Y(n_5329)
);

OA21x2_ASAP7_75t_L g5330 ( 
.A1(n_4947),
.A2(n_4160),
.B(n_4189),
.Y(n_5330)
);

A2O1A1Ixp33_ASAP7_75t_L g5331 ( 
.A1(n_4834),
.A2(n_4277),
.B(n_4348),
.C(n_4252),
.Y(n_5331)
);

AO21x2_ASAP7_75t_L g5332 ( 
.A1(n_4686),
.A2(n_4189),
.B(n_4160),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_4702),
.Y(n_5333)
);

OA21x2_ASAP7_75t_L g5334 ( 
.A1(n_4949),
.A2(n_4189),
.B(n_4063),
.Y(n_5334)
);

OAI21x1_ASAP7_75t_L g5335 ( 
.A1(n_4651),
.A2(n_4063),
.B(n_4070),
.Y(n_5335)
);

INVx1_ASAP7_75t_L g5336 ( 
.A(n_4702),
.Y(n_5336)
);

AOI21xp5_ASAP7_75t_L g5337 ( 
.A1(n_4945),
.A2(n_4252),
.B(n_4277),
.Y(n_5337)
);

INVx1_ASAP7_75t_L g5338 ( 
.A(n_4737),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_4737),
.Y(n_5339)
);

BUFx3_ASAP7_75t_L g5340 ( 
.A(n_4761),
.Y(n_5340)
);

INVx1_ASAP7_75t_L g5341 ( 
.A(n_4756),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_4862),
.B(n_3806),
.Y(n_5342)
);

AOI21x1_ASAP7_75t_L g5343 ( 
.A1(n_4825),
.A2(n_3981),
.B(n_4340),
.Y(n_5343)
);

OAI21x1_ASAP7_75t_L g5344 ( 
.A1(n_4981),
.A2(n_4005),
.B(n_4121),
.Y(n_5344)
);

INVx2_ASAP7_75t_L g5345 ( 
.A(n_4610),
.Y(n_5345)
);

INVx1_ASAP7_75t_L g5346 ( 
.A(n_4756),
.Y(n_5346)
);

INVx2_ASAP7_75t_L g5347 ( 
.A(n_4610),
.Y(n_5347)
);

AND2x2_ASAP7_75t_L g5348 ( 
.A(n_4872),
.B(n_4005),
.Y(n_5348)
);

INVx2_ASAP7_75t_SL g5349 ( 
.A(n_4669),
.Y(n_5349)
);

AOI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_4945),
.A2(n_4247),
.B(n_4129),
.Y(n_5350)
);

AND2x4_ASAP7_75t_L g5351 ( 
.A(n_4600),
.B(n_4074),
.Y(n_5351)
);

AO31x2_ASAP7_75t_L g5352 ( 
.A1(n_5010),
.A2(n_4005),
.A3(n_4213),
.B(n_3979),
.Y(n_5352)
);

AOI21xp5_ASAP7_75t_L g5353 ( 
.A1(n_4689),
.A2(n_4247),
.B(n_4129),
.Y(n_5353)
);

NOR2x1_ASAP7_75t_SL g5354 ( 
.A(n_4555),
.B(n_4074),
.Y(n_5354)
);

AOI21xp5_ASAP7_75t_L g5355 ( 
.A1(n_4738),
.A2(n_4247),
.B(n_4129),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_4738),
.A2(n_4247),
.B(n_4129),
.Y(n_5356)
);

NAND2xp5_ASAP7_75t_L g5357 ( 
.A(n_4876),
.B(n_3806),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_4760),
.Y(n_5358)
);

INVx3_ASAP7_75t_L g5359 ( 
.A(n_4920),
.Y(n_5359)
);

BUFx2_ASAP7_75t_R g5360 ( 
.A(n_4591),
.Y(n_5360)
);

OA21x2_ASAP7_75t_L g5361 ( 
.A1(n_4949),
.A2(n_4260),
.B(n_4266),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_L g5362 ( 
.A(n_4876),
.B(n_3806),
.Y(n_5362)
);

OA21x2_ASAP7_75t_L g5363 ( 
.A1(n_4949),
.A2(n_4958),
.B(n_4968),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_4738),
.A2(n_4247),
.B(n_4129),
.Y(n_5364)
);

OAI21x1_ASAP7_75t_SL g5365 ( 
.A1(n_4871),
.A2(n_4005),
.B(n_3979),
.Y(n_5365)
);

NAND3xp33_ASAP7_75t_SL g5366 ( 
.A(n_4655),
.B(n_4005),
.C(n_4364),
.Y(n_5366)
);

AND2x2_ASAP7_75t_L g5367 ( 
.A(n_4872),
.B(n_4696),
.Y(n_5367)
);

AND2x4_ASAP7_75t_L g5368 ( 
.A(n_4600),
.B(n_4623),
.Y(n_5368)
);

AOI21xp5_ASAP7_75t_L g5369 ( 
.A1(n_4738),
.A2(n_4425),
.B(n_4395),
.Y(n_5369)
);

AOI221xp5_ASAP7_75t_L g5370 ( 
.A1(n_4552),
.A2(n_4085),
.B1(n_4074),
.B2(n_4317),
.C(n_4395),
.Y(n_5370)
);

AOI21xp5_ASAP7_75t_L g5371 ( 
.A1(n_4796),
.A2(n_4425),
.B(n_4395),
.Y(n_5371)
);

AOI21xp5_ASAP7_75t_L g5372 ( 
.A1(n_4796),
.A2(n_4425),
.B(n_4395),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_4760),
.Y(n_5373)
);

INVx2_ASAP7_75t_L g5374 ( 
.A(n_4610),
.Y(n_5374)
);

NAND2xp5_ASAP7_75t_L g5375 ( 
.A(n_4879),
.B(n_3806),
.Y(n_5375)
);

OAI21xp5_ASAP7_75t_L g5376 ( 
.A1(n_4582),
.A2(n_2810),
.B(n_4293),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_4763),
.Y(n_5377)
);

NOR2xp33_ASAP7_75t_L g5378 ( 
.A(n_4626),
.B(n_4085),
.Y(n_5378)
);

AND2x4_ASAP7_75t_L g5379 ( 
.A(n_4600),
.B(n_4085),
.Y(n_5379)
);

HB1xp67_ASAP7_75t_L g5380 ( 
.A(n_4692),
.Y(n_5380)
);

AOI21xp5_ASAP7_75t_L g5381 ( 
.A1(n_4743),
.A2(n_4942),
.B(n_4642),
.Y(n_5381)
);

INVx1_ASAP7_75t_L g5382 ( 
.A(n_4763),
.Y(n_5382)
);

AOI21xp33_ASAP7_75t_SL g5383 ( 
.A1(n_4669),
.A2(n_4395),
.B(n_4317),
.Y(n_5383)
);

AND2x2_ASAP7_75t_L g5384 ( 
.A(n_4872),
.B(n_4262),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4770),
.Y(n_5385)
);

AOI21xp5_ASAP7_75t_L g5386 ( 
.A1(n_4942),
.A2(n_4425),
.B(n_4317),
.Y(n_5386)
);

AOI21xp5_ASAP7_75t_L g5387 ( 
.A1(n_4642),
.A2(n_4425),
.B(n_4317),
.Y(n_5387)
);

AOI221xp5_ASAP7_75t_L g5388 ( 
.A1(n_4768),
.A2(n_4085),
.B1(n_4317),
.B2(n_4501),
.C(n_4493),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_4770),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_4771),
.Y(n_5390)
);

OR2x6_ASAP7_75t_L g5391 ( 
.A(n_4636),
.B(n_2419),
.Y(n_5391)
);

OAI21x1_ASAP7_75t_SL g5392 ( 
.A1(n_4871),
.A2(n_4311),
.B(n_4262),
.Y(n_5392)
);

NAND2xp5_ASAP7_75t_L g5393 ( 
.A(n_4879),
.B(n_3806),
.Y(n_5393)
);

OR2x2_ASAP7_75t_L g5394 ( 
.A(n_4971),
.B(n_4293),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_4771),
.Y(n_5395)
);

INVx1_ASAP7_75t_L g5396 ( 
.A(n_4783),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_4783),
.Y(n_5397)
);

NAND2xp5_ASAP7_75t_L g5398 ( 
.A(n_4818),
.B(n_3806),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_4818),
.B(n_4337),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_4613),
.Y(n_5400)
);

INVx3_ASAP7_75t_L g5401 ( 
.A(n_4911),
.Y(n_5401)
);

BUFx2_ASAP7_75t_L g5402 ( 
.A(n_4889),
.Y(n_5402)
);

AOI21x1_ASAP7_75t_L g5403 ( 
.A1(n_4930),
.A2(n_4311),
.B(n_4291),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_4787),
.Y(n_5404)
);

AOI21xp5_ASAP7_75t_L g5405 ( 
.A1(n_4989),
.A2(n_2464),
.B(n_2466),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_4787),
.Y(n_5406)
);

OR2x2_ASAP7_75t_L g5407 ( 
.A(n_4692),
.B(n_4293),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_4790),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_4790),
.Y(n_5409)
);

AND2x4_ASAP7_75t_SL g5410 ( 
.A(n_4994),
.B(n_4291),
.Y(n_5410)
);

AND2x4_ASAP7_75t_L g5411 ( 
.A(n_4600),
.B(n_4337),
.Y(n_5411)
);

AOI21x1_ASAP7_75t_L g5412 ( 
.A1(n_4930),
.A2(n_4311),
.B(n_4291),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_4793),
.Y(n_5413)
);

INVx8_ASAP7_75t_L g5414 ( 
.A(n_4534),
.Y(n_5414)
);

NAND2xp5_ASAP7_75t_L g5415 ( 
.A(n_4678),
.B(n_4679),
.Y(n_5415)
);

OAI21x1_ASAP7_75t_L g5416 ( 
.A1(n_4981),
.A2(n_4121),
.B(n_4135),
.Y(n_5416)
);

AND2x2_ASAP7_75t_L g5417 ( 
.A(n_4696),
.B(n_4291),
.Y(n_5417)
);

OR2x2_ASAP7_75t_L g5418 ( 
.A(n_4705),
.B(n_4293),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_4793),
.Y(n_5419)
);

OAI21x1_ASAP7_75t_L g5420 ( 
.A1(n_4981),
.A2(n_4121),
.B(n_4135),
.Y(n_5420)
);

NAND2xp5_ASAP7_75t_L g5421 ( 
.A(n_4679),
.B(n_4337),
.Y(n_5421)
);

BUFx2_ASAP7_75t_L g5422 ( 
.A(n_4555),
.Y(n_5422)
);

OR2x6_ASAP7_75t_L g5423 ( 
.A(n_4555),
.B(n_2464),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_4613),
.Y(n_5424)
);

OR2x2_ASAP7_75t_L g5425 ( 
.A(n_4705),
.B(n_4293),
.Y(n_5425)
);

CKINVDCx5p33_ASAP7_75t_R g5426 ( 
.A(n_4936),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_4613),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_4800),
.Y(n_5428)
);

A2O1A1Ixp33_ASAP7_75t_L g5429 ( 
.A1(n_4849),
.A2(n_4655),
.B(n_4614),
.C(n_4819),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_4800),
.Y(n_5430)
);

HB1xp67_ASAP7_75t_L g5431 ( 
.A(n_4812),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_4812),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_4816),
.Y(n_5433)
);

INVx1_ASAP7_75t_L g5434 ( 
.A(n_4816),
.Y(n_5434)
);

INVx1_ASAP7_75t_L g5435 ( 
.A(n_4829),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_4829),
.Y(n_5436)
);

BUFx8_ASAP7_75t_SL g5437 ( 
.A(n_4639),
.Y(n_5437)
);

OAI21xp5_ASAP7_75t_L g5438 ( 
.A1(n_4582),
.A2(n_4666),
.B(n_4628),
.Y(n_5438)
);

BUFx6f_ASAP7_75t_L g5439 ( 
.A(n_4639),
.Y(n_5439)
);

INVx2_ASAP7_75t_SL g5440 ( 
.A(n_4669),
.Y(n_5440)
);

HB1xp67_ASAP7_75t_L g5441 ( 
.A(n_4844),
.Y(n_5441)
);

INVx1_ASAP7_75t_L g5442 ( 
.A(n_4844),
.Y(n_5442)
);

BUFx2_ASAP7_75t_L g5443 ( 
.A(n_4555),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_4751),
.B(n_4337),
.Y(n_5444)
);

NAND2xp5_ASAP7_75t_L g5445 ( 
.A(n_4751),
.B(n_4337),
.Y(n_5445)
);

INVx3_ASAP7_75t_L g5446 ( 
.A(n_4638),
.Y(n_5446)
);

A2O1A1Ixp33_ASAP7_75t_L g5447 ( 
.A1(n_4849),
.A2(n_4501),
.B(n_4493),
.C(n_4311),
.Y(n_5447)
);

NAND2xp5_ASAP7_75t_L g5448 ( 
.A(n_4820),
.B(n_4400),
.Y(n_5448)
);

CKINVDCx11_ASAP7_75t_R g5449 ( 
.A(n_4656),
.Y(n_5449)
);

NOR2xp33_ASAP7_75t_L g5450 ( 
.A(n_4639),
.B(n_4340),
.Y(n_5450)
);

INVx2_ASAP7_75t_SL g5451 ( 
.A(n_4669),
.Y(n_5451)
);

BUFx6f_ASAP7_75t_L g5452 ( 
.A(n_4716),
.Y(n_5452)
);

OR2x2_ASAP7_75t_L g5453 ( 
.A(n_4948),
.B(n_4501),
.Y(n_5453)
);

INVx1_ASAP7_75t_L g5454 ( 
.A(n_4847),
.Y(n_5454)
);

A2O1A1Ixp33_ASAP7_75t_L g5455 ( 
.A1(n_4614),
.A2(n_4501),
.B(n_4493),
.C(n_4340),
.Y(n_5455)
);

OA21x2_ASAP7_75t_L g5456 ( 
.A1(n_4958),
.A2(n_4260),
.B(n_4266),
.Y(n_5456)
);

AOI21xp5_ASAP7_75t_SL g5457 ( 
.A1(n_4869),
.A2(n_2464),
.B(n_2466),
.Y(n_5457)
);

BUFx12f_ASAP7_75t_L g5458 ( 
.A(n_4568),
.Y(n_5458)
);

OR2x2_ASAP7_75t_L g5459 ( 
.A(n_4948),
.B(n_4501),
.Y(n_5459)
);

AO21x2_ASAP7_75t_L g5460 ( 
.A1(n_4745),
.A2(n_4213),
.B(n_4266),
.Y(n_5460)
);

AOI22xp33_ASAP7_75t_L g5461 ( 
.A1(n_4584),
.A2(n_4340),
.B1(n_4364),
.B2(n_4389),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4847),
.Y(n_5462)
);

AOI21xp33_ASAP7_75t_SL g5463 ( 
.A1(n_4534),
.A2(n_4364),
.B(n_4389),
.Y(n_5463)
);

INVx1_ASAP7_75t_L g5464 ( 
.A(n_4850),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_4850),
.Y(n_5465)
);

NAND2xp5_ASAP7_75t_L g5466 ( 
.A(n_4820),
.B(n_4400),
.Y(n_5466)
);

NAND2xp5_ASAP7_75t_L g5467 ( 
.A(n_4736),
.B(n_4400),
.Y(n_5467)
);

AOI21x1_ASAP7_75t_L g5468 ( 
.A1(n_4660),
.A2(n_4389),
.B(n_4364),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_4630),
.Y(n_5469)
);

NAND2xp5_ASAP7_75t_L g5470 ( 
.A(n_4819),
.B(n_4400),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_4630),
.Y(n_5471)
);

NAND2xp5_ASAP7_75t_L g5472 ( 
.A(n_4837),
.B(n_4727),
.Y(n_5472)
);

INVx2_ASAP7_75t_L g5473 ( 
.A(n_4630),
.Y(n_5473)
);

INVx1_ASAP7_75t_L g5474 ( 
.A(n_4853),
.Y(n_5474)
);

AO21x2_ASAP7_75t_L g5475 ( 
.A1(n_4685),
.A2(n_4213),
.B(n_4260),
.Y(n_5475)
);

OAI21xp5_ASAP7_75t_L g5476 ( 
.A1(n_4681),
.A2(n_4765),
.B(n_4654),
.Y(n_5476)
);

AOI21xp5_ASAP7_75t_L g5477 ( 
.A1(n_4989),
.A2(n_2466),
.B(n_2501),
.Y(n_5477)
);

BUFx2_ASAP7_75t_L g5478 ( 
.A(n_4555),
.Y(n_5478)
);

INVx1_ASAP7_75t_SL g5479 ( 
.A(n_4961),
.Y(n_5479)
);

OAI21x1_ASAP7_75t_L g5480 ( 
.A1(n_4997),
.A2(n_4986),
.B(n_4806),
.Y(n_5480)
);

BUFx3_ASAP7_75t_L g5481 ( 
.A(n_4534),
.Y(n_5481)
);

NAND2x1p5_ASAP7_75t_L g5482 ( 
.A(n_4739),
.B(n_2466),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_4853),
.Y(n_5483)
);

OA21x2_ASAP7_75t_L g5484 ( 
.A1(n_4958),
.A2(n_4260),
.B(n_4266),
.Y(n_5484)
);

AOI22xp33_ASAP7_75t_L g5485 ( 
.A1(n_4554),
.A2(n_4389),
.B1(n_2810),
.B2(n_2536),
.Y(n_5485)
);

AOI21x1_ASAP7_75t_L g5486 ( 
.A1(n_4660),
.A2(n_4266),
.B(n_4260),
.Y(n_5486)
);

OAI21x1_ASAP7_75t_L g5487 ( 
.A1(n_4997),
.A2(n_4151),
.B(n_4121),
.Y(n_5487)
);

OAI21xp5_ASAP7_75t_L g5488 ( 
.A1(n_4654),
.A2(n_2810),
.B(n_4493),
.Y(n_5488)
);

NAND2xp5_ASAP7_75t_L g5489 ( 
.A(n_4727),
.B(n_4400),
.Y(n_5489)
);

NOR2xp67_ASAP7_75t_R g5490 ( 
.A(n_4568),
.B(n_2466),
.Y(n_5490)
);

OAI21xp5_ASAP7_75t_L g5491 ( 
.A1(n_4654),
.A2(n_2810),
.B(n_4493),
.Y(n_5491)
);

OAI21x1_ASAP7_75t_L g5492 ( 
.A1(n_4997),
.A2(n_4176),
.B(n_4151),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_4632),
.Y(n_5493)
);

HB1xp67_ASAP7_75t_L g5494 ( 
.A(n_4867),
.Y(n_5494)
);

INVx2_ASAP7_75t_L g5495 ( 
.A(n_4632),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_4867),
.Y(n_5496)
);

NAND2xp5_ASAP7_75t_L g5497 ( 
.A(n_4730),
.B(n_3737),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_4870),
.Y(n_5498)
);

NAND2xp5_ASAP7_75t_L g5499 ( 
.A(n_4730),
.B(n_4750),
.Y(n_5499)
);

AOI21x1_ASAP7_75t_L g5500 ( 
.A1(n_4711),
.A2(n_4272),
.B(n_4283),
.Y(n_5500)
);

AOI221xp5_ASAP7_75t_L g5501 ( 
.A1(n_4752),
.A2(n_4460),
.B1(n_4451),
.B2(n_4445),
.C(n_4440),
.Y(n_5501)
);

AO21x2_ASAP7_75t_L g5502 ( 
.A1(n_4685),
.A2(n_4272),
.B(n_4451),
.Y(n_5502)
);

AOI21xp5_ASAP7_75t_L g5503 ( 
.A1(n_4694),
.A2(n_2466),
.B(n_2501),
.Y(n_5503)
);

OA21x2_ASAP7_75t_L g5504 ( 
.A1(n_4968),
.A2(n_4272),
.B(n_4283),
.Y(n_5504)
);

NAND2xp5_ASAP7_75t_L g5505 ( 
.A(n_4730),
.B(n_3737),
.Y(n_5505)
);

OAI22xp5_ASAP7_75t_L g5506 ( 
.A1(n_4688),
.A2(n_2466),
.B1(n_2501),
.B2(n_2536),
.Y(n_5506)
);

INVx1_ASAP7_75t_SL g5507 ( 
.A(n_4961),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_4750),
.B(n_3706),
.Y(n_5508)
);

NAND2xp5_ASAP7_75t_L g5509 ( 
.A(n_4750),
.B(n_3706),
.Y(n_5509)
);

HB1xp67_ASAP7_75t_L g5510 ( 
.A(n_4870),
.Y(n_5510)
);

INVx2_ASAP7_75t_L g5511 ( 
.A(n_4632),
.Y(n_5511)
);

NAND2xp5_ASAP7_75t_SL g5512 ( 
.A(n_4528),
.B(n_2466),
.Y(n_5512)
);

AOI21xp5_ASAP7_75t_L g5513 ( 
.A1(n_4717),
.A2(n_4943),
.B(n_4903),
.Y(n_5513)
);

OA21x2_ASAP7_75t_L g5514 ( 
.A1(n_4968),
.A2(n_4272),
.B(n_4283),
.Y(n_5514)
);

AND2x2_ASAP7_75t_L g5515 ( 
.A(n_4731),
.B(n_4324),
.Y(n_5515)
);

OAI21x1_ASAP7_75t_L g5516 ( 
.A1(n_4986),
.A2(n_4176),
.B(n_4151),
.Y(n_5516)
);

AO21x2_ASAP7_75t_L g5517 ( 
.A1(n_4685),
.A2(n_4272),
.B(n_4445),
.Y(n_5517)
);

OAI21x1_ASAP7_75t_L g5518 ( 
.A1(n_4986),
.A2(n_4151),
.B(n_4176),
.Y(n_5518)
);

AO21x2_ASAP7_75t_L g5519 ( 
.A1(n_4685),
.A2(n_4460),
.B(n_4445),
.Y(n_5519)
);

AND2x6_ASAP7_75t_L g5520 ( 
.A(n_4716),
.B(n_2501),
.Y(n_5520)
);

AOI21xp5_ASAP7_75t_L g5521 ( 
.A1(n_4903),
.A2(n_2501),
.B(n_2536),
.Y(n_5521)
);

AOI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_4943),
.A2(n_2501),
.B(n_2536),
.Y(n_5522)
);

OAI21x1_ASAP7_75t_L g5523 ( 
.A1(n_4986),
.A2(n_4151),
.B(n_4176),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_4757),
.B(n_3706),
.Y(n_5524)
);

NAND2xp5_ASAP7_75t_L g5525 ( 
.A(n_4757),
.B(n_3706),
.Y(n_5525)
);

OR2x6_ASAP7_75t_L g5526 ( 
.A(n_4555),
.B(n_2501),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_4634),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_4878),
.Y(n_5528)
);

INVx2_ASAP7_75t_L g5529 ( 
.A(n_4634),
.Y(n_5529)
);

INVx2_ASAP7_75t_SL g5530 ( 
.A(n_4993),
.Y(n_5530)
);

AOI22xp5_ASAP7_75t_L g5531 ( 
.A1(n_4895),
.A2(n_2501),
.B1(n_2536),
.B2(n_2540),
.Y(n_5531)
);

AO21x2_ASAP7_75t_L g5532 ( 
.A1(n_4699),
.A2(n_4445),
.B(n_4440),
.Y(n_5532)
);

OR2x2_ASAP7_75t_L g5533 ( 
.A(n_4801),
.B(n_4440),
.Y(n_5533)
);

NAND2xp5_ASAP7_75t_L g5534 ( 
.A(n_4757),
.B(n_3706),
.Y(n_5534)
);

OAI21x1_ASAP7_75t_L g5535 ( 
.A1(n_4788),
.A2(n_4135),
.B(n_4121),
.Y(n_5535)
);

AO21x2_ASAP7_75t_L g5536 ( 
.A1(n_4699),
.A2(n_4440),
.B(n_4437),
.Y(n_5536)
);

OR2x2_ASAP7_75t_L g5537 ( 
.A(n_4801),
.B(n_4440),
.Y(n_5537)
);

NOR2x1_ASAP7_75t_SL g5538 ( 
.A(n_4638),
.B(n_4135),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_L g5539 ( 
.A(n_4782),
.B(n_3787),
.Y(n_5539)
);

INVxp67_ASAP7_75t_SL g5540 ( 
.A(n_4927),
.Y(n_5540)
);

AOI21xp5_ASAP7_75t_L g5541 ( 
.A1(n_5007),
.A2(n_2536),
.B(n_2540),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_4782),
.B(n_3787),
.Y(n_5542)
);

BUFx2_ASAP7_75t_L g5543 ( 
.A(n_4712),
.Y(n_5543)
);

AND2x4_ASAP7_75t_L g5544 ( 
.A(n_4623),
.B(n_4330),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_4878),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_L g5546 ( 
.A(n_4782),
.B(n_3787),
.Y(n_5546)
);

INVx3_ASAP7_75t_L g5547 ( 
.A(n_4638),
.Y(n_5547)
);

AOI21xp5_ASAP7_75t_L g5548 ( 
.A1(n_5007),
.A2(n_2536),
.B(n_2540),
.Y(n_5548)
);

AOI21x1_ASAP7_75t_L g5549 ( 
.A1(n_4711),
.A2(n_4283),
.B(n_4330),
.Y(n_5549)
);

AOI21xp5_ASAP7_75t_L g5550 ( 
.A1(n_4817),
.A2(n_2536),
.B(n_2540),
.Y(n_5550)
);

INVx1_ASAP7_75t_L g5551 ( 
.A(n_4884),
.Y(n_5551)
);

NAND2xp5_ASAP7_75t_L g5552 ( 
.A(n_4838),
.B(n_3787),
.Y(n_5552)
);

OA21x2_ASAP7_75t_L g5553 ( 
.A1(n_4939),
.A2(n_5011),
.B(n_5008),
.Y(n_5553)
);

AOI22xp33_ASAP7_75t_L g5554 ( 
.A1(n_4802),
.A2(n_2540),
.B1(n_2549),
.B2(n_2551),
.Y(n_5554)
);

OAI21x1_ASAP7_75t_L g5555 ( 
.A1(n_4806),
.A2(n_4690),
.B(n_4602),
.Y(n_5555)
);

OAI21x1_ASAP7_75t_L g5556 ( 
.A1(n_4690),
.A2(n_4330),
.B(n_4324),
.Y(n_5556)
);

OR2x2_ASAP7_75t_L g5557 ( 
.A(n_4842),
.B(n_4437),
.Y(n_5557)
);

AOI21x1_ASAP7_75t_L g5558 ( 
.A1(n_4854),
.A2(n_4753),
.B(n_4746),
.Y(n_5558)
);

NAND2xp5_ASAP7_75t_L g5559 ( 
.A(n_4838),
.B(n_3787),
.Y(n_5559)
);

INVx2_ASAP7_75t_L g5560 ( 
.A(n_5079),
.Y(n_5560)
);

CKINVDCx5p33_ASAP7_75t_R g5561 ( 
.A(n_5249),
.Y(n_5561)
);

NAND2xp5_ASAP7_75t_L g5562 ( 
.A(n_5092),
.B(n_4838),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_5431),
.Y(n_5563)
);

BUFx2_ASAP7_75t_L g5564 ( 
.A(n_5321),
.Y(n_5564)
);

AOI22xp33_ASAP7_75t_SL g5565 ( 
.A1(n_5186),
.A2(n_4739),
.B1(n_4677),
.B2(n_4638),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_5075),
.A2(n_4972),
.B1(n_4832),
.B2(n_4573),
.Y(n_5566)
);

AOI211xp5_ASAP7_75t_L g5567 ( 
.A1(n_5198),
.A2(n_4845),
.B(n_4836),
.C(n_4960),
.Y(n_5567)
);

OAI21xp5_ASAP7_75t_SL g5568 ( 
.A1(n_5176),
.A2(n_4604),
.B(n_4590),
.Y(n_5568)
);

BUFx3_ASAP7_75t_L g5569 ( 
.A(n_5055),
.Y(n_5569)
);

AOI22xp33_ASAP7_75t_SL g5570 ( 
.A1(n_5476),
.A2(n_4739),
.B1(n_4677),
.B2(n_4638),
.Y(n_5570)
);

AOI22xp33_ASAP7_75t_L g5571 ( 
.A1(n_5077),
.A2(n_4972),
.B1(n_4832),
.B2(n_4577),
.Y(n_5571)
);

INVx1_ASAP7_75t_L g5572 ( 
.A(n_5023),
.Y(n_5572)
);

OAI22xp5_ASAP7_75t_L g5573 ( 
.A1(n_5429),
.A2(n_4604),
.B1(n_4688),
.B2(n_4822),
.Y(n_5573)
);

AOI22xp33_ASAP7_75t_L g5574 ( 
.A1(n_5053),
.A2(n_4817),
.B1(n_4802),
.B2(n_4719),
.Y(n_5574)
);

INVx3_ASAP7_75t_L g5575 ( 
.A(n_5150),
.Y(n_5575)
);

AOI22xp33_ASAP7_75t_SL g5576 ( 
.A1(n_5122),
.A2(n_4739),
.B1(n_4677),
.B2(n_4638),
.Y(n_5576)
);

INVx2_ASAP7_75t_L g5577 ( 
.A(n_5079),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_5023),
.Y(n_5578)
);

INVx3_ASAP7_75t_L g5579 ( 
.A(n_5150),
.Y(n_5579)
);

NAND2xp5_ASAP7_75t_L g5580 ( 
.A(n_5178),
.B(n_4840),
.Y(n_5580)
);

CKINVDCx11_ASAP7_75t_R g5581 ( 
.A(n_5055),
.Y(n_5581)
);

CKINVDCx5p33_ASAP7_75t_R g5582 ( 
.A(n_5260),
.Y(n_5582)
);

AOI22xp33_ASAP7_75t_L g5583 ( 
.A1(n_5141),
.A2(n_4817),
.B1(n_4752),
.B2(n_4778),
.Y(n_5583)
);

INVx2_ASAP7_75t_L g5584 ( 
.A(n_5079),
.Y(n_5584)
);

OAI22xp5_ASAP7_75t_L g5585 ( 
.A1(n_5168),
.A2(n_5062),
.B1(n_5059),
.B2(n_5123),
.Y(n_5585)
);

OAI222xp33_ASAP7_75t_L g5586 ( 
.A1(n_5381),
.A2(n_4895),
.B1(n_4836),
.B2(n_4863),
.C1(n_4842),
.C2(n_4905),
.Y(n_5586)
);

OAI22xp5_ASAP7_75t_L g5587 ( 
.A1(n_5168),
.A2(n_5331),
.B1(n_5472),
.B2(n_5076),
.Y(n_5587)
);

AOI22xp33_ASAP7_75t_L g5588 ( 
.A1(n_5032),
.A2(n_4817),
.B1(n_4677),
.B2(n_4638),
.Y(n_5588)
);

AOI22xp33_ASAP7_75t_L g5589 ( 
.A1(n_5041),
.A2(n_4677),
.B1(n_4733),
.B2(n_4621),
.Y(n_5589)
);

CKINVDCx20_ASAP7_75t_R g5590 ( 
.A(n_5129),
.Y(n_5590)
);

OAI211xp5_ASAP7_75t_SL g5591 ( 
.A1(n_5028),
.A2(n_4845),
.B(n_4900),
.C(n_4918),
.Y(n_5591)
);

OAI21xp33_ASAP7_75t_L g5592 ( 
.A1(n_5115),
.A2(n_4905),
.B(n_4969),
.Y(n_5592)
);

INVx3_ASAP7_75t_L g5593 ( 
.A(n_5164),
.Y(n_5593)
);

AND2x2_ASAP7_75t_L g5594 ( 
.A(n_5016),
.B(n_4731),
.Y(n_5594)
);

AOI22xp5_ASAP7_75t_L g5595 ( 
.A1(n_5071),
.A2(n_4875),
.B1(n_4858),
.B2(n_4956),
.Y(n_5595)
);

INVx2_ASAP7_75t_L g5596 ( 
.A(n_5079),
.Y(n_5596)
);

OAI22xp5_ASAP7_75t_L g5597 ( 
.A1(n_5201),
.A2(n_4906),
.B1(n_4803),
.B2(n_4805),
.Y(n_5597)
);

AOI22xp5_ASAP7_75t_L g5598 ( 
.A1(n_5117),
.A2(n_4956),
.B1(n_4749),
.B2(n_4906),
.Y(n_5598)
);

OAI21xp33_ASAP7_75t_L g5599 ( 
.A1(n_5142),
.A2(n_4969),
.B(n_4830),
.Y(n_5599)
);

INVx2_ASAP7_75t_L g5600 ( 
.A(n_5098),
.Y(n_5600)
);

INVx2_ASAP7_75t_SL g5601 ( 
.A(n_5281),
.Y(n_5601)
);

INVx1_ASAP7_75t_L g5602 ( 
.A(n_5441),
.Y(n_5602)
);

NAND3xp33_ASAP7_75t_L g5603 ( 
.A(n_5151),
.B(n_4982),
.C(n_4960),
.Y(n_5603)
);

AOI22xp5_ASAP7_75t_L g5604 ( 
.A1(n_5051),
.A2(n_4749),
.B1(n_4726),
.B2(n_4928),
.Y(n_5604)
);

OAI22xp5_ASAP7_75t_L g5605 ( 
.A1(n_5185),
.A2(n_4748),
.B1(n_4901),
.B2(n_4898),
.Y(n_5605)
);

BUFx4f_ASAP7_75t_SL g5606 ( 
.A(n_5157),
.Y(n_5606)
);

AOI22xp33_ASAP7_75t_L g5607 ( 
.A1(n_5438),
.A2(n_4677),
.B1(n_4621),
.B2(n_4568),
.Y(n_5607)
);

INVx1_ASAP7_75t_L g5608 ( 
.A(n_5494),
.Y(n_5608)
);

CKINVDCx8_ASAP7_75t_R g5609 ( 
.A(n_5054),
.Y(n_5609)
);

AOI22xp33_ASAP7_75t_L g5610 ( 
.A1(n_5183),
.A2(n_4677),
.B1(n_4621),
.B2(n_4568),
.Y(n_5610)
);

OAI21xp33_ASAP7_75t_L g5611 ( 
.A1(n_5025),
.A2(n_4969),
.B(n_4830),
.Y(n_5611)
);

AOI22xp33_ASAP7_75t_L g5612 ( 
.A1(n_5018),
.A2(n_4621),
.B1(n_4952),
.B2(n_4839),
.Y(n_5612)
);

OAI21xp33_ASAP7_75t_L g5613 ( 
.A1(n_5128),
.A2(n_4830),
.B(n_4900),
.Y(n_5613)
);

INVx4_ASAP7_75t_L g5614 ( 
.A(n_5054),
.Y(n_5614)
);

AOI22xp33_ASAP7_75t_L g5615 ( 
.A1(n_5144),
.A2(n_4621),
.B1(n_4839),
.B2(n_4868),
.Y(n_5615)
);

AOI22xp33_ASAP7_75t_L g5616 ( 
.A1(n_5026),
.A2(n_4868),
.B1(n_4672),
.B2(n_4921),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5510),
.Y(n_5617)
);

OAI22xp5_ASAP7_75t_L g5618 ( 
.A1(n_5203),
.A2(n_4866),
.B1(n_4975),
.B2(n_4780),
.Y(n_5618)
);

INVx1_ASAP7_75t_L g5619 ( 
.A(n_5029),
.Y(n_5619)
);

INVx2_ASAP7_75t_L g5620 ( 
.A(n_5098),
.Y(n_5620)
);

OR2x2_ASAP7_75t_SL g5621 ( 
.A(n_5366),
.B(n_4529),
.Y(n_5621)
);

AOI22xp33_ASAP7_75t_L g5622 ( 
.A1(n_5026),
.A2(n_4640),
.B1(n_4641),
.B2(n_4623),
.Y(n_5622)
);

AOI22xp33_ASAP7_75t_L g5623 ( 
.A1(n_5026),
.A2(n_4640),
.B1(n_4641),
.B2(n_4623),
.Y(n_5623)
);

AOI22xp33_ASAP7_75t_L g5624 ( 
.A1(n_5026),
.A2(n_4641),
.B1(n_4653),
.B2(n_4640),
.Y(n_5624)
);

AND2x4_ASAP7_75t_L g5625 ( 
.A(n_5368),
.B(n_4541),
.Y(n_5625)
);

INVx1_ASAP7_75t_L g5626 ( 
.A(n_5029),
.Y(n_5626)
);

INVx2_ASAP7_75t_L g5627 ( 
.A(n_5098),
.Y(n_5627)
);

AOI22xp33_ASAP7_75t_L g5628 ( 
.A1(n_5174),
.A2(n_4641),
.B1(n_4653),
.B2(n_4640),
.Y(n_5628)
);

INVx1_ASAP7_75t_L g5629 ( 
.A(n_5038),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_5038),
.Y(n_5630)
);

NAND2xp5_ASAP7_75t_L g5631 ( 
.A(n_5027),
.B(n_4840),
.Y(n_5631)
);

BUFx2_ASAP7_75t_L g5632 ( 
.A(n_5321),
.Y(n_5632)
);

BUFx6f_ASAP7_75t_L g5633 ( 
.A(n_5054),
.Y(n_5633)
);

INVx2_ASAP7_75t_L g5634 ( 
.A(n_5098),
.Y(n_5634)
);

NAND2xp5_ASAP7_75t_L g5635 ( 
.A(n_5088),
.B(n_4840),
.Y(n_5635)
);

INVx1_ASAP7_75t_L g5636 ( 
.A(n_5042),
.Y(n_5636)
);

INVx2_ASAP7_75t_L g5637 ( 
.A(n_5104),
.Y(n_5637)
);

OAI22xp5_ASAP7_75t_L g5638 ( 
.A1(n_5078),
.A2(n_5485),
.B1(n_5507),
.B2(n_5479),
.Y(n_5638)
);

INVx1_ASAP7_75t_L g5639 ( 
.A(n_5042),
.Y(n_5639)
);

AND2x2_ASAP7_75t_L g5640 ( 
.A(n_5016),
.B(n_4735),
.Y(n_5640)
);

CKINVDCx5p33_ASAP7_75t_R g5641 ( 
.A(n_5260),
.Y(n_5641)
);

OAI222xp33_ASAP7_75t_L g5642 ( 
.A1(n_5037),
.A2(n_4927),
.B1(n_4712),
.B2(n_5014),
.C1(n_4953),
.C2(n_4808),
.Y(n_5642)
);

AOI22xp5_ASAP7_75t_L g5643 ( 
.A1(n_5060),
.A2(n_4556),
.B1(n_4580),
.B2(n_4547),
.Y(n_5643)
);

AOI22xp5_ASAP7_75t_L g5644 ( 
.A1(n_5033),
.A2(n_4615),
.B1(n_4622),
.B2(n_4603),
.Y(n_5644)
);

INVx2_ASAP7_75t_L g5645 ( 
.A(n_5104),
.Y(n_5645)
);

OAI21xp33_ASAP7_75t_L g5646 ( 
.A1(n_5223),
.A2(n_5014),
.B(n_4784),
.Y(n_5646)
);

CKINVDCx14_ASAP7_75t_R g5647 ( 
.A(n_5024),
.Y(n_5647)
);

NAND2xp5_ASAP7_75t_L g5648 ( 
.A(n_5415),
.B(n_4855),
.Y(n_5648)
);

AOI22xp33_ASAP7_75t_L g5649 ( 
.A1(n_5170),
.A2(n_4653),
.B1(n_4716),
.B2(n_4729),
.Y(n_5649)
);

INVx2_ASAP7_75t_L g5650 ( 
.A(n_5104),
.Y(n_5650)
);

CKINVDCx5p33_ASAP7_75t_R g5651 ( 
.A(n_5157),
.Y(n_5651)
);

AOI22xp33_ASAP7_75t_L g5652 ( 
.A1(n_5034),
.A2(n_5439),
.B1(n_5452),
.B2(n_5230),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_5045),
.Y(n_5653)
);

CKINVDCx20_ASAP7_75t_R g5654 ( 
.A(n_5319),
.Y(n_5654)
);

CKINVDCx20_ASAP7_75t_R g5655 ( 
.A(n_5426),
.Y(n_5655)
);

AOI22xp33_ASAP7_75t_L g5656 ( 
.A1(n_5034),
.A2(n_4653),
.B1(n_4723),
.B2(n_4722),
.Y(n_5656)
);

AOI22xp33_ASAP7_75t_L g5657 ( 
.A1(n_5034),
.A2(n_4722),
.B1(n_4723),
.B2(n_4880),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5039),
.B(n_4735),
.Y(n_5658)
);

OAI222xp33_ASAP7_75t_L g5659 ( 
.A1(n_5017),
.A2(n_4712),
.B1(n_4953),
.B2(n_4808),
.C1(n_4880),
.C2(n_4908),
.Y(n_5659)
);

BUFx2_ASAP7_75t_L g5660 ( 
.A(n_5321),
.Y(n_5660)
);

AOI22xp33_ASAP7_75t_L g5661 ( 
.A1(n_5034),
.A2(n_4722),
.B1(n_4723),
.B2(n_4880),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5045),
.Y(n_5662)
);

BUFx12f_ASAP7_75t_L g5663 ( 
.A(n_5243),
.Y(n_5663)
);

OAI22xp5_ASAP7_75t_L g5664 ( 
.A1(n_5259),
.A2(n_4975),
.B1(n_4522),
.B2(n_4712),
.Y(n_5664)
);

INVx4_ASAP7_75t_L g5665 ( 
.A(n_5054),
.Y(n_5665)
);

BUFx6f_ASAP7_75t_L g5666 ( 
.A(n_5054),
.Y(n_5666)
);

OAI22xp5_ASAP7_75t_L g5667 ( 
.A1(n_5252),
.A2(n_4522),
.B1(n_4541),
.B2(n_4532),
.Y(n_5667)
);

AOI22xp33_ASAP7_75t_SL g5668 ( 
.A1(n_5057),
.A2(n_4683),
.B1(n_4704),
.B2(n_4671),
.Y(n_5668)
);

BUFx6f_ASAP7_75t_L g5669 ( 
.A(n_5020),
.Y(n_5669)
);

INVx1_ASAP7_75t_L g5670 ( 
.A(n_5050),
.Y(n_5670)
);

INVx2_ASAP7_75t_L g5671 ( 
.A(n_5104),
.Y(n_5671)
);

AOI22xp33_ASAP7_75t_L g5672 ( 
.A1(n_5439),
.A2(n_4723),
.B1(n_4722),
.B2(n_4880),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_5125),
.Y(n_5673)
);

NAND2xp5_ASAP7_75t_L g5674 ( 
.A(n_5056),
.B(n_4855),
.Y(n_5674)
);

INVx1_ASAP7_75t_L g5675 ( 
.A(n_5050),
.Y(n_5675)
);

OAI22xp5_ASAP7_75t_L g5676 ( 
.A1(n_5258),
.A2(n_4541),
.B1(n_4618),
.B2(n_4532),
.Y(n_5676)
);

INVx1_ASAP7_75t_L g5677 ( 
.A(n_5061),
.Y(n_5677)
);

AOI22xp33_ASAP7_75t_L g5678 ( 
.A1(n_5439),
.A2(n_4880),
.B1(n_5002),
.B2(n_4896),
.Y(n_5678)
);

INVx1_ASAP7_75t_L g5679 ( 
.A(n_5061),
.Y(n_5679)
);

AOI22xp33_ASAP7_75t_L g5680 ( 
.A1(n_5439),
.A2(n_4880),
.B1(n_5002),
.B2(n_4896),
.Y(n_5680)
);

INVx3_ASAP7_75t_SL g5681 ( 
.A(n_5243),
.Y(n_5681)
);

AOI22xp33_ASAP7_75t_L g5682 ( 
.A1(n_5439),
.A2(n_4896),
.B1(n_5002),
.B2(n_4954),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_5073),
.Y(n_5683)
);

AOI22xp33_ASAP7_75t_L g5684 ( 
.A1(n_5452),
.A2(n_4896),
.B1(n_5002),
.B2(n_4954),
.Y(n_5684)
);

INVxp67_ASAP7_75t_L g5685 ( 
.A(n_5131),
.Y(n_5685)
);

OAI22xp5_ASAP7_75t_SL g5686 ( 
.A1(n_5230),
.A2(n_4848),
.B1(n_4954),
.B2(n_4855),
.Y(n_5686)
);

INVx2_ASAP7_75t_L g5687 ( 
.A(n_5125),
.Y(n_5687)
);

AOI22xp33_ASAP7_75t_L g5688 ( 
.A1(n_5452),
.A2(n_4991),
.B1(n_4534),
.B2(n_4841),
.Y(n_5688)
);

AOI22xp33_ASAP7_75t_L g5689 ( 
.A1(n_5452),
.A2(n_4991),
.B1(n_4534),
.B2(n_4841),
.Y(n_5689)
);

AOI22xp33_ASAP7_75t_L g5690 ( 
.A1(n_5452),
.A2(n_4991),
.B1(n_4534),
.B2(n_4841),
.Y(n_5690)
);

OAI22xp5_ASAP7_75t_L g5691 ( 
.A1(n_5039),
.A2(n_4541),
.B1(n_4618),
.B2(n_4532),
.Y(n_5691)
);

NAND2xp5_ASAP7_75t_L g5692 ( 
.A(n_5080),
.B(n_4864),
.Y(n_5692)
);

OAI22x1_ASAP7_75t_L g5693 ( 
.A1(n_5540),
.A2(n_4531),
.B1(n_4637),
.B2(n_4881),
.Y(n_5693)
);

AOI211xp5_ASAP7_75t_L g5694 ( 
.A1(n_5188),
.A2(n_4982),
.B(n_4590),
.C(n_4762),
.Y(n_5694)
);

BUFx8_ASAP7_75t_L g5695 ( 
.A(n_5020),
.Y(n_5695)
);

AOI22xp33_ASAP7_75t_L g5696 ( 
.A1(n_5230),
.A2(n_4841),
.B1(n_4856),
.B2(n_4835),
.Y(n_5696)
);

BUFx12f_ASAP7_75t_L g5697 ( 
.A(n_5024),
.Y(n_5697)
);

BUFx6f_ASAP7_75t_L g5698 ( 
.A(n_5108),
.Y(n_5698)
);

HB1xp67_ASAP7_75t_L g5699 ( 
.A(n_5175),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5073),
.Y(n_5700)
);

INVx4_ASAP7_75t_L g5701 ( 
.A(n_5108),
.Y(n_5701)
);

OAI22xp5_ASAP7_75t_L g5702 ( 
.A1(n_5083),
.A2(n_4541),
.B1(n_4618),
.B2(n_4532),
.Y(n_5702)
);

AOI22xp33_ASAP7_75t_L g5703 ( 
.A1(n_5458),
.A2(n_4856),
.B1(n_4835),
.B2(n_4541),
.Y(n_5703)
);

OAI22xp5_ASAP7_75t_L g5704 ( 
.A1(n_5083),
.A2(n_4629),
.B1(n_4618),
.B2(n_4885),
.Y(n_5704)
);

CKINVDCx5p33_ASAP7_75t_R g5705 ( 
.A(n_5437),
.Y(n_5705)
);

BUFx4f_ASAP7_75t_SL g5706 ( 
.A(n_5311),
.Y(n_5706)
);

AND2x2_ASAP7_75t_L g5707 ( 
.A(n_5086),
.B(n_4881),
.Y(n_5707)
);

AND2x2_ASAP7_75t_L g5708 ( 
.A(n_5086),
.B(n_4923),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_5074),
.Y(n_5709)
);

AOI22xp33_ASAP7_75t_L g5710 ( 
.A1(n_5458),
.A2(n_4856),
.B1(n_4835),
.B2(n_4965),
.Y(n_5710)
);

OAI22xp5_ASAP7_75t_SL g5711 ( 
.A1(n_5138),
.A2(n_4531),
.B1(n_4637),
.B2(n_5009),
.Y(n_5711)
);

INVx1_ASAP7_75t_L g5712 ( 
.A(n_5074),
.Y(n_5712)
);

AOI22xp33_ASAP7_75t_SL g5713 ( 
.A1(n_5365),
.A2(n_4671),
.B1(n_4704),
.B2(n_4683),
.Y(n_5713)
);

INVx1_ASAP7_75t_L g5714 ( 
.A(n_5082),
.Y(n_5714)
);

BUFx8_ASAP7_75t_SL g5715 ( 
.A(n_5311),
.Y(n_5715)
);

BUFx3_ASAP7_75t_L g5716 ( 
.A(n_5304),
.Y(n_5716)
);

OAI21xp5_ASAP7_75t_L g5717 ( 
.A1(n_5022),
.A2(n_4753),
.B(n_4746),
.Y(n_5717)
);

CKINVDCx5p33_ASAP7_75t_R g5718 ( 
.A(n_5426),
.Y(n_5718)
);

HB1xp67_ASAP7_75t_L g5719 ( 
.A(n_5191),
.Y(n_5719)
);

OAI21xp5_ASAP7_75t_SL g5720 ( 
.A1(n_5237),
.A2(n_5004),
.B(n_4885),
.Y(n_5720)
);

OAI222xp33_ASAP7_75t_L g5721 ( 
.A1(n_5531),
.A2(n_4908),
.B1(n_4923),
.B2(n_4815),
.C1(n_4683),
.C2(n_4704),
.Y(n_5721)
);

AOI22xp33_ASAP7_75t_L g5722 ( 
.A1(n_5281),
.A2(n_4856),
.B1(n_4835),
.B2(n_4965),
.Y(n_5722)
);

AOI22xp33_ASAP7_75t_SL g5723 ( 
.A1(n_5365),
.A2(n_4671),
.B1(n_4815),
.B2(n_4977),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5082),
.Y(n_5724)
);

OAI21xp5_ASAP7_75t_SL g5725 ( 
.A1(n_5337),
.A2(n_5004),
.B(n_4885),
.Y(n_5725)
);

AOI22xp33_ASAP7_75t_L g5726 ( 
.A1(n_5281),
.A2(n_4965),
.B1(n_4924),
.B2(n_4663),
.Y(n_5726)
);

AOI22xp33_ASAP7_75t_L g5727 ( 
.A1(n_5281),
.A2(n_5298),
.B1(n_5368),
.B2(n_5052),
.Y(n_5727)
);

AOI22xp33_ASAP7_75t_L g5728 ( 
.A1(n_5368),
.A2(n_4965),
.B1(n_4924),
.B2(n_4663),
.Y(n_5728)
);

INVx2_ASAP7_75t_L g5729 ( 
.A(n_5125),
.Y(n_5729)
);

AND2x4_ASAP7_75t_L g5730 ( 
.A(n_5211),
.B(n_5213),
.Y(n_5730)
);

INVx4_ASAP7_75t_L g5731 ( 
.A(n_5449),
.Y(n_5731)
);

AND2x2_ASAP7_75t_L g5732 ( 
.A(n_5091),
.B(n_4929),
.Y(n_5732)
);

OAI21xp5_ASAP7_75t_SL g5733 ( 
.A1(n_5031),
.A2(n_5004),
.B(n_4799),
.Y(n_5733)
);

AOI22xp33_ASAP7_75t_SL g5734 ( 
.A1(n_5091),
.A2(n_4815),
.B1(n_4977),
.B2(n_4965),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5090),
.Y(n_5735)
);

OAI22xp5_ASAP7_75t_L g5736 ( 
.A1(n_5167),
.A2(n_4629),
.B1(n_5009),
.B2(n_4924),
.Y(n_5736)
);

AOI22xp33_ASAP7_75t_SL g5737 ( 
.A1(n_5167),
.A2(n_4977),
.B1(n_5005),
.B2(n_4996),
.Y(n_5737)
);

AND2x2_ASAP7_75t_L g5738 ( 
.A(n_5267),
.B(n_4929),
.Y(n_5738)
);

BUFx6f_ASAP7_75t_L g5739 ( 
.A(n_5340),
.Y(n_5739)
);

BUFx6f_ASAP7_75t_L g5740 ( 
.A(n_5340),
.Y(n_5740)
);

INVx1_ASAP7_75t_L g5741 ( 
.A(n_5090),
.Y(n_5741)
);

OAI222xp33_ASAP7_75t_L g5742 ( 
.A1(n_5040),
.A2(n_4908),
.B1(n_4929),
.B2(n_4937),
.C1(n_4941),
.C2(n_4924),
.Y(n_5742)
);

AOI22xp33_ASAP7_75t_SL g5743 ( 
.A1(n_5267),
.A2(n_4977),
.B1(n_5005),
.B2(n_4996),
.Y(n_5743)
);

INVx1_ASAP7_75t_L g5744 ( 
.A(n_5094),
.Y(n_5744)
);

AOI22xp33_ASAP7_75t_L g5745 ( 
.A1(n_5318),
.A2(n_4924),
.B1(n_4629),
.B2(n_4612),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_5094),
.Y(n_5746)
);

BUFx12f_ASAP7_75t_L g5747 ( 
.A(n_5304),
.Y(n_5747)
);

HB1xp67_ASAP7_75t_L g5748 ( 
.A(n_5209),
.Y(n_5748)
);

INVx2_ASAP7_75t_L g5749 ( 
.A(n_5125),
.Y(n_5749)
);

AOI22xp33_ASAP7_75t_L g5750 ( 
.A1(n_5481),
.A2(n_4924),
.B1(n_4629),
.B2(n_4612),
.Y(n_5750)
);

AOI22xp33_ASAP7_75t_L g5751 ( 
.A1(n_5481),
.A2(n_4612),
.B1(n_4908),
.B2(n_4852),
.Y(n_5751)
);

NAND2xp5_ASAP7_75t_L g5752 ( 
.A(n_5019),
.B(n_4553),
.Y(n_5752)
);

INVx4_ASAP7_75t_L g5753 ( 
.A(n_5291),
.Y(n_5753)
);

BUFx12f_ASAP7_75t_L g5754 ( 
.A(n_5304),
.Y(n_5754)
);

OAI22xp33_ASAP7_75t_L g5755 ( 
.A1(n_5093),
.A2(n_4908),
.B1(n_5009),
.B2(n_4531),
.Y(n_5755)
);

NAND3xp33_ASAP7_75t_L g5756 ( 
.A(n_5265),
.B(n_4548),
.C(n_4918),
.Y(n_5756)
);

AND2x2_ASAP7_75t_L g5757 ( 
.A(n_5402),
.B(n_4877),
.Y(n_5757)
);

BUFx6f_ASAP7_75t_L g5758 ( 
.A(n_5291),
.Y(n_5758)
);

AND2x2_ASAP7_75t_L g5759 ( 
.A(n_5402),
.B(n_4877),
.Y(n_5759)
);

OAI222xp33_ASAP7_75t_L g5760 ( 
.A1(n_5289),
.A2(n_5387),
.B1(n_5303),
.B2(n_5300),
.C1(n_5398),
.C2(n_5263),
.Y(n_5760)
);

CKINVDCx14_ASAP7_75t_R g5761 ( 
.A(n_5288),
.Y(n_5761)
);

OR2x2_ASAP7_75t_L g5762 ( 
.A(n_5116),
.B(n_4983),
.Y(n_5762)
);

INVx1_ASAP7_75t_L g5763 ( 
.A(n_5105),
.Y(n_5763)
);

OAI22xp5_ASAP7_75t_L g5764 ( 
.A1(n_5461),
.A2(n_4967),
.B1(n_4773),
.B2(n_4828),
.Y(n_5764)
);

OAI222xp33_ASAP7_75t_L g5765 ( 
.A1(n_5513),
.A2(n_4908),
.B1(n_4937),
.B2(n_4941),
.C1(n_4773),
.C2(n_4828),
.Y(n_5765)
);

AOI22xp33_ASAP7_75t_L g5766 ( 
.A1(n_5048),
.A2(n_4612),
.B1(n_4852),
.B2(n_4769),
.Y(n_5766)
);

AOI22xp33_ASAP7_75t_L g5767 ( 
.A1(n_5048),
.A2(n_4612),
.B1(n_4852),
.B2(n_4769),
.Y(n_5767)
);

AOI22xp33_ASAP7_75t_L g5768 ( 
.A1(n_5048),
.A2(n_4612),
.B1(n_4852),
.B2(n_4769),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_5105),
.Y(n_5769)
);

INVx2_ASAP7_75t_L g5770 ( 
.A(n_5133),
.Y(n_5770)
);

AOI22xp33_ASAP7_75t_L g5771 ( 
.A1(n_5048),
.A2(n_4612),
.B1(n_4769),
.B2(n_4987),
.Y(n_5771)
);

INVx2_ASAP7_75t_L g5772 ( 
.A(n_5133),
.Y(n_5772)
);

NAND2xp5_ASAP7_75t_L g5773 ( 
.A(n_5233),
.B(n_4553),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5109),
.Y(n_5774)
);

CKINVDCx14_ASAP7_75t_R g5775 ( 
.A(n_5378),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5109),
.Y(n_5776)
);

OAI22xp5_ASAP7_75t_L g5777 ( 
.A1(n_5554),
.A2(n_4967),
.B1(n_4773),
.B2(n_4828),
.Y(n_5777)
);

OR2x2_ASAP7_75t_L g5778 ( 
.A(n_5116),
.B(n_4983),
.Y(n_5778)
);

INVx5_ASAP7_75t_SL g5779 ( 
.A(n_5269),
.Y(n_5779)
);

INVx2_ASAP7_75t_SL g5780 ( 
.A(n_5269),
.Y(n_5780)
);

HB1xp67_ASAP7_75t_L g5781 ( 
.A(n_5064),
.Y(n_5781)
);

AOI222xp33_ASAP7_75t_L g5782 ( 
.A1(n_5470),
.A2(n_4890),
.B1(n_4774),
.B2(n_4656),
.C1(n_4922),
.C2(n_4941),
.Y(n_5782)
);

AOI22xp33_ASAP7_75t_SL g5783 ( 
.A1(n_5242),
.A2(n_4977),
.B1(n_5005),
.B2(n_4996),
.Y(n_5783)
);

INVx1_ASAP7_75t_L g5784 ( 
.A(n_5112),
.Y(n_5784)
);

INVx1_ASAP7_75t_L g5785 ( 
.A(n_5112),
.Y(n_5785)
);

AOI22xp33_ASAP7_75t_L g5786 ( 
.A1(n_5279),
.A2(n_4612),
.B1(n_4769),
.B2(n_4987),
.Y(n_5786)
);

AOI22xp33_ASAP7_75t_L g5787 ( 
.A1(n_5279),
.A2(n_4612),
.B1(n_4769),
.B2(n_4987),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5193),
.B(n_5367),
.Y(n_5788)
);

AOI22xp33_ASAP7_75t_SL g5789 ( 
.A1(n_5242),
.A2(n_4996),
.B1(n_5005),
.B2(n_4922),
.Y(n_5789)
);

AND2x2_ASAP7_75t_L g5790 ( 
.A(n_5193),
.B(n_4877),
.Y(n_5790)
);

NAND2xp5_ASAP7_75t_L g5791 ( 
.A(n_5277),
.B(n_4670),
.Y(n_5791)
);

INVxp67_ASAP7_75t_SL g5792 ( 
.A(n_5312),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_5134),
.Y(n_5793)
);

BUFx12f_ASAP7_75t_L g5794 ( 
.A(n_5036),
.Y(n_5794)
);

AOI22xp33_ASAP7_75t_L g5795 ( 
.A1(n_5279),
.A2(n_4612),
.B1(n_4769),
.B2(n_4987),
.Y(n_5795)
);

OAI222xp33_ASAP7_75t_L g5796 ( 
.A1(n_5246),
.A2(n_4773),
.B1(n_4813),
.B2(n_4828),
.C1(n_4912),
.C2(n_4877),
.Y(n_5796)
);

INVx2_ASAP7_75t_L g5797 ( 
.A(n_5133),
.Y(n_5797)
);

INVxp67_ASAP7_75t_L g5798 ( 
.A(n_5087),
.Y(n_5798)
);

AOI22xp33_ASAP7_75t_L g5799 ( 
.A1(n_5297),
.A2(n_4612),
.B1(n_4769),
.B2(n_4992),
.Y(n_5799)
);

OAI22xp5_ASAP7_75t_L g5800 ( 
.A1(n_5058),
.A2(n_4967),
.B1(n_4813),
.B2(n_4637),
.Y(n_5800)
);

INVx1_ASAP7_75t_SL g5801 ( 
.A(n_5360),
.Y(n_5801)
);

AOI22xp33_ASAP7_75t_L g5802 ( 
.A1(n_5297),
.A2(n_4769),
.B1(n_4992),
.B2(n_4775),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5134),
.Y(n_5803)
);

AND2x2_ASAP7_75t_L g5804 ( 
.A(n_5367),
.B(n_4955),
.Y(n_5804)
);

AOI22xp33_ASAP7_75t_L g5805 ( 
.A1(n_5297),
.A2(n_4769),
.B1(n_4992),
.B2(n_4775),
.Y(n_5805)
);

NOR2x1p5_ASAP7_75t_L g5806 ( 
.A(n_5305),
.B(n_4656),
.Y(n_5806)
);

INVx1_ASAP7_75t_L g5807 ( 
.A(n_5135),
.Y(n_5807)
);

AOI22xp33_ASAP7_75t_SL g5808 ( 
.A1(n_5354),
.A2(n_4996),
.B1(n_5005),
.B2(n_4922),
.Y(n_5808)
);

INVx2_ASAP7_75t_L g5809 ( 
.A(n_5133),
.Y(n_5809)
);

NAND3xp33_ASAP7_75t_L g5810 ( 
.A(n_5455),
.B(n_4548),
.C(n_4762),
.Y(n_5810)
);

AOI222xp33_ASAP7_75t_L g5811 ( 
.A1(n_5399),
.A2(n_4774),
.B1(n_4922),
.B2(n_4799),
.C1(n_4913),
.C2(n_4709),
.Y(n_5811)
);

INVx1_ASAP7_75t_L g5812 ( 
.A(n_5135),
.Y(n_5812)
);

INVx2_ASAP7_75t_L g5813 ( 
.A(n_5143),
.Y(n_5813)
);

BUFx2_ASAP7_75t_L g5814 ( 
.A(n_5305),
.Y(n_5814)
);

OAI22xp33_ASAP7_75t_L g5815 ( 
.A1(n_5305),
.A2(n_4993),
.B1(n_4813),
.B2(n_4824),
.Y(n_5815)
);

AOI22xp33_ASAP7_75t_L g5816 ( 
.A1(n_5392),
.A2(n_4769),
.B1(n_4992),
.B2(n_4814),
.Y(n_5816)
);

AOI22xp33_ASAP7_75t_L g5817 ( 
.A1(n_5392),
.A2(n_4755),
.B1(n_4814),
.B2(n_4699),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5148),
.Y(n_5818)
);

OAI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_5058),
.A2(n_4967),
.B1(n_4813),
.B2(n_4993),
.Y(n_5819)
);

OAI22xp5_ASAP7_75t_L g5820 ( 
.A1(n_5072),
.A2(n_4993),
.B1(n_4814),
.B2(n_4755),
.Y(n_5820)
);

AND2x2_ASAP7_75t_L g5821 ( 
.A(n_5211),
.B(n_5213),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5148),
.Y(n_5822)
);

INVx3_ASAP7_75t_L g5823 ( 
.A(n_5164),
.Y(n_5823)
);

AOI22xp33_ASAP7_75t_L g5824 ( 
.A1(n_5211),
.A2(n_4755),
.B1(n_4814),
.B2(n_4699),
.Y(n_5824)
);

OAI22xp5_ASAP7_75t_L g5825 ( 
.A1(n_5072),
.A2(n_4993),
.B1(n_4755),
.B2(n_4824),
.Y(n_5825)
);

BUFx8_ASAP7_75t_SL g5826 ( 
.A(n_5310),
.Y(n_5826)
);

CKINVDCx11_ASAP7_75t_R g5827 ( 
.A(n_5036),
.Y(n_5827)
);

INVx1_ASAP7_75t_L g5828 ( 
.A(n_5154),
.Y(n_5828)
);

INVx2_ASAP7_75t_L g5829 ( 
.A(n_5143),
.Y(n_5829)
);

INVx3_ASAP7_75t_L g5830 ( 
.A(n_5164),
.Y(n_5830)
);

INVx4_ASAP7_75t_L g5831 ( 
.A(n_5114),
.Y(n_5831)
);

OAI22xp5_ASAP7_75t_L g5832 ( 
.A1(n_5195),
.A2(n_4993),
.B1(n_4824),
.B2(n_4946),
.Y(n_5832)
);

AND2x2_ASAP7_75t_L g5833 ( 
.A(n_5213),
.B(n_5351),
.Y(n_5833)
);

AOI22xp33_ASAP7_75t_L g5834 ( 
.A1(n_5351),
.A2(n_4980),
.B1(n_4955),
.B2(n_4535),
.Y(n_5834)
);

OR2x2_ASAP7_75t_L g5835 ( 
.A(n_5210),
.B(n_4670),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_5154),
.Y(n_5836)
);

HB1xp67_ASAP7_75t_L g5837 ( 
.A(n_5107),
.Y(n_5837)
);

INVx1_ASAP7_75t_L g5838 ( 
.A(n_5161),
.Y(n_5838)
);

AOI22xp33_ASAP7_75t_L g5839 ( 
.A1(n_5351),
.A2(n_4980),
.B1(n_4955),
.B2(n_4535),
.Y(n_5839)
);

AOI22xp33_ASAP7_75t_SL g5840 ( 
.A1(n_5354),
.A2(n_4922),
.B1(n_4548),
.B2(n_4873),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5161),
.Y(n_5841)
);

AOI22xp33_ASAP7_75t_L g5842 ( 
.A1(n_5379),
.A2(n_4980),
.B1(n_4955),
.B2(n_4535),
.Y(n_5842)
);

OAI21xp5_ASAP7_75t_SL g5843 ( 
.A1(n_5031),
.A2(n_4913),
.B(n_4970),
.Y(n_5843)
);

OAI21xp5_ASAP7_75t_SL g5844 ( 
.A1(n_5067),
.A2(n_4970),
.B(n_5013),
.Y(n_5844)
);

AOI21xp33_ASAP7_75t_L g5845 ( 
.A1(n_5240),
.A2(n_4980),
.B(n_4914),
.Y(n_5845)
);

AOI22xp33_ASAP7_75t_L g5846 ( 
.A1(n_5379),
.A2(n_4548),
.B1(n_4909),
.B2(n_4740),
.Y(n_5846)
);

AND2x2_ASAP7_75t_L g5847 ( 
.A(n_5379),
.B(n_5013),
.Y(n_5847)
);

NOR2x1_ASAP7_75t_L g5848 ( 
.A(n_5499),
.B(n_4676),
.Y(n_5848)
);

OAI21xp5_ASAP7_75t_SL g5849 ( 
.A1(n_5067),
.A2(n_4959),
.B(n_4995),
.Y(n_5849)
);

INVx2_ASAP7_75t_L g5850 ( 
.A(n_5143),
.Y(n_5850)
);

AND2x2_ASAP7_75t_L g5851 ( 
.A(n_5180),
.B(n_4627),
.Y(n_5851)
);

AND2x2_ASAP7_75t_L g5852 ( 
.A(n_5180),
.B(n_4627),
.Y(n_5852)
);

NOR2xp33_ASAP7_75t_L g5853 ( 
.A(n_5099),
.B(n_4676),
.Y(n_5853)
);

HB1xp67_ASAP7_75t_L g5854 ( 
.A(n_5113),
.Y(n_5854)
);

AND2x2_ASAP7_75t_L g5855 ( 
.A(n_5180),
.B(n_4657),
.Y(n_5855)
);

AOI222xp33_ASAP7_75t_L g5856 ( 
.A1(n_5370),
.A2(n_4709),
.B1(n_4646),
.B2(n_4611),
.C1(n_4938),
.C2(n_4916),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5163),
.Y(n_5857)
);

CKINVDCx8_ASAP7_75t_R g5858 ( 
.A(n_5414),
.Y(n_5858)
);

AOI22xp33_ASAP7_75t_SL g5859 ( 
.A1(n_5310),
.A2(n_4548),
.B1(n_4873),
.B2(n_5006),
.Y(n_5859)
);

AOI22xp33_ASAP7_75t_L g5860 ( 
.A1(n_5015),
.A2(n_4909),
.B1(n_4740),
.B2(n_4873),
.Y(n_5860)
);

AOI22xp33_ASAP7_75t_L g5861 ( 
.A1(n_5414),
.A2(n_4909),
.B1(n_4740),
.B2(n_4873),
.Y(n_5861)
);

AOI22xp33_ASAP7_75t_L g5862 ( 
.A1(n_5414),
.A2(n_4909),
.B1(n_4740),
.B2(n_4601),
.Y(n_5862)
);

INVx2_ASAP7_75t_L g5863 ( 
.A(n_5143),
.Y(n_5863)
);

AOI22xp33_ASAP7_75t_L g5864 ( 
.A1(n_5414),
.A2(n_5181),
.B1(n_5350),
.B2(n_5327),
.Y(n_5864)
);

BUFx3_ASAP7_75t_L g5865 ( 
.A(n_5195),
.Y(n_5865)
);

BUFx4f_ASAP7_75t_SL g5866 ( 
.A(n_5036),
.Y(n_5866)
);

AOI22xp33_ASAP7_75t_L g5867 ( 
.A1(n_5181),
.A2(n_4601),
.B1(n_4914),
.B2(n_4804),
.Y(n_5867)
);

AOI22xp33_ASAP7_75t_L g5868 ( 
.A1(n_5181),
.A2(n_4601),
.B1(n_4914),
.B2(n_4804),
.Y(n_5868)
);

OR2x2_ASAP7_75t_L g5869 ( 
.A(n_5210),
.B(n_4611),
.Y(n_5869)
);

BUFx2_ASAP7_75t_L g5870 ( 
.A(n_5310),
.Y(n_5870)
);

AOI222xp33_ASAP7_75t_L g5871 ( 
.A1(n_5489),
.A2(n_4646),
.B1(n_4938),
.B2(n_4916),
.C1(n_4865),
.C2(n_4675),
.Y(n_5871)
);

NAND2xp5_ASAP7_75t_L g5872 ( 
.A(n_5306),
.B(n_4884),
.Y(n_5872)
);

INVx2_ASAP7_75t_SL g5873 ( 
.A(n_5269),
.Y(n_5873)
);

AOI22xp33_ASAP7_75t_L g5874 ( 
.A1(n_5273),
.A2(n_4601),
.B1(n_4914),
.B2(n_4804),
.Y(n_5874)
);

AOI22xp33_ASAP7_75t_L g5875 ( 
.A1(n_5273),
.A2(n_4804),
.B1(n_4647),
.B2(n_4831),
.Y(n_5875)
);

NAND2xp5_ASAP7_75t_L g5876 ( 
.A(n_5286),
.B(n_4887),
.Y(n_5876)
);

CKINVDCx5p33_ASAP7_75t_R g5877 ( 
.A(n_5089),
.Y(n_5877)
);

AOI22xp33_ASAP7_75t_L g5878 ( 
.A1(n_5327),
.A2(n_4647),
.B1(n_4831),
.B2(n_4824),
.Y(n_5878)
);

INVx2_ASAP7_75t_L g5879 ( 
.A(n_5401),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5163),
.Y(n_5880)
);

AOI22xp33_ASAP7_75t_L g5881 ( 
.A1(n_5349),
.A2(n_4647),
.B1(n_4831),
.B2(n_4824),
.Y(n_5881)
);

AOI22xp33_ASAP7_75t_L g5882 ( 
.A1(n_5349),
.A2(n_4647),
.B1(n_4831),
.B2(n_4824),
.Y(n_5882)
);

NAND2xp5_ASAP7_75t_L g5883 ( 
.A(n_5290),
.B(n_4887),
.Y(n_5883)
);

INVx2_ASAP7_75t_SL g5884 ( 
.A(n_5269),
.Y(n_5884)
);

AOI22xp33_ASAP7_75t_L g5885 ( 
.A1(n_5440),
.A2(n_4824),
.B1(n_4946),
.B2(n_4759),
.Y(n_5885)
);

AOI22xp33_ASAP7_75t_SL g5886 ( 
.A1(n_5359),
.A2(n_5006),
.B1(n_4925),
.B2(n_4938),
.Y(n_5886)
);

BUFx4f_ASAP7_75t_SL g5887 ( 
.A(n_5440),
.Y(n_5887)
);

BUFx3_ASAP7_75t_L g5888 ( 
.A(n_5451),
.Y(n_5888)
);

OAI21xp5_ASAP7_75t_SL g5889 ( 
.A1(n_5488),
.A2(n_4959),
.B(n_4995),
.Y(n_5889)
);

OAI21xp33_ASAP7_75t_L g5890 ( 
.A1(n_5421),
.A2(n_5491),
.B(n_5156),
.Y(n_5890)
);

INVx1_ASAP7_75t_L g5891 ( 
.A(n_5169),
.Y(n_5891)
);

INVx4_ASAP7_75t_L g5892 ( 
.A(n_5269),
.Y(n_5892)
);

OAI22xp5_ASAP7_75t_L g5893 ( 
.A1(n_5359),
.A2(n_4946),
.B1(n_4759),
.B2(n_4809),
.Y(n_5893)
);

INVx2_ASAP7_75t_SL g5894 ( 
.A(n_5301),
.Y(n_5894)
);

OR2x2_ASAP7_75t_L g5895 ( 
.A(n_5192),
.B(n_4536),
.Y(n_5895)
);

AOI22xp33_ASAP7_75t_L g5896 ( 
.A1(n_5451),
.A2(n_5359),
.B1(n_5152),
.B2(n_5124),
.Y(n_5896)
);

INVx3_ASAP7_75t_L g5897 ( 
.A(n_5164),
.Y(n_5897)
);

AOI22xp33_ASAP7_75t_SL g5898 ( 
.A1(n_5376),
.A2(n_5006),
.B1(n_4925),
.B2(n_4916),
.Y(n_5898)
);

AOI22xp5_ASAP7_75t_L g5899 ( 
.A1(n_5096),
.A2(n_4865),
.B1(n_4675),
.B2(n_4718),
.Y(n_5899)
);

AND2x2_ASAP7_75t_L g5900 ( 
.A(n_5124),
.B(n_4657),
.Y(n_5900)
);

INVx1_ASAP7_75t_L g5901 ( 
.A(n_5169),
.Y(n_5901)
);

AND2x2_ASAP7_75t_L g5902 ( 
.A(n_5124),
.B(n_4718),
.Y(n_5902)
);

OAI21xp5_ASAP7_75t_SL g5903 ( 
.A1(n_5283),
.A2(n_5003),
.B(n_4995),
.Y(n_5903)
);

BUFx3_ASAP7_75t_L g5904 ( 
.A(n_5301),
.Y(n_5904)
);

BUFx12f_ASAP7_75t_L g5905 ( 
.A(n_5301),
.Y(n_5905)
);

INVx2_ASAP7_75t_L g5906 ( 
.A(n_5401),
.Y(n_5906)
);

INVx1_ASAP7_75t_L g5907 ( 
.A(n_5173),
.Y(n_5907)
);

AOI22xp33_ASAP7_75t_L g5908 ( 
.A1(n_5152),
.A2(n_4759),
.B1(n_4946),
.B2(n_4827),
.Y(n_5908)
);

NAND2xp5_ASAP7_75t_L g5909 ( 
.A(n_5156),
.B(n_4894),
.Y(n_5909)
);

INVx2_ASAP7_75t_L g5910 ( 
.A(n_5401),
.Y(n_5910)
);

AOI22xp33_ASAP7_75t_L g5911 ( 
.A1(n_5309),
.A2(n_4759),
.B1(n_4946),
.B2(n_4827),
.Y(n_5911)
);

CKINVDCx20_ASAP7_75t_R g5912 ( 
.A(n_5450),
.Y(n_5912)
);

AOI22xp33_ASAP7_75t_L g5913 ( 
.A1(n_5309),
.A2(n_4759),
.B1(n_4946),
.B2(n_4827),
.Y(n_5913)
);

AOI22xp33_ASAP7_75t_L g5914 ( 
.A1(n_5309),
.A2(n_4759),
.B1(n_4946),
.B2(n_4827),
.Y(n_5914)
);

OAI22xp5_ASAP7_75t_SL g5915 ( 
.A1(n_5312),
.A2(n_4759),
.B1(n_4809),
.B2(n_4764),
.Y(n_5915)
);

AOI22xp33_ASAP7_75t_L g5916 ( 
.A1(n_5422),
.A2(n_4962),
.B1(n_4865),
.B2(n_4675),
.Y(n_5916)
);

INVx1_ASAP7_75t_L g5917 ( 
.A(n_5173),
.Y(n_5917)
);

AOI22xp33_ASAP7_75t_L g5918 ( 
.A1(n_5422),
.A2(n_4962),
.B1(n_4865),
.B2(n_4675),
.Y(n_5918)
);

AOI22xp33_ASAP7_75t_L g5919 ( 
.A1(n_5443),
.A2(n_4962),
.B1(n_4865),
.B2(n_4675),
.Y(n_5919)
);

NOR2x1_ASAP7_75t_L g5920 ( 
.A(n_5095),
.B(n_4676),
.Y(n_5920)
);

OAI22xp33_ASAP7_75t_L g5921 ( 
.A1(n_5353),
.A2(n_4809),
.B1(n_4810),
.B2(n_4764),
.Y(n_5921)
);

AOI22xp33_ASAP7_75t_L g5922 ( 
.A1(n_5443),
.A2(n_4962),
.B1(n_4741),
.B2(n_4995),
.Y(n_5922)
);

INVx4_ASAP7_75t_L g5923 ( 
.A(n_5301),
.Y(n_5923)
);

INVx2_ASAP7_75t_L g5924 ( 
.A(n_5097),
.Y(n_5924)
);

INVx2_ASAP7_75t_SL g5925 ( 
.A(n_5301),
.Y(n_5925)
);

INVx1_ASAP7_75t_L g5926 ( 
.A(n_5182),
.Y(n_5926)
);

AOI22xp33_ASAP7_75t_SL g5927 ( 
.A1(n_5102),
.A2(n_5006),
.B1(n_4925),
.B2(n_4916),
.Y(n_5927)
);

INVx1_ASAP7_75t_L g5928 ( 
.A(n_5182),
.Y(n_5928)
);

HB1xp67_ASAP7_75t_L g5929 ( 
.A(n_5047),
.Y(n_5929)
);

AOI22xp33_ASAP7_75t_SL g5930 ( 
.A1(n_5102),
.A2(n_5006),
.B1(n_4925),
.B2(n_4916),
.Y(n_5930)
);

INVx1_ASAP7_75t_L g5931 ( 
.A(n_5196),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5196),
.Y(n_5932)
);

BUFx3_ASAP7_75t_L g5933 ( 
.A(n_5095),
.Y(n_5933)
);

HB1xp67_ASAP7_75t_L g5934 ( 
.A(n_5047),
.Y(n_5934)
);

AOI22xp33_ASAP7_75t_L g5935 ( 
.A1(n_5478),
.A2(n_5102),
.B1(n_5543),
.B2(n_5520),
.Y(n_5935)
);

INVx2_ASAP7_75t_L g5936 ( 
.A(n_5097),
.Y(n_5936)
);

NAND2xp5_ASAP7_75t_L g5937 ( 
.A(n_5244),
.B(n_4894),
.Y(n_5937)
);

OAI22xp5_ASAP7_75t_SL g5938 ( 
.A1(n_5312),
.A2(n_4764),
.B1(n_4810),
.B2(n_4529),
.Y(n_5938)
);

INVx2_ASAP7_75t_L g5939 ( 
.A(n_5100),
.Y(n_5939)
);

BUFx6f_ASAP7_75t_L g5940 ( 
.A(n_5220),
.Y(n_5940)
);

AOI22xp33_ASAP7_75t_L g5941 ( 
.A1(n_5478),
.A2(n_5543),
.B1(n_5520),
.B2(n_5332),
.Y(n_5941)
);

AOI22xp33_ASAP7_75t_L g5942 ( 
.A1(n_5520),
.A2(n_5332),
.B1(n_5372),
.B2(n_5371),
.Y(n_5942)
);

INVx1_ASAP7_75t_L g5943 ( 
.A(n_5197),
.Y(n_5943)
);

AOI22xp33_ASAP7_75t_L g5944 ( 
.A1(n_5520),
.A2(n_4741),
.B1(n_5003),
.B2(n_4823),
.Y(n_5944)
);

AOI22xp33_ASAP7_75t_L g5945 ( 
.A1(n_5520),
.A2(n_4741),
.B1(n_5003),
.B2(n_4823),
.Y(n_5945)
);

AND2x2_ASAP7_75t_L g5946 ( 
.A(n_5348),
.B(n_4728),
.Y(n_5946)
);

OAI21xp5_ASAP7_75t_SL g5947 ( 
.A1(n_5245),
.A2(n_5003),
.B(n_4728),
.Y(n_5947)
);

BUFx3_ASAP7_75t_L g5948 ( 
.A(n_5095),
.Y(n_5948)
);

OAI22xp5_ASAP7_75t_L g5949 ( 
.A1(n_5214),
.A2(n_4810),
.B1(n_4747),
.B2(n_4676),
.Y(n_5949)
);

AOI22xp33_ASAP7_75t_L g5950 ( 
.A1(n_5520),
.A2(n_4741),
.B1(n_4851),
.B2(n_4925),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5197),
.Y(n_5951)
);

BUFx6f_ASAP7_75t_L g5952 ( 
.A(n_5220),
.Y(n_5952)
);

CKINVDCx11_ASAP7_75t_R g5953 ( 
.A(n_5220),
.Y(n_5953)
);

INVx1_ASAP7_75t_L g5954 ( 
.A(n_5202),
.Y(n_5954)
);

BUFx4f_ASAP7_75t_SL g5955 ( 
.A(n_5530),
.Y(n_5955)
);

AOI222xp33_ASAP7_75t_L g5956 ( 
.A1(n_5501),
.A2(n_4944),
.B1(n_4939),
.B2(n_4974),
.C1(n_5000),
.C2(n_4931),
.Y(n_5956)
);

AOI22xp33_ASAP7_75t_L g5957 ( 
.A1(n_5520),
.A2(n_5332),
.B1(n_5063),
.B2(n_5160),
.Y(n_5957)
);

AOI22xp33_ASAP7_75t_L g5958 ( 
.A1(n_5063),
.A2(n_4851),
.B1(n_4944),
.B2(n_4963),
.Y(n_5958)
);

AOI22xp33_ASAP7_75t_L g5959 ( 
.A1(n_5063),
.A2(n_4851),
.B1(n_4944),
.B2(n_4963),
.Y(n_5959)
);

BUFx5_ASAP7_75t_L g5960 ( 
.A(n_5544),
.Y(n_5960)
);

OAI22xp5_ASAP7_75t_L g5961 ( 
.A1(n_5530),
.A2(n_4821),
.B1(n_4932),
.B2(n_4747),
.Y(n_5961)
);

INVx2_ASAP7_75t_SL g5962 ( 
.A(n_5220),
.Y(n_5962)
);

INVx1_ASAP7_75t_L g5963 ( 
.A(n_5202),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5208),
.Y(n_5964)
);

AND2x2_ASAP7_75t_L g5965 ( 
.A(n_5348),
.B(n_4747),
.Y(n_5965)
);

OR2x2_ASAP7_75t_L g5966 ( 
.A(n_5192),
.B(n_4536),
.Y(n_5966)
);

OAI22xp5_ASAP7_75t_L g5967 ( 
.A1(n_5035),
.A2(n_4821),
.B1(n_4932),
.B2(n_4747),
.Y(n_5967)
);

INVx2_ASAP7_75t_L g5968 ( 
.A(n_5100),
.Y(n_5968)
);

OR2x2_ASAP7_75t_L g5969 ( 
.A(n_5207),
.B(n_4536),
.Y(n_5969)
);

AOI22xp33_ASAP7_75t_SL g5970 ( 
.A1(n_5172),
.A2(n_5538),
.B1(n_5547),
.B2(n_5446),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5208),
.Y(n_5971)
);

AOI22xp33_ASAP7_75t_L g5972 ( 
.A1(n_5063),
.A2(n_4851),
.B1(n_4963),
.B2(n_4893),
.Y(n_5972)
);

INVx3_ASAP7_75t_L g5973 ( 
.A(n_5164),
.Y(n_5973)
);

AOI22xp33_ASAP7_75t_L g5974 ( 
.A1(n_5224),
.A2(n_5547),
.B1(n_5446),
.B2(n_5512),
.Y(n_5974)
);

HB1xp67_ASAP7_75t_L g5975 ( 
.A(n_5047),
.Y(n_5975)
);

OAI22xp5_ASAP7_75t_L g5976 ( 
.A1(n_5383),
.A2(n_4932),
.B1(n_4935),
.B2(n_4821),
.Y(n_5976)
);

NAND2xp5_ASAP7_75t_L g5977 ( 
.A(n_5271),
.B(n_4904),
.Y(n_5977)
);

AOI22xp33_ASAP7_75t_L g5978 ( 
.A1(n_5446),
.A2(n_4851),
.B1(n_4963),
.B2(n_4893),
.Y(n_5978)
);

OAI22xp5_ASAP7_75t_L g5979 ( 
.A1(n_5383),
.A2(n_4932),
.B1(n_4935),
.B2(n_4821),
.Y(n_5979)
);

AOI22xp33_ASAP7_75t_SL g5980 ( 
.A1(n_5172),
.A2(n_4680),
.B1(n_4605),
.B2(n_4635),
.Y(n_5980)
);

BUFx4f_ASAP7_75t_SL g5981 ( 
.A(n_5547),
.Y(n_5981)
);

BUFx2_ASAP7_75t_L g5982 ( 
.A(n_5285),
.Y(n_5982)
);

NAND2xp5_ASAP7_75t_L g5983 ( 
.A(n_5121),
.B(n_4904),
.Y(n_5983)
);

INVx1_ASAP7_75t_L g5984 ( 
.A(n_5217),
.Y(n_5984)
);

OAI22xp5_ASAP7_75t_L g5985 ( 
.A1(n_5044),
.A2(n_5012),
.B1(n_4935),
.B2(n_4910),
.Y(n_5985)
);

AOI222xp33_ASAP7_75t_L g5986 ( 
.A1(n_5212),
.A2(n_4915),
.B1(n_4951),
.B2(n_4966),
.C1(n_4910),
.C2(n_5000),
.Y(n_5986)
);

INVx1_ASAP7_75t_L g5987 ( 
.A(n_5217),
.Y(n_5987)
);

AOI22xp33_ASAP7_75t_L g5988 ( 
.A1(n_5278),
.A2(n_4963),
.B1(n_4893),
.B2(n_4935),
.Y(n_5988)
);

CKINVDCx5p33_ASAP7_75t_R g5989 ( 
.A(n_5285),
.Y(n_5989)
);

AND2x4_ASAP7_75t_L g5990 ( 
.A(n_5200),
.B(n_4658),
.Y(n_5990)
);

BUFx6f_ASAP7_75t_SL g5991 ( 
.A(n_5285),
.Y(n_5991)
);

AOI22xp33_ASAP7_75t_SL g5992 ( 
.A1(n_5538),
.A2(n_4680),
.B1(n_4605),
.B2(n_4635),
.Y(n_5992)
);

INVx2_ASAP7_75t_L g5993 ( 
.A(n_5021),
.Y(n_5993)
);

BUFx2_ASAP7_75t_L g5994 ( 
.A(n_5285),
.Y(n_5994)
);

HB1xp67_ASAP7_75t_L g5995 ( 
.A(n_5153),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5222),
.Y(n_5996)
);

AOI22xp33_ASAP7_75t_L g5997 ( 
.A1(n_5110),
.A2(n_5386),
.B1(n_5526),
.B2(n_5423),
.Y(n_5997)
);

AOI22xp33_ASAP7_75t_L g5998 ( 
.A1(n_5110),
.A2(n_4893),
.B1(n_5012),
.B2(n_4605),
.Y(n_5998)
);

AOI22xp33_ASAP7_75t_SL g5999 ( 
.A1(n_5334),
.A2(n_4680),
.B1(n_4605),
.B2(n_4635),
.Y(n_5999)
);

NOR2xp33_ASAP7_75t_L g6000 ( 
.A(n_5231),
.B(n_5012),
.Y(n_6000)
);

INVx3_ASAP7_75t_L g6001 ( 
.A(n_5155),
.Y(n_6001)
);

OAI22xp33_ASAP7_75t_L g6002 ( 
.A1(n_5044),
.A2(n_5012),
.B1(n_4893),
.B2(n_4605),
.Y(n_6002)
);

INVx2_ASAP7_75t_L g6003 ( 
.A(n_5021),
.Y(n_6003)
);

INVx3_ASAP7_75t_L g6004 ( 
.A(n_5155),
.Y(n_6004)
);

AOI22xp33_ASAP7_75t_L g6005 ( 
.A1(n_5110),
.A2(n_4994),
.B1(n_4843),
.B2(n_4786),
.Y(n_6005)
);

INVx1_ASAP7_75t_L g6006 ( 
.A(n_5222),
.Y(n_6006)
);

AND2x2_ASAP7_75t_L g6007 ( 
.A(n_5384),
.B(n_4536),
.Y(n_6007)
);

OAI21xp33_ASAP7_75t_L g6008 ( 
.A1(n_5328),
.A2(n_5467),
.B(n_5447),
.Y(n_6008)
);

BUFx2_ASAP7_75t_L g6009 ( 
.A(n_5044),
.Y(n_6009)
);

AOI22xp33_ASAP7_75t_SL g6010 ( 
.A1(n_5334),
.A2(n_4680),
.B1(n_4635),
.B2(n_4843),
.Y(n_6010)
);

OAI21xp5_ASAP7_75t_SL g6011 ( 
.A1(n_5503),
.A2(n_4536),
.B(n_4607),
.Y(n_6011)
);

OAI22xp5_ASAP7_75t_L g6012 ( 
.A1(n_5457),
.A2(n_4915),
.B1(n_4931),
.B2(n_4907),
.Y(n_6012)
);

AOI22xp33_ASAP7_75t_L g6013 ( 
.A1(n_5423),
.A2(n_4994),
.B1(n_4843),
.B2(n_4791),
.Y(n_6013)
);

OAI21xp33_ASAP7_75t_L g6014 ( 
.A1(n_5482),
.A2(n_4926),
.B(n_4594),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5619),
.Y(n_6015)
);

AND2x2_ASAP7_75t_L g6016 ( 
.A(n_5831),
.B(n_5159),
.Y(n_6016)
);

NAND2xp5_ASAP7_75t_L g6017 ( 
.A(n_5937),
.B(n_5205),
.Y(n_6017)
);

INVx2_ASAP7_75t_L g6018 ( 
.A(n_5814),
.Y(n_6018)
);

OAI21xp5_ASAP7_75t_L g6019 ( 
.A1(n_5573),
.A2(n_5356),
.B(n_5355),
.Y(n_6019)
);

AND2x2_ASAP7_75t_L g6020 ( 
.A(n_5831),
.B(n_5159),
.Y(n_6020)
);

INVx1_ASAP7_75t_L g6021 ( 
.A(n_5619),
.Y(n_6021)
);

OR2x2_ASAP7_75t_L g6022 ( 
.A(n_5781),
.B(n_5068),
.Y(n_6022)
);

INVx3_ASAP7_75t_L g6023 ( 
.A(n_5609),
.Y(n_6023)
);

INVx2_ASAP7_75t_L g6024 ( 
.A(n_5814),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5626),
.Y(n_6025)
);

AO21x2_ASAP7_75t_L g6026 ( 
.A1(n_5642),
.A2(n_5065),
.B(n_5322),
.Y(n_6026)
);

INVx3_ASAP7_75t_SL g6027 ( 
.A(n_5651),
.Y(n_6027)
);

AND2x4_ASAP7_75t_L g6028 ( 
.A(n_5730),
.B(n_5200),
.Y(n_6028)
);

BUFx6f_ASAP7_75t_L g6029 ( 
.A(n_5581),
.Y(n_6029)
);

INVx2_ASAP7_75t_L g6030 ( 
.A(n_5870),
.Y(n_6030)
);

HB1xp67_ASAP7_75t_L g6031 ( 
.A(n_5699),
.Y(n_6031)
);

OAI22xp5_ASAP7_75t_L g6032 ( 
.A1(n_5570),
.A2(n_5457),
.B1(n_5132),
.B2(n_5189),
.Y(n_6032)
);

INVxp67_ASAP7_75t_R g6033 ( 
.A(n_5686),
.Y(n_6033)
);

INVx1_ASAP7_75t_SL g6034 ( 
.A(n_5681),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5626),
.Y(n_6035)
);

AND2x4_ASAP7_75t_L g6036 ( 
.A(n_5730),
.B(n_5423),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5629),
.Y(n_6037)
);

INVx1_ASAP7_75t_L g6038 ( 
.A(n_5629),
.Y(n_6038)
);

INVx1_ASAP7_75t_L g6039 ( 
.A(n_5630),
.Y(n_6039)
);

INVx2_ASAP7_75t_SL g6040 ( 
.A(n_5806),
.Y(n_6040)
);

CKINVDCx5p33_ASAP7_75t_R g6041 ( 
.A(n_5715),
.Y(n_6041)
);

INVx2_ASAP7_75t_L g6042 ( 
.A(n_5870),
.Y(n_6042)
);

INVx2_ASAP7_75t_SL g6043 ( 
.A(n_5940),
.Y(n_6043)
);

AO21x2_ASAP7_75t_L g6044 ( 
.A1(n_5756),
.A2(n_5065),
.B(n_5322),
.Y(n_6044)
);

INVx1_ASAP7_75t_L g6045 ( 
.A(n_5630),
.Y(n_6045)
);

INVx2_ASAP7_75t_L g6046 ( 
.A(n_5965),
.Y(n_6046)
);

INVxp67_ASAP7_75t_L g6047 ( 
.A(n_5826),
.Y(n_6047)
);

INVx2_ASAP7_75t_SL g6048 ( 
.A(n_5940),
.Y(n_6048)
);

INVx1_ASAP7_75t_L g6049 ( 
.A(n_5636),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5965),
.Y(n_6050)
);

INVx2_ASAP7_75t_L g6051 ( 
.A(n_6001),
.Y(n_6051)
);

CKINVDCx5p33_ASAP7_75t_R g6052 ( 
.A(n_5715),
.Y(n_6052)
);

INVx5_ASAP7_75t_L g6053 ( 
.A(n_5633),
.Y(n_6053)
);

INVx2_ASAP7_75t_L g6054 ( 
.A(n_6001),
.Y(n_6054)
);

BUFx2_ASAP7_75t_L g6055 ( 
.A(n_5826),
.Y(n_6055)
);

NOR2x1_ASAP7_75t_L g6056 ( 
.A(n_5831),
.B(n_5322),
.Y(n_6056)
);

BUFx6f_ASAP7_75t_L g6057 ( 
.A(n_5581),
.Y(n_6057)
);

BUFx3_ASAP7_75t_L g6058 ( 
.A(n_5747),
.Y(n_6058)
);

AND2x2_ASAP7_75t_L g6059 ( 
.A(n_5788),
.B(n_5166),
.Y(n_6059)
);

INVx1_ASAP7_75t_L g6060 ( 
.A(n_5636),
.Y(n_6060)
);

INVx2_ASAP7_75t_L g6061 ( 
.A(n_6001),
.Y(n_6061)
);

INVx1_ASAP7_75t_L g6062 ( 
.A(n_5639),
.Y(n_6062)
);

AND2x2_ASAP7_75t_L g6063 ( 
.A(n_5788),
.B(n_5166),
.Y(n_6063)
);

INVx1_ASAP7_75t_L g6064 ( 
.A(n_5639),
.Y(n_6064)
);

BUFx8_ASAP7_75t_SL g6065 ( 
.A(n_5697),
.Y(n_6065)
);

OR2x2_ASAP7_75t_L g6066 ( 
.A(n_5837),
.B(n_5854),
.Y(n_6066)
);

INVx2_ASAP7_75t_L g6067 ( 
.A(n_6004),
.Y(n_6067)
);

AND2x2_ASAP7_75t_L g6068 ( 
.A(n_5833),
.B(n_5229),
.Y(n_6068)
);

INVx2_ASAP7_75t_L g6069 ( 
.A(n_6004),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_6004),
.Y(n_6070)
);

HB1xp67_ASAP7_75t_L g6071 ( 
.A(n_5719),
.Y(n_6071)
);

INVx1_ASAP7_75t_L g6072 ( 
.A(n_5653),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5653),
.Y(n_6073)
);

INVx1_ASAP7_75t_L g6074 ( 
.A(n_5662),
.Y(n_6074)
);

AOI21xp5_ASAP7_75t_SL g6075 ( 
.A1(n_5580),
.A2(n_5369),
.B(n_5364),
.Y(n_6075)
);

OA21x2_ASAP7_75t_L g6076 ( 
.A1(n_5845),
.A2(n_5555),
.B(n_5251),
.Y(n_6076)
);

INVx1_ASAP7_75t_L g6077 ( 
.A(n_5662),
.Y(n_6077)
);

HB1xp67_ASAP7_75t_L g6078 ( 
.A(n_5748),
.Y(n_6078)
);

INVx2_ASAP7_75t_SL g6079 ( 
.A(n_5940),
.Y(n_6079)
);

INVx5_ASAP7_75t_SL g6080 ( 
.A(n_5758),
.Y(n_6080)
);

INVx1_ASAP7_75t_L g6081 ( 
.A(n_5670),
.Y(n_6081)
);

INVx2_ASAP7_75t_L g6082 ( 
.A(n_5879),
.Y(n_6082)
);

OR2x2_ASAP7_75t_L g6083 ( 
.A(n_5909),
.B(n_5068),
.Y(n_6083)
);

BUFx2_ASAP7_75t_L g6084 ( 
.A(n_5731),
.Y(n_6084)
);

OR2x2_ASAP7_75t_L g6085 ( 
.A(n_5876),
.B(n_5068),
.Y(n_6085)
);

INVx2_ASAP7_75t_L g6086 ( 
.A(n_5879),
.Y(n_6086)
);

INVx2_ASAP7_75t_L g6087 ( 
.A(n_5906),
.Y(n_6087)
);

INVx2_ASAP7_75t_L g6088 ( 
.A(n_5906),
.Y(n_6088)
);

INVx4_ASAP7_75t_L g6089 ( 
.A(n_5747),
.Y(n_6089)
);

INVx2_ASAP7_75t_L g6090 ( 
.A(n_5910),
.Y(n_6090)
);

AO21x2_ASAP7_75t_L g6091 ( 
.A1(n_5810),
.A2(n_5070),
.B(n_5066),
.Y(n_6091)
);

INVx1_ASAP7_75t_L g6092 ( 
.A(n_5670),
.Y(n_6092)
);

INVx2_ASAP7_75t_L g6093 ( 
.A(n_5910),
.Y(n_6093)
);

NAND2xp5_ASAP7_75t_L g6094 ( 
.A(n_5674),
.B(n_5692),
.Y(n_6094)
);

OAI21x1_ASAP7_75t_L g6095 ( 
.A1(n_5920),
.A2(n_5149),
.B(n_5343),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_5675),
.Y(n_6096)
);

INVx1_ASAP7_75t_L g6097 ( 
.A(n_5675),
.Y(n_6097)
);

AOI21xp5_ASAP7_75t_L g6098 ( 
.A1(n_5568),
.A2(n_5760),
.B(n_5585),
.Y(n_6098)
);

AND2x4_ASAP7_75t_L g6099 ( 
.A(n_5730),
.B(n_5423),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_5833),
.B(n_5229),
.Y(n_6100)
);

AO21x2_ASAP7_75t_L g6101 ( 
.A1(n_5929),
.A2(n_5070),
.B(n_5066),
.Y(n_6101)
);

OAI21x1_ASAP7_75t_L g6102 ( 
.A1(n_5717),
.A2(n_5149),
.B(n_5343),
.Y(n_6102)
);

AND2x2_ASAP7_75t_L g6103 ( 
.A(n_5821),
.B(n_5238),
.Y(n_6103)
);

INVx2_ASAP7_75t_L g6104 ( 
.A(n_5904),
.Y(n_6104)
);

AND2x2_ASAP7_75t_L g6105 ( 
.A(n_5821),
.B(n_5238),
.Y(n_6105)
);

HB1xp67_ASAP7_75t_L g6106 ( 
.A(n_5685),
.Y(n_6106)
);

AO21x2_ASAP7_75t_L g6107 ( 
.A1(n_5934),
.A2(n_5101),
.B(n_5085),
.Y(n_6107)
);

OR2x2_ASAP7_75t_L g6108 ( 
.A(n_5798),
.B(n_5068),
.Y(n_6108)
);

AO21x2_ASAP7_75t_L g6109 ( 
.A1(n_5975),
.A2(n_5101),
.B(n_5085),
.Y(n_6109)
);

AO21x2_ASAP7_75t_L g6110 ( 
.A1(n_6011),
.A2(n_5139),
.B(n_5106),
.Y(n_6110)
);

INVx1_ASAP7_75t_L g6111 ( 
.A(n_5677),
.Y(n_6111)
);

INVx2_ASAP7_75t_SL g6112 ( 
.A(n_5940),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5904),
.Y(n_6113)
);

AO21x2_ASAP7_75t_L g6114 ( 
.A1(n_5659),
.A2(n_5139),
.B(n_5106),
.Y(n_6114)
);

INVx2_ASAP7_75t_L g6115 ( 
.A(n_5594),
.Y(n_6115)
);

AOI21xp5_ASAP7_75t_SL g6116 ( 
.A1(n_5731),
.A2(n_5334),
.B(n_5482),
.Y(n_6116)
);

INVx1_ASAP7_75t_L g6117 ( 
.A(n_5677),
.Y(n_6117)
);

AOI22xp33_ASAP7_75t_L g6118 ( 
.A1(n_5613),
.A2(n_5526),
.B1(n_5179),
.B2(n_5460),
.Y(n_6118)
);

AND2x2_ASAP7_75t_L g6119 ( 
.A(n_5732),
.B(n_5250),
.Y(n_6119)
);

INVx1_ASAP7_75t_L g6120 ( 
.A(n_5679),
.Y(n_6120)
);

INVx2_ASAP7_75t_L g6121 ( 
.A(n_5594),
.Y(n_6121)
);

BUFx2_ASAP7_75t_L g6122 ( 
.A(n_5731),
.Y(n_6122)
);

AND2x2_ASAP7_75t_L g6123 ( 
.A(n_5732),
.B(n_5250),
.Y(n_6123)
);

INVx1_ASAP7_75t_SL g6124 ( 
.A(n_5681),
.Y(n_6124)
);

BUFx3_ASAP7_75t_L g6125 ( 
.A(n_5754),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5679),
.Y(n_6126)
);

AO21x2_ASAP7_75t_L g6127 ( 
.A1(n_5742),
.A2(n_5165),
.B(n_5145),
.Y(n_6127)
);

INVx1_ASAP7_75t_L g6128 ( 
.A(n_5700),
.Y(n_6128)
);

AND2x2_ASAP7_75t_L g6129 ( 
.A(n_5738),
.B(n_5324),
.Y(n_6129)
);

HB1xp67_ASAP7_75t_L g6130 ( 
.A(n_5640),
.Y(n_6130)
);

BUFx2_ASAP7_75t_L g6131 ( 
.A(n_5794),
.Y(n_6131)
);

NAND2xp5_ASAP7_75t_L g6132 ( 
.A(n_5635),
.B(n_5205),
.Y(n_6132)
);

NAND2xp5_ASAP7_75t_L g6133 ( 
.A(n_5648),
.B(n_5324),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_5640),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_5738),
.B(n_5126),
.Y(n_6135)
);

HB1xp67_ASAP7_75t_L g6136 ( 
.A(n_5658),
.Y(n_6136)
);

BUFx3_ASAP7_75t_L g6137 ( 
.A(n_5754),
.Y(n_6137)
);

BUFx6f_ASAP7_75t_L g6138 ( 
.A(n_5663),
.Y(n_6138)
);

INVx1_ASAP7_75t_L g6139 ( 
.A(n_5700),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_5658),
.Y(n_6140)
);

HB1xp67_ASAP7_75t_L g6141 ( 
.A(n_5707),
.Y(n_6141)
);

INVx1_ASAP7_75t_L g6142 ( 
.A(n_5709),
.Y(n_6142)
);

INVx2_ASAP7_75t_L g6143 ( 
.A(n_5707),
.Y(n_6143)
);

INVx1_ASAP7_75t_L g6144 ( 
.A(n_5709),
.Y(n_6144)
);

AND2x2_ASAP7_75t_L g6145 ( 
.A(n_5851),
.B(n_5126),
.Y(n_6145)
);

AND2x4_ASAP7_75t_L g6146 ( 
.A(n_5625),
.B(n_5526),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_5712),
.Y(n_6147)
);

OAI21x1_ASAP7_75t_L g6148 ( 
.A1(n_5848),
.A2(n_5468),
.B(n_5558),
.Y(n_6148)
);

AOI21x1_ASAP7_75t_L g6149 ( 
.A1(n_5564),
.A2(n_5660),
.B(n_5632),
.Y(n_6149)
);

INVx2_ASAP7_75t_L g6150 ( 
.A(n_5708),
.Y(n_6150)
);

AND2x2_ASAP7_75t_L g6151 ( 
.A(n_5851),
.B(n_5126),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_5708),
.Y(n_6152)
);

AOI21x1_ASAP7_75t_L g6153 ( 
.A1(n_5564),
.A2(n_5468),
.B(n_5558),
.Y(n_6153)
);

INVx1_ASAP7_75t_L g6154 ( 
.A(n_5712),
.Y(n_6154)
);

NAND2xp5_ASAP7_75t_L g6155 ( 
.A(n_5872),
.B(n_5068),
.Y(n_6155)
);

HB1xp67_ASAP7_75t_L g6156 ( 
.A(n_5995),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5746),
.Y(n_6157)
);

INVx1_ASAP7_75t_L g6158 ( 
.A(n_5746),
.Y(n_6158)
);

AND2x2_ASAP7_75t_L g6159 ( 
.A(n_5852),
.B(n_5132),
.Y(n_6159)
);

OR2x2_ASAP7_75t_L g6160 ( 
.A(n_5977),
.B(n_5207),
.Y(n_6160)
);

INVx1_ASAP7_75t_L g6161 ( 
.A(n_5763),
.Y(n_6161)
);

INVx3_ASAP7_75t_L g6162 ( 
.A(n_5609),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_L g6163 ( 
.A(n_5562),
.B(n_5329),
.Y(n_6163)
);

INVx2_ASAP7_75t_L g6164 ( 
.A(n_5946),
.Y(n_6164)
);

OR2x6_ASAP7_75t_L g6165 ( 
.A(n_5632),
.B(n_5482),
.Y(n_6165)
);

AND2x2_ASAP7_75t_SL g6166 ( 
.A(n_5607),
.B(n_5334),
.Y(n_6166)
);

OR2x2_ASAP7_75t_SL g6167 ( 
.A(n_5603),
.B(n_5030),
.Y(n_6167)
);

AND2x4_ASAP7_75t_L g6168 ( 
.A(n_5625),
.B(n_5526),
.Y(n_6168)
);

INVx1_ASAP7_75t_L g6169 ( 
.A(n_5763),
.Y(n_6169)
);

AO21x2_ASAP7_75t_L g6170 ( 
.A1(n_5765),
.A2(n_5165),
.B(n_5145),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_5769),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_5769),
.Y(n_6172)
);

INVx2_ASAP7_75t_L g6173 ( 
.A(n_5946),
.Y(n_6173)
);

AO31x2_ASAP7_75t_L g6174 ( 
.A1(n_5587),
.A2(n_5184),
.A3(n_5199),
.B(n_5177),
.Y(n_6174)
);

HB1xp67_ASAP7_75t_L g6175 ( 
.A(n_5660),
.Y(n_6175)
);

INVx2_ASAP7_75t_L g6176 ( 
.A(n_5933),
.Y(n_6176)
);

INVx2_ASAP7_75t_L g6177 ( 
.A(n_5933),
.Y(n_6177)
);

NOR2xp33_ASAP7_75t_R g6178 ( 
.A(n_5705),
.B(n_4994),
.Y(n_6178)
);

INVx2_ASAP7_75t_L g6179 ( 
.A(n_5948),
.Y(n_6179)
);

AND2x2_ASAP7_75t_L g6180 ( 
.A(n_5852),
.B(n_5132),
.Y(n_6180)
);

AO21x2_ASAP7_75t_L g6181 ( 
.A1(n_6002),
.A2(n_5184),
.B(n_5177),
.Y(n_6181)
);

AO21x2_ASAP7_75t_L g6182 ( 
.A1(n_5646),
.A2(n_5218),
.B(n_5199),
.Y(n_6182)
);

BUFx6f_ASAP7_75t_L g6183 ( 
.A(n_5663),
.Y(n_6183)
);

INVx1_ASAP7_75t_L g6184 ( 
.A(n_5774),
.Y(n_6184)
);

NOR2xp33_ASAP7_75t_L g6185 ( 
.A(n_5606),
.B(n_5130),
.Y(n_6185)
);

OA21x2_ASAP7_75t_L g6186 ( 
.A1(n_5860),
.A2(n_5555),
.B(n_5251),
.Y(n_6186)
);

INVx2_ASAP7_75t_L g6187 ( 
.A(n_5948),
.Y(n_6187)
);

HB1xp67_ASAP7_75t_L g6188 ( 
.A(n_5563),
.Y(n_6188)
);

AO21x2_ASAP7_75t_L g6189 ( 
.A1(n_5755),
.A2(n_5227),
.B(n_5218),
.Y(n_6189)
);

AND2x2_ASAP7_75t_L g6190 ( 
.A(n_5855),
.B(n_5189),
.Y(n_6190)
);

CKINVDCx20_ASAP7_75t_R g6191 ( 
.A(n_5655),
.Y(n_6191)
);

OAI21xp5_ASAP7_75t_L g6192 ( 
.A1(n_5565),
.A2(n_5550),
.B(n_5282),
.Y(n_6192)
);

OAI21x1_ASAP7_75t_L g6193 ( 
.A1(n_5911),
.A2(n_5118),
.B(n_5103),
.Y(n_6193)
);

INVx3_ASAP7_75t_L g6194 ( 
.A(n_5940),
.Y(n_6194)
);

INVx2_ASAP7_75t_L g6195 ( 
.A(n_5892),
.Y(n_6195)
);

INVx1_ASAP7_75t_L g6196 ( 
.A(n_5774),
.Y(n_6196)
);

INVx1_ASAP7_75t_L g6197 ( 
.A(n_5776),
.Y(n_6197)
);

OA21x2_ASAP7_75t_L g6198 ( 
.A1(n_5972),
.A2(n_5241),
.B(n_5416),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_5776),
.Y(n_6199)
);

AO21x2_ASAP7_75t_L g6200 ( 
.A1(n_5843),
.A2(n_5248),
.B(n_5227),
.Y(n_6200)
);

NAND2xp5_ASAP7_75t_L g6201 ( 
.A(n_5567),
.B(n_5219),
.Y(n_6201)
);

AO21x2_ASAP7_75t_L g6202 ( 
.A1(n_5792),
.A2(n_5248),
.B(n_5460),
.Y(n_6202)
);

NOR2xp67_ASAP7_75t_L g6203 ( 
.A(n_5693),
.B(n_5463),
.Y(n_6203)
);

INVx2_ASAP7_75t_L g6204 ( 
.A(n_5892),
.Y(n_6204)
);

INVx3_ASAP7_75t_L g6205 ( 
.A(n_5952),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_5784),
.Y(n_6206)
);

AND2x4_ASAP7_75t_L g6207 ( 
.A(n_5625),
.B(n_5120),
.Y(n_6207)
);

INVx2_ASAP7_75t_L g6208 ( 
.A(n_5892),
.Y(n_6208)
);

OR2x2_ASAP7_75t_L g6209 ( 
.A(n_5791),
.B(n_5497),
.Y(n_6209)
);

AND2x4_ASAP7_75t_L g6210 ( 
.A(n_5982),
.B(n_5120),
.Y(n_6210)
);

INVx1_ASAP7_75t_L g6211 ( 
.A(n_5784),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_5785),
.Y(n_6212)
);

INVx1_ASAP7_75t_L g6213 ( 
.A(n_5785),
.Y(n_6213)
);

OAI21x1_ASAP7_75t_L g6214 ( 
.A1(n_5913),
.A2(n_5118),
.B(n_5103),
.Y(n_6214)
);

BUFx2_ASAP7_75t_L g6215 ( 
.A(n_5794),
.Y(n_6215)
);

INVxp67_ASAP7_75t_SL g6216 ( 
.A(n_5669),
.Y(n_6216)
);

INVx2_ASAP7_75t_L g6217 ( 
.A(n_5923),
.Y(n_6217)
);

HB1xp67_ASAP7_75t_L g6218 ( 
.A(n_5563),
.Y(n_6218)
);

CKINVDCx5p33_ASAP7_75t_R g6219 ( 
.A(n_5705),
.Y(n_6219)
);

HB1xp67_ASAP7_75t_L g6220 ( 
.A(n_5602),
.Y(n_6220)
);

INVx2_ASAP7_75t_L g6221 ( 
.A(n_5923),
.Y(n_6221)
);

HB1xp67_ASAP7_75t_L g6222 ( 
.A(n_5602),
.Y(n_6222)
);

INVx2_ASAP7_75t_L g6223 ( 
.A(n_5923),
.Y(n_6223)
);

INVx2_ASAP7_75t_L g6224 ( 
.A(n_5575),
.Y(n_6224)
);

AND2x4_ASAP7_75t_L g6225 ( 
.A(n_5982),
.B(n_5120),
.Y(n_6225)
);

BUFx2_ASAP7_75t_SL g6226 ( 
.A(n_5991),
.Y(n_6226)
);

AND2x2_ASAP7_75t_L g6227 ( 
.A(n_5855),
.B(n_5189),
.Y(n_6227)
);

HB1xp67_ASAP7_75t_L g6228 ( 
.A(n_5608),
.Y(n_6228)
);

AND2x2_ASAP7_75t_L g6229 ( 
.A(n_5900),
.B(n_5194),
.Y(n_6229)
);

INVx1_ASAP7_75t_L g6230 ( 
.A(n_5793),
.Y(n_6230)
);

AO21x2_ASAP7_75t_L g6231 ( 
.A1(n_5591),
.A2(n_5460),
.B(n_5344),
.Y(n_6231)
);

OR2x2_ASAP7_75t_L g6232 ( 
.A(n_5762),
.B(n_5505),
.Y(n_6232)
);

INVx1_ASAP7_75t_L g6233 ( 
.A(n_5793),
.Y(n_6233)
);

AOI21x1_ASAP7_75t_L g6234 ( 
.A1(n_5994),
.A2(n_5693),
.B(n_5949),
.Y(n_6234)
);

INVx1_ASAP7_75t_L g6235 ( 
.A(n_5803),
.Y(n_6235)
);

INVx2_ASAP7_75t_L g6236 ( 
.A(n_5575),
.Y(n_6236)
);

HB1xp67_ASAP7_75t_L g6237 ( 
.A(n_5608),
.Y(n_6237)
);

INVx3_ASAP7_75t_L g6238 ( 
.A(n_5952),
.Y(n_6238)
);

OAI21xp5_ASAP7_75t_L g6239 ( 
.A1(n_5576),
.A2(n_5282),
.B(n_5276),
.Y(n_6239)
);

AND2x2_ASAP7_75t_L g6240 ( 
.A(n_5900),
.B(n_5194),
.Y(n_6240)
);

AND2x2_ASAP7_75t_L g6241 ( 
.A(n_5902),
.B(n_5194),
.Y(n_6241)
);

INVx2_ASAP7_75t_L g6242 ( 
.A(n_5575),
.Y(n_6242)
);

INVx2_ASAP7_75t_L g6243 ( 
.A(n_5579),
.Y(n_6243)
);

INVx1_ASAP7_75t_L g6244 ( 
.A(n_5803),
.Y(n_6244)
);

CKINVDCx11_ASAP7_75t_R g6245 ( 
.A(n_5697),
.Y(n_6245)
);

NAND2xp5_ASAP7_75t_L g6246 ( 
.A(n_5727),
.B(n_5219),
.Y(n_6246)
);

INVx1_ASAP7_75t_L g6247 ( 
.A(n_5807),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5579),
.Y(n_6248)
);

AND2x2_ASAP7_75t_L g6249 ( 
.A(n_5902),
.B(n_5384),
.Y(n_6249)
);

HB1xp67_ASAP7_75t_L g6250 ( 
.A(n_5617),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_5579),
.Y(n_6251)
);

OA21x2_ASAP7_75t_L g6252 ( 
.A1(n_5560),
.A2(n_5241),
.B(n_5416),
.Y(n_6252)
);

INVx1_ASAP7_75t_L g6253 ( 
.A(n_5807),
.Y(n_6253)
);

BUFx2_ASAP7_75t_L g6254 ( 
.A(n_5905),
.Y(n_6254)
);

INVx2_ASAP7_75t_L g6255 ( 
.A(n_5993),
.Y(n_6255)
);

NAND2xp5_ASAP7_75t_L g6256 ( 
.A(n_6008),
.B(n_5255),
.Y(n_6256)
);

INVx3_ASAP7_75t_L g6257 ( 
.A(n_5952),
.Y(n_6257)
);

INVx1_ASAP7_75t_L g6258 ( 
.A(n_5838),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_5838),
.Y(n_6259)
);

AND2x4_ASAP7_75t_L g6260 ( 
.A(n_5994),
.B(n_5120),
.Y(n_6260)
);

OAI21xp5_ASAP7_75t_L g6261 ( 
.A1(n_5583),
.A2(n_5276),
.B(n_5294),
.Y(n_6261)
);

INVx3_ASAP7_75t_L g6262 ( 
.A(n_5952),
.Y(n_6262)
);

AO21x2_ASAP7_75t_L g6263 ( 
.A1(n_5611),
.A2(n_5344),
.B(n_5475),
.Y(n_6263)
);

NAND2xp5_ASAP7_75t_L g6264 ( 
.A(n_5631),
.B(n_5255),
.Y(n_6264)
);

NAND2xp5_ASAP7_75t_SL g6265 ( 
.A(n_5877),
.B(n_5463),
.Y(n_6265)
);

AND2x4_ASAP7_75t_L g6266 ( 
.A(n_5952),
.B(n_5120),
.Y(n_6266)
);

AO21x2_ASAP7_75t_L g6267 ( 
.A1(n_5947),
.A2(n_5475),
.B(n_5486),
.Y(n_6267)
);

HB1xp67_ASAP7_75t_L g6268 ( 
.A(n_5617),
.Y(n_6268)
);

INVxp67_ASAP7_75t_L g6269 ( 
.A(n_5669),
.Y(n_6269)
);

OA21x2_ASAP7_75t_L g6270 ( 
.A1(n_5560),
.A2(n_5487),
.B(n_5420),
.Y(n_6270)
);

NAND2xp5_ASAP7_75t_L g6271 ( 
.A(n_5986),
.B(n_5255),
.Y(n_6271)
);

INVx2_ASAP7_75t_L g6272 ( 
.A(n_5993),
.Y(n_6272)
);

INVxp67_ASAP7_75t_L g6273 ( 
.A(n_5669),
.Y(n_6273)
);

INVx3_ASAP7_75t_L g6274 ( 
.A(n_5991),
.Y(n_6274)
);

AND2x2_ASAP7_75t_L g6275 ( 
.A(n_5601),
.B(n_5847),
.Y(n_6275)
);

BUFx2_ASAP7_75t_SL g6276 ( 
.A(n_5991),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_6003),
.Y(n_6277)
);

INVx2_ASAP7_75t_L g6278 ( 
.A(n_6003),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_5780),
.Y(n_6279)
);

BUFx3_ASAP7_75t_L g6280 ( 
.A(n_5695),
.Y(n_6280)
);

INVx4_ASAP7_75t_SL g6281 ( 
.A(n_5706),
.Y(n_6281)
);

AND2x2_ASAP7_75t_L g6282 ( 
.A(n_5601),
.B(n_5187),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_5841),
.Y(n_6283)
);

AOI21xp5_ASAP7_75t_SL g6284 ( 
.A1(n_5753),
.A2(n_5522),
.B(n_5521),
.Y(n_6284)
);

OR2x6_ASAP7_75t_L g6285 ( 
.A(n_5758),
.B(n_5221),
.Y(n_6285)
);

INVx1_ASAP7_75t_L g6286 ( 
.A(n_5841),
.Y(n_6286)
);

INVx2_ASAP7_75t_SL g6287 ( 
.A(n_5669),
.Y(n_6287)
);

CKINVDCx6p67_ASAP7_75t_R g6288 ( 
.A(n_5569),
.Y(n_6288)
);

AND2x2_ASAP7_75t_L g6289 ( 
.A(n_5847),
.B(n_5757),
.Y(n_6289)
);

OA21x2_ASAP7_75t_L g6290 ( 
.A1(n_5577),
.A2(n_5487),
.B(n_5420),
.Y(n_6290)
);

BUFx6f_ASAP7_75t_L g6291 ( 
.A(n_5716),
.Y(n_6291)
);

INVx3_ASAP7_75t_L g6292 ( 
.A(n_5905),
.Y(n_6292)
);

INVx1_ASAP7_75t_L g6293 ( 
.A(n_5880),
.Y(n_6293)
);

INVx1_ASAP7_75t_L g6294 ( 
.A(n_5880),
.Y(n_6294)
);

HB1xp67_ASAP7_75t_L g6295 ( 
.A(n_5780),
.Y(n_6295)
);

INVx2_ASAP7_75t_L g6296 ( 
.A(n_5873),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_5891),
.Y(n_6297)
);

HB1xp67_ASAP7_75t_L g6298 ( 
.A(n_5873),
.Y(n_6298)
);

INVx2_ASAP7_75t_L g6299 ( 
.A(n_5884),
.Y(n_6299)
);

AOI21xp5_ASAP7_75t_SL g6300 ( 
.A1(n_5753),
.A2(n_5030),
.B(n_5162),
.Y(n_6300)
);

AND2x2_ASAP7_75t_L g6301 ( 
.A(n_5757),
.B(n_5187),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_5891),
.Y(n_6302)
);

OAI21xp5_ASAP7_75t_L g6303 ( 
.A1(n_5574),
.A2(n_5294),
.B(n_5253),
.Y(n_6303)
);

INVx2_ASAP7_75t_L g6304 ( 
.A(n_5884),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_5894),
.Y(n_6305)
);

BUFx4f_ASAP7_75t_L g6306 ( 
.A(n_5758),
.Y(n_6306)
);

OR2x2_ASAP7_75t_L g6307 ( 
.A(n_5762),
.B(n_5508),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_5901),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_5894),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_5759),
.B(n_5187),
.Y(n_6310)
);

INVx2_ASAP7_75t_L g6311 ( 
.A(n_5925),
.Y(n_6311)
);

BUFx3_ASAP7_75t_L g6312 ( 
.A(n_5695),
.Y(n_6312)
);

INVx1_ASAP7_75t_L g6313 ( 
.A(n_5901),
.Y(n_6313)
);

BUFx6f_ASAP7_75t_L g6314 ( 
.A(n_5716),
.Y(n_6314)
);

AND2x2_ASAP7_75t_L g6315 ( 
.A(n_5759),
.B(n_5187),
.Y(n_6315)
);

BUFx2_ASAP7_75t_L g6316 ( 
.A(n_5695),
.Y(n_6316)
);

AO21x2_ASAP7_75t_L g6317 ( 
.A1(n_5849),
.A2(n_5475),
.B(n_5486),
.Y(n_6317)
);

INVxp67_ASAP7_75t_L g6318 ( 
.A(n_5669),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_5779),
.B(n_5187),
.Y(n_6319)
);

OR2x6_ASAP7_75t_L g6320 ( 
.A(n_5758),
.B(n_5753),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5926),
.Y(n_6321)
);

AND2x2_ASAP7_75t_L g6322 ( 
.A(n_5779),
.B(n_5140),
.Y(n_6322)
);

HB1xp67_ASAP7_75t_L g6323 ( 
.A(n_5925),
.Y(n_6323)
);

AND2x2_ASAP7_75t_L g6324 ( 
.A(n_5779),
.B(n_5140),
.Y(n_6324)
);

AOI21x1_ASAP7_75t_L g6325 ( 
.A1(n_6009),
.A2(n_5412),
.B(n_5403),
.Y(n_6325)
);

OR2x2_ASAP7_75t_L g6326 ( 
.A(n_5778),
.B(n_5509),
.Y(n_6326)
);

INVx1_ASAP7_75t_L g6327 ( 
.A(n_5926),
.Y(n_6327)
);

AND2x2_ASAP7_75t_L g6328 ( 
.A(n_5779),
.B(n_5140),
.Y(n_6328)
);

OA21x2_ASAP7_75t_L g6329 ( 
.A1(n_5577),
.A2(n_5492),
.B(n_5232),
.Y(n_6329)
);

INVx1_ASAP7_75t_L g6330 ( 
.A(n_5951),
.Y(n_6330)
);

HB1xp67_ASAP7_75t_L g6331 ( 
.A(n_5865),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_5593),
.Y(n_6332)
);

INVx2_ASAP7_75t_L g6333 ( 
.A(n_5593),
.Y(n_6333)
);

OR2x2_ASAP7_75t_L g6334 ( 
.A(n_5778),
.B(n_5524),
.Y(n_6334)
);

NOR2xp33_ASAP7_75t_L g6335 ( 
.A(n_5582),
.B(n_5239),
.Y(n_6335)
);

INVx3_ASAP7_75t_L g6336 ( 
.A(n_5633),
.Y(n_6336)
);

AND2x2_ASAP7_75t_L g6337 ( 
.A(n_5865),
.B(n_5140),
.Y(n_6337)
);

BUFx2_ASAP7_75t_L g6338 ( 
.A(n_5701),
.Y(n_6338)
);

INVx1_ASAP7_75t_L g6339 ( 
.A(n_5951),
.Y(n_6339)
);

INVx2_ASAP7_75t_L g6340 ( 
.A(n_5593),
.Y(n_6340)
);

BUFx3_ASAP7_75t_L g6341 ( 
.A(n_5582),
.Y(n_6341)
);

AND2x2_ASAP7_75t_L g6342 ( 
.A(n_5804),
.B(n_5140),
.Y(n_6342)
);

INVx2_ASAP7_75t_L g6343 ( 
.A(n_5823),
.Y(n_6343)
);

AND2x2_ASAP7_75t_L g6344 ( 
.A(n_5804),
.B(n_5417),
.Y(n_6344)
);

INVx2_ASAP7_75t_L g6345 ( 
.A(n_5823),
.Y(n_6345)
);

HB1xp67_ASAP7_75t_L g6346 ( 
.A(n_5954),
.Y(n_6346)
);

INVx3_ASAP7_75t_L g6347 ( 
.A(n_5614),
.Y(n_6347)
);

OA21x2_ASAP7_75t_L g6348 ( 
.A1(n_5584),
.A2(n_5492),
.B(n_5232),
.Y(n_6348)
);

NAND2xp5_ASAP7_75t_L g6349 ( 
.A(n_5599),
.B(n_5255),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_5954),
.Y(n_6350)
);

INVx2_ASAP7_75t_L g6351 ( 
.A(n_5823),
.Y(n_6351)
);

INVx2_ASAP7_75t_L g6352 ( 
.A(n_5830),
.Y(n_6352)
);

AND2x2_ASAP7_75t_L g6353 ( 
.A(n_5953),
.B(n_5417),
.Y(n_6353)
);

INVx2_ASAP7_75t_L g6354 ( 
.A(n_5830),
.Y(n_6354)
);

INVx1_ASAP7_75t_L g6355 ( 
.A(n_5963),
.Y(n_6355)
);

AO21x2_ASAP7_75t_L g6356 ( 
.A1(n_5733),
.A2(n_5445),
.B(n_5444),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_5830),
.Y(n_6357)
);

OA21x2_ASAP7_75t_L g6358 ( 
.A1(n_5584),
.A2(n_5480),
.B(n_5556),
.Y(n_6358)
);

INVx2_ASAP7_75t_SL g6359 ( 
.A(n_5698),
.Y(n_6359)
);

INVx2_ASAP7_75t_L g6360 ( 
.A(n_5897),
.Y(n_6360)
);

AND2x2_ASAP7_75t_L g6361 ( 
.A(n_5953),
.B(n_5049),
.Y(n_6361)
);

AND2x2_ASAP7_75t_L g6362 ( 
.A(n_5888),
.B(n_5049),
.Y(n_6362)
);

AO21x2_ASAP7_75t_L g6363 ( 
.A1(n_6012),
.A2(n_5466),
.B(n_5448),
.Y(n_6363)
);

NAND2xp5_ASAP7_75t_L g6364 ( 
.A(n_5589),
.B(n_5255),
.Y(n_6364)
);

BUFx2_ASAP7_75t_L g6365 ( 
.A(n_5701),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_5963),
.Y(n_6366)
);

OR2x2_ASAP7_75t_L g6367 ( 
.A(n_5869),
.B(n_5525),
.Y(n_6367)
);

HB1xp67_ASAP7_75t_L g6368 ( 
.A(n_5964),
.Y(n_6368)
);

OA21x2_ASAP7_75t_L g6369 ( 
.A1(n_5596),
.A2(n_5480),
.B(n_5556),
.Y(n_6369)
);

OR2x2_ASAP7_75t_L g6370 ( 
.A(n_5869),
.B(n_5534),
.Y(n_6370)
);

INVx1_ASAP7_75t_L g6371 ( 
.A(n_5964),
.Y(n_6371)
);

INVx2_ASAP7_75t_L g6372 ( 
.A(n_5897),
.Y(n_6372)
);

AND2x2_ASAP7_75t_L g6373 ( 
.A(n_5888),
.B(n_5049),
.Y(n_6373)
);

BUFx12f_ASAP7_75t_L g6374 ( 
.A(n_5641),
.Y(n_6374)
);

AND2x4_ASAP7_75t_L g6375 ( 
.A(n_5962),
.B(n_5049),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_5971),
.Y(n_6376)
);

INVx1_ASAP7_75t_L g6377 ( 
.A(n_5971),
.Y(n_6377)
);

INVx1_ASAP7_75t_L g6378 ( 
.A(n_5984),
.Y(n_6378)
);

HB1xp67_ASAP7_75t_L g6379 ( 
.A(n_5984),
.Y(n_6379)
);

INVx1_ASAP7_75t_L g6380 ( 
.A(n_5987),
.Y(n_6380)
);

AO21x2_ASAP7_75t_L g6381 ( 
.A1(n_5921),
.A2(n_5592),
.B(n_5721),
.Y(n_6381)
);

AND2x2_ASAP7_75t_L g6382 ( 
.A(n_5790),
.B(n_5962),
.Y(n_6382)
);

INVx2_ASAP7_75t_L g6383 ( 
.A(n_5897),
.Y(n_6383)
);

AND2x2_ASAP7_75t_L g6384 ( 
.A(n_5790),
.B(n_5049),
.Y(n_6384)
);

BUFx4f_ASAP7_75t_SL g6385 ( 
.A(n_5655),
.Y(n_6385)
);

NAND2xp5_ASAP7_75t_L g6386 ( 
.A(n_5883),
.B(n_5877),
.Y(n_6386)
);

INVx2_ASAP7_75t_L g6387 ( 
.A(n_5973),
.Y(n_6387)
);

INVx2_ASAP7_75t_L g6388 ( 
.A(n_5973),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_5987),
.Y(n_6389)
);

AO21x2_ASAP7_75t_L g6390 ( 
.A1(n_5924),
.A2(n_5517),
.B(n_5502),
.Y(n_6390)
);

INVx2_ASAP7_75t_SL g6391 ( 
.A(n_5698),
.Y(n_6391)
);

AND2x2_ASAP7_75t_L g6392 ( 
.A(n_6009),
.B(n_5411),
.Y(n_6392)
);

INVx1_ASAP7_75t_L g6393 ( 
.A(n_5572),
.Y(n_6393)
);

OR2x6_ASAP7_75t_L g6394 ( 
.A(n_5758),
.B(n_5221),
.Y(n_6394)
);

INVx2_ASAP7_75t_L g6395 ( 
.A(n_5973),
.Y(n_6395)
);

OR2x2_ASAP7_75t_L g6396 ( 
.A(n_5835),
.B(n_5216),
.Y(n_6396)
);

INVx1_ASAP7_75t_L g6397 ( 
.A(n_5578),
.Y(n_6397)
);

HB1xp67_ASAP7_75t_L g6398 ( 
.A(n_6130),
.Y(n_6398)
);

INVx1_ASAP7_75t_L g6399 ( 
.A(n_6346),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6368),
.Y(n_6400)
);

NOR2xp33_ASAP7_75t_L g6401 ( 
.A(n_6041),
.B(n_5569),
.Y(n_6401)
);

AND2x4_ASAP7_75t_L g6402 ( 
.A(n_6053),
.B(n_5614),
.Y(n_6402)
);

BUFx6f_ASAP7_75t_L g6403 ( 
.A(n_6029),
.Y(n_6403)
);

AND2x2_ASAP7_75t_L g6404 ( 
.A(n_6016),
.B(n_5701),
.Y(n_6404)
);

NAND2xp5_ASAP7_75t_L g6405 ( 
.A(n_6098),
.B(n_5698),
.Y(n_6405)
);

NAND2xp5_ASAP7_75t_L g6406 ( 
.A(n_6216),
.B(n_5698),
.Y(n_6406)
);

OR2x2_ASAP7_75t_L g6407 ( 
.A(n_6066),
.B(n_5683),
.Y(n_6407)
);

BUFx3_ASAP7_75t_L g6408 ( 
.A(n_6029),
.Y(n_6408)
);

INVx2_ASAP7_75t_SL g6409 ( 
.A(n_6053),
.Y(n_6409)
);

NAND2xp5_ASAP7_75t_L g6410 ( 
.A(n_6269),
.B(n_5698),
.Y(n_6410)
);

AND2x2_ASAP7_75t_L g6411 ( 
.A(n_6016),
.B(n_5614),
.Y(n_6411)
);

BUFx12f_ASAP7_75t_L g6412 ( 
.A(n_6029),
.Y(n_6412)
);

INVx2_ASAP7_75t_L g6413 ( 
.A(n_6149),
.Y(n_6413)
);

INVx1_ASAP7_75t_SL g6414 ( 
.A(n_6385),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_6149),
.Y(n_6415)
);

AND2x2_ASAP7_75t_L g6416 ( 
.A(n_6020),
.B(n_5665),
.Y(n_6416)
);

INVx2_ASAP7_75t_L g6417 ( 
.A(n_6084),
.Y(n_6417)
);

INVx2_ASAP7_75t_L g6418 ( 
.A(n_6084),
.Y(n_6418)
);

INVx1_ASAP7_75t_L g6419 ( 
.A(n_6379),
.Y(n_6419)
);

INVxp67_ASAP7_75t_L g6420 ( 
.A(n_6055),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_L g6421 ( 
.A(n_6273),
.B(n_5739),
.Y(n_6421)
);

OR2x2_ASAP7_75t_L g6422 ( 
.A(n_6066),
.B(n_5714),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_6015),
.Y(n_6423)
);

OR2x6_ASAP7_75t_L g6424 ( 
.A(n_6226),
.B(n_5665),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_6020),
.B(n_5665),
.Y(n_6425)
);

AND2x2_ASAP7_75t_L g6426 ( 
.A(n_6353),
.B(n_5739),
.Y(n_6426)
);

AND2x2_ASAP7_75t_L g6427 ( 
.A(n_6353),
.B(n_5739),
.Y(n_6427)
);

NAND2xp5_ASAP7_75t_L g6428 ( 
.A(n_6318),
.B(n_5739),
.Y(n_6428)
);

AND2x2_ASAP7_75t_L g6429 ( 
.A(n_6289),
.B(n_6119),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_6015),
.Y(n_6430)
);

OR2x2_ASAP7_75t_L g6431 ( 
.A(n_6031),
.B(n_5724),
.Y(n_6431)
);

BUFx3_ASAP7_75t_L g6432 ( 
.A(n_6029),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_6021),
.Y(n_6433)
);

AND2x4_ASAP7_75t_L g6434 ( 
.A(n_6053),
.B(n_5633),
.Y(n_6434)
);

AND2x2_ASAP7_75t_L g6435 ( 
.A(n_6289),
.B(n_5739),
.Y(n_6435)
);

INVx1_ASAP7_75t_L g6436 ( 
.A(n_6021),
.Y(n_6436)
);

NAND2xp5_ASAP7_75t_L g6437 ( 
.A(n_6106),
.B(n_5740),
.Y(n_6437)
);

OR2x2_ASAP7_75t_L g6438 ( 
.A(n_6071),
.B(n_5735),
.Y(n_6438)
);

INVx1_ASAP7_75t_SL g6439 ( 
.A(n_6191),
.Y(n_6439)
);

INVx1_ASAP7_75t_L g6440 ( 
.A(n_6025),
.Y(n_6440)
);

INVx1_ASAP7_75t_L g6441 ( 
.A(n_6025),
.Y(n_6441)
);

NOR2xp67_ASAP7_75t_L g6442 ( 
.A(n_6047),
.B(n_5725),
.Y(n_6442)
);

AOI22xp33_ASAP7_75t_L g6443 ( 
.A1(n_6381),
.A2(n_5811),
.B1(n_5588),
.B2(n_5890),
.Y(n_6443)
);

AOI22xp33_ASAP7_75t_L g6444 ( 
.A1(n_6381),
.A2(n_5638),
.B1(n_5610),
.B2(n_5713),
.Y(n_6444)
);

AO21x2_ASAP7_75t_L g6445 ( 
.A1(n_6234),
.A2(n_5936),
.B(n_5924),
.Y(n_6445)
);

INVx2_ASAP7_75t_L g6446 ( 
.A(n_6122),
.Y(n_6446)
);

INVx1_ASAP7_75t_L g6447 ( 
.A(n_6035),
.Y(n_6447)
);

INVx2_ASAP7_75t_L g6448 ( 
.A(n_6122),
.Y(n_6448)
);

INVx2_ASAP7_75t_L g6449 ( 
.A(n_6194),
.Y(n_6449)
);

AND2x2_ASAP7_75t_L g6450 ( 
.A(n_6119),
.B(n_5740),
.Y(n_6450)
);

INVx1_ASAP7_75t_L g6451 ( 
.A(n_6035),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_6037),
.Y(n_6452)
);

INVx1_ASAP7_75t_L g6453 ( 
.A(n_6037),
.Y(n_6453)
);

NAND2xp5_ASAP7_75t_L g6454 ( 
.A(n_6078),
.B(n_5740),
.Y(n_6454)
);

CKINVDCx5p33_ASAP7_75t_R g6455 ( 
.A(n_6245),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6038),
.Y(n_6456)
);

NAND2xp5_ASAP7_75t_L g6457 ( 
.A(n_6136),
.B(n_5740),
.Y(n_6457)
);

INVx1_ASAP7_75t_L g6458 ( 
.A(n_6038),
.Y(n_6458)
);

HB1xp67_ASAP7_75t_L g6459 ( 
.A(n_6141),
.Y(n_6459)
);

INVx1_ASAP7_75t_L g6460 ( 
.A(n_6039),
.Y(n_6460)
);

HB1xp67_ASAP7_75t_L g6461 ( 
.A(n_6175),
.Y(n_6461)
);

OR2x2_ASAP7_75t_L g6462 ( 
.A(n_6018),
.B(n_5741),
.Y(n_6462)
);

OR2x2_ASAP7_75t_L g6463 ( 
.A(n_6018),
.B(n_5744),
.Y(n_6463)
);

INVx1_ASAP7_75t_L g6464 ( 
.A(n_6039),
.Y(n_6464)
);

INVx2_ASAP7_75t_L g6465 ( 
.A(n_6194),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_6156),
.B(n_5740),
.Y(n_6466)
);

INVx1_ASAP7_75t_L g6467 ( 
.A(n_6045),
.Y(n_6467)
);

AND2x2_ASAP7_75t_L g6468 ( 
.A(n_6123),
.B(n_5896),
.Y(n_6468)
);

INVx2_ASAP7_75t_L g6469 ( 
.A(n_6194),
.Y(n_6469)
);

OR2x2_ASAP7_75t_L g6470 ( 
.A(n_6024),
.B(n_6030),
.Y(n_6470)
);

INVx2_ASAP7_75t_L g6471 ( 
.A(n_6194),
.Y(n_6471)
);

AO21x2_ASAP7_75t_L g6472 ( 
.A1(n_6234),
.A2(n_5939),
.B(n_5936),
.Y(n_6472)
);

INVx2_ASAP7_75t_L g6473 ( 
.A(n_6205),
.Y(n_6473)
);

AOI22xp33_ASAP7_75t_L g6474 ( 
.A1(n_6381),
.A2(n_5782),
.B1(n_5856),
.B2(n_5612),
.Y(n_6474)
);

INVx1_ASAP7_75t_L g6475 ( 
.A(n_6045),
.Y(n_6475)
);

AND2x4_ASAP7_75t_L g6476 ( 
.A(n_6053),
.B(n_5633),
.Y(n_6476)
);

INVx2_ASAP7_75t_L g6477 ( 
.A(n_6205),
.Y(n_6477)
);

AND2x2_ASAP7_75t_L g6478 ( 
.A(n_6123),
.B(n_5652),
.Y(n_6478)
);

AND2x2_ASAP7_75t_L g6479 ( 
.A(n_6129),
.B(n_5989),
.Y(n_6479)
);

OR2x2_ASAP7_75t_L g6480 ( 
.A(n_6024),
.B(n_6030),
.Y(n_6480)
);

INVx2_ASAP7_75t_L g6481 ( 
.A(n_6205),
.Y(n_6481)
);

HB1xp67_ASAP7_75t_L g6482 ( 
.A(n_6042),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6129),
.B(n_5989),
.Y(n_6483)
);

INVx2_ASAP7_75t_L g6484 ( 
.A(n_6205),
.Y(n_6484)
);

INVx1_ASAP7_75t_L g6485 ( 
.A(n_6049),
.Y(n_6485)
);

AND2x4_ASAP7_75t_L g6486 ( 
.A(n_6053),
.B(n_5633),
.Y(n_6486)
);

AND2x4_ASAP7_75t_L g6487 ( 
.A(n_6053),
.B(n_5666),
.Y(n_6487)
);

AND2x4_ASAP7_75t_L g6488 ( 
.A(n_6023),
.B(n_5666),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_6238),
.Y(n_6489)
);

AND2x4_ASAP7_75t_L g6490 ( 
.A(n_6023),
.B(n_6162),
.Y(n_6490)
);

AND2x2_ASAP7_75t_L g6491 ( 
.A(n_6226),
.B(n_5864),
.Y(n_6491)
);

BUFx2_ASAP7_75t_L g6492 ( 
.A(n_6055),
.Y(n_6492)
);

NAND2xp5_ASAP7_75t_L g6493 ( 
.A(n_6094),
.B(n_5666),
.Y(n_6493)
);

INVx1_ASAP7_75t_L g6494 ( 
.A(n_6049),
.Y(n_6494)
);

AND2x2_ASAP7_75t_L g6495 ( 
.A(n_6276),
.B(n_5628),
.Y(n_6495)
);

AND2x2_ASAP7_75t_SL g6496 ( 
.A(n_6029),
.B(n_5666),
.Y(n_6496)
);

INVx1_ASAP7_75t_SL g6497 ( 
.A(n_6027),
.Y(n_6497)
);

AND2x4_ASAP7_75t_L g6498 ( 
.A(n_6023),
.B(n_5666),
.Y(n_6498)
);

INVxp67_ASAP7_75t_SL g6499 ( 
.A(n_6023),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_L g6500 ( 
.A(n_6162),
.B(n_5761),
.Y(n_6500)
);

BUFx3_ASAP7_75t_L g6501 ( 
.A(n_6057),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6238),
.Y(n_6502)
);

INVx1_ASAP7_75t_L g6503 ( 
.A(n_6060),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6060),
.Y(n_6504)
);

OR2x2_ASAP7_75t_L g6505 ( 
.A(n_6042),
.B(n_5812),
.Y(n_6505)
);

AND2x2_ASAP7_75t_L g6506 ( 
.A(n_6276),
.B(n_5899),
.Y(n_6506)
);

INVx2_ASAP7_75t_SL g6507 ( 
.A(n_6306),
.Y(n_6507)
);

INVx1_ASAP7_75t_L g6508 ( 
.A(n_6062),
.Y(n_6508)
);

NAND3xp33_ASAP7_75t_L g6509 ( 
.A(n_6019),
.B(n_5694),
.C(n_5956),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6062),
.Y(n_6510)
);

BUFx2_ASAP7_75t_L g6511 ( 
.A(n_6320),
.Y(n_6511)
);

INVx1_ASAP7_75t_L g6512 ( 
.A(n_6064),
.Y(n_6512)
);

INVx1_ASAP7_75t_L g6513 ( 
.A(n_6064),
.Y(n_6513)
);

INVx1_ASAP7_75t_L g6514 ( 
.A(n_6072),
.Y(n_6514)
);

INVx2_ASAP7_75t_L g6515 ( 
.A(n_6238),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_6072),
.Y(n_6516)
);

AND2x2_ASAP7_75t_L g6517 ( 
.A(n_6382),
.B(n_5696),
.Y(n_6517)
);

AND2x2_ASAP7_75t_L g6518 ( 
.A(n_6382),
.B(n_5916),
.Y(n_6518)
);

AND2x2_ASAP7_75t_L g6519 ( 
.A(n_6103),
.B(n_6105),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_6073),
.Y(n_6520)
);

BUFx2_ASAP7_75t_L g6521 ( 
.A(n_6320),
.Y(n_6521)
);

OR2x2_ASAP7_75t_L g6522 ( 
.A(n_6115),
.B(n_6121),
.Y(n_6522)
);

NAND2xp5_ASAP7_75t_L g6523 ( 
.A(n_6162),
.B(n_5775),
.Y(n_6523)
);

AND2x4_ASAP7_75t_L g6524 ( 
.A(n_6162),
.B(n_5818),
.Y(n_6524)
);

HB1xp67_ASAP7_75t_L g6525 ( 
.A(n_6331),
.Y(n_6525)
);

BUFx3_ASAP7_75t_L g6526 ( 
.A(n_6057),
.Y(n_6526)
);

INVx5_ASAP7_75t_L g6527 ( 
.A(n_6057),
.Y(n_6527)
);

AOI22xp33_ASAP7_75t_L g6528 ( 
.A1(n_6364),
.A2(n_5571),
.B1(n_5597),
.B2(n_5618),
.Y(n_6528)
);

HB1xp67_ASAP7_75t_L g6529 ( 
.A(n_6115),
.Y(n_6529)
);

NAND2xp5_ASAP7_75t_L g6530 ( 
.A(n_6121),
.B(n_5566),
.Y(n_6530)
);

AO21x2_ASAP7_75t_L g6531 ( 
.A1(n_6075),
.A2(n_5968),
.B(n_5939),
.Y(n_6531)
);

AND2x2_ASAP7_75t_L g6532 ( 
.A(n_6103),
.B(n_5918),
.Y(n_6532)
);

NOR2xp67_ASAP7_75t_L g6533 ( 
.A(n_6374),
.B(n_5720),
.Y(n_6533)
);

AND2x2_ASAP7_75t_L g6534 ( 
.A(n_6105),
.B(n_5919),
.Y(n_6534)
);

AND2x4_ASAP7_75t_L g6535 ( 
.A(n_6347),
.B(n_5822),
.Y(n_6535)
);

INVx4_ASAP7_75t_L g6536 ( 
.A(n_6057),
.Y(n_6536)
);

INVx2_ASAP7_75t_L g6537 ( 
.A(n_6257),
.Y(n_6537)
);

NAND2xp5_ASAP7_75t_L g6538 ( 
.A(n_6134),
.B(n_5682),
.Y(n_6538)
);

INVx3_ASAP7_75t_L g6539 ( 
.A(n_6057),
.Y(n_6539)
);

INVx2_ASAP7_75t_L g6540 ( 
.A(n_6257),
.Y(n_6540)
);

AND2x2_ASAP7_75t_L g6541 ( 
.A(n_6068),
.B(n_5672),
.Y(n_6541)
);

INVx1_ASAP7_75t_L g6542 ( 
.A(n_6073),
.Y(n_6542)
);

INVx1_ASAP7_75t_L g6543 ( 
.A(n_6074),
.Y(n_6543)
);

INVx2_ASAP7_75t_L g6544 ( 
.A(n_6257),
.Y(n_6544)
);

AND2x2_ASAP7_75t_L g6545 ( 
.A(n_6068),
.B(n_5668),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_6074),
.Y(n_6546)
);

AND2x4_ASAP7_75t_SL g6547 ( 
.A(n_6320),
.B(n_5912),
.Y(n_6547)
);

AND2x2_ASAP7_75t_L g6548 ( 
.A(n_6100),
.B(n_5615),
.Y(n_6548)
);

HB1xp67_ASAP7_75t_L g6549 ( 
.A(n_6134),
.Y(n_6549)
);

BUFx3_ASAP7_75t_L g6550 ( 
.A(n_6374),
.Y(n_6550)
);

NAND2xp5_ASAP7_75t_L g6551 ( 
.A(n_6140),
.B(n_5684),
.Y(n_6551)
);

AOI22xp33_ASAP7_75t_SL g6552 ( 
.A1(n_6201),
.A2(n_6166),
.B1(n_6182),
.B2(n_6361),
.Y(n_6552)
);

AND2x2_ASAP7_75t_L g6553 ( 
.A(n_6100),
.B(n_5942),
.Y(n_6553)
);

AO31x2_ASAP7_75t_L g6554 ( 
.A1(n_6338),
.A2(n_5893),
.A3(n_5832),
.B(n_5676),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_6275),
.B(n_6007),
.Y(n_6555)
);

INVx2_ASAP7_75t_L g6556 ( 
.A(n_6262),
.Y(n_6556)
);

NAND2xp5_ASAP7_75t_L g6557 ( 
.A(n_6140),
.B(n_5912),
.Y(n_6557)
);

NAND2xp5_ASAP7_75t_L g6558 ( 
.A(n_6143),
.B(n_5649),
.Y(n_6558)
);

OAI211xp5_ASAP7_75t_L g6559 ( 
.A1(n_6075),
.A2(n_5871),
.B(n_5914),
.C(n_5988),
.Y(n_6559)
);

INVxp67_ASAP7_75t_SL g6560 ( 
.A(n_6203),
.Y(n_6560)
);

NOR2xp33_ASAP7_75t_L g6561 ( 
.A(n_6041),
.B(n_5641),
.Y(n_6561)
);

AO21x2_ASAP7_75t_L g6562 ( 
.A1(n_6116),
.A2(n_5968),
.B(n_5903),
.Y(n_6562)
);

AND2x2_ASAP7_75t_L g6563 ( 
.A(n_6275),
.B(n_6135),
.Y(n_6563)
);

OAI22xp33_ASAP7_75t_L g6564 ( 
.A1(n_6033),
.A2(n_5595),
.B1(n_5604),
.B2(n_5598),
.Y(n_6564)
);

INVx3_ASAP7_75t_L g6565 ( 
.A(n_6028),
.Y(n_6565)
);

INVx2_ASAP7_75t_L g6566 ( 
.A(n_6262),
.Y(n_6566)
);

AND2x2_ASAP7_75t_L g6567 ( 
.A(n_6135),
.B(n_6007),
.Y(n_6567)
);

NOR4xp25_ASAP7_75t_SL g6568 ( 
.A(n_6265),
.B(n_5844),
.C(n_5889),
.D(n_5561),
.Y(n_6568)
);

AND2x2_ASAP7_75t_L g6569 ( 
.A(n_6344),
.B(n_5688),
.Y(n_6569)
);

INVx2_ASAP7_75t_L g6570 ( 
.A(n_6262),
.Y(n_6570)
);

INVxp67_ASAP7_75t_SL g6571 ( 
.A(n_6203),
.Y(n_6571)
);

INVx2_ASAP7_75t_L g6572 ( 
.A(n_6347),
.Y(n_6572)
);

AND2x2_ASAP7_75t_L g6573 ( 
.A(n_6344),
.B(n_5689),
.Y(n_6573)
);

OR2x2_ASAP7_75t_L g6574 ( 
.A(n_6143),
.B(n_5828),
.Y(n_6574)
);

OR2x2_ASAP7_75t_SL g6575 ( 
.A(n_6138),
.B(n_5895),
.Y(n_6575)
);

INVx1_ASAP7_75t_L g6576 ( 
.A(n_6077),
.Y(n_6576)
);

OR2x2_ASAP7_75t_L g6577 ( 
.A(n_6150),
.B(n_5836),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_6077),
.Y(n_6578)
);

INVx1_ASAP7_75t_SL g6579 ( 
.A(n_6027),
.Y(n_6579)
);

AND2x4_ASAP7_75t_L g6580 ( 
.A(n_6347),
.B(n_5857),
.Y(n_6580)
);

AND2x4_ASAP7_75t_L g6581 ( 
.A(n_6274),
.B(n_5907),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6081),
.Y(n_6582)
);

INVx1_ASAP7_75t_L g6583 ( 
.A(n_6081),
.Y(n_6583)
);

AND2x2_ASAP7_75t_L g6584 ( 
.A(n_6249),
.B(n_6059),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_L g6585 ( 
.A(n_6150),
.B(n_6000),
.Y(n_6585)
);

AND2x4_ASAP7_75t_L g6586 ( 
.A(n_6274),
.B(n_5917),
.Y(n_6586)
);

AND2x2_ASAP7_75t_L g6587 ( 
.A(n_6249),
.B(n_5690),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6092),
.Y(n_6588)
);

AND2x2_ASAP7_75t_L g6589 ( 
.A(n_6059),
.B(n_5703),
.Y(n_6589)
);

AND2x2_ASAP7_75t_L g6590 ( 
.A(n_6063),
.B(n_5970),
.Y(n_6590)
);

INVx2_ASAP7_75t_L g6591 ( 
.A(n_6336),
.Y(n_6591)
);

AND2x4_ASAP7_75t_L g6592 ( 
.A(n_6274),
.B(n_6287),
.Y(n_6592)
);

NOR2xp33_ASAP7_75t_L g6593 ( 
.A(n_6052),
.B(n_5561),
.Y(n_6593)
);

AND2x2_ASAP7_75t_L g6594 ( 
.A(n_6063),
.B(n_5997),
.Y(n_6594)
);

INVx1_ASAP7_75t_L g6595 ( 
.A(n_6092),
.Y(n_6595)
);

INVx2_ASAP7_75t_L g6596 ( 
.A(n_6336),
.Y(n_6596)
);

AOI22xp33_ASAP7_75t_L g6597 ( 
.A1(n_6131),
.A2(n_5764),
.B1(n_5605),
.B2(n_5616),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_L g6598 ( 
.A(n_6052),
.B(n_6065),
.Y(n_6598)
);

INVx1_ASAP7_75t_L g6599 ( 
.A(n_6096),
.Y(n_6599)
);

INVx2_ASAP7_75t_L g6600 ( 
.A(n_6336),
.Y(n_6600)
);

INVx1_ASAP7_75t_L g6601 ( 
.A(n_6096),
.Y(n_6601)
);

BUFx3_ASAP7_75t_L g6602 ( 
.A(n_6316),
.Y(n_6602)
);

AND2x4_ASAP7_75t_L g6603 ( 
.A(n_6274),
.B(n_5928),
.Y(n_6603)
);

NOR2xp33_ASAP7_75t_L g6604 ( 
.A(n_6027),
.B(n_5651),
.Y(n_6604)
);

AND2x2_ASAP7_75t_L g6605 ( 
.A(n_6229),
.B(n_5801),
.Y(n_6605)
);

INVx2_ASAP7_75t_L g6606 ( 
.A(n_6336),
.Y(n_6606)
);

INVx1_ASAP7_75t_L g6607 ( 
.A(n_6097),
.Y(n_6607)
);

AND2x2_ASAP7_75t_L g6608 ( 
.A(n_6229),
.B(n_5817),
.Y(n_6608)
);

INVx2_ASAP7_75t_L g6609 ( 
.A(n_6338),
.Y(n_6609)
);

INVx1_ASAP7_75t_L g6610 ( 
.A(n_6097),
.Y(n_6610)
);

INVx1_ASAP7_75t_L g6611 ( 
.A(n_6111),
.Y(n_6611)
);

HB1xp67_ASAP7_75t_L g6612 ( 
.A(n_6152),
.Y(n_6612)
);

OR2x2_ASAP7_75t_SL g6613 ( 
.A(n_6138),
.B(n_6183),
.Y(n_6613)
);

INVx1_ASAP7_75t_L g6614 ( 
.A(n_6111),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_6117),
.Y(n_6615)
);

INVx2_ASAP7_75t_SL g6616 ( 
.A(n_6306),
.Y(n_6616)
);

AO31x2_ASAP7_75t_L g6617 ( 
.A1(n_6365),
.A2(n_5825),
.A3(n_5667),
.B(n_5985),
.Y(n_6617)
);

AND2x2_ASAP7_75t_L g6618 ( 
.A(n_6240),
.B(n_5853),
.Y(n_6618)
);

INVx2_ASAP7_75t_L g6619 ( 
.A(n_6365),
.Y(n_6619)
);

NAND2xp5_ASAP7_75t_L g6620 ( 
.A(n_6152),
.B(n_5752),
.Y(n_6620)
);

BUFx2_ASAP7_75t_L g6621 ( 
.A(n_6320),
.Y(n_6621)
);

INVx2_ASAP7_75t_L g6622 ( 
.A(n_6287),
.Y(n_6622)
);

AND2x2_ASAP7_75t_L g6623 ( 
.A(n_6240),
.B(n_5941),
.Y(n_6623)
);

INVx1_ASAP7_75t_L g6624 ( 
.A(n_6117),
.Y(n_6624)
);

INVx2_ASAP7_75t_L g6625 ( 
.A(n_6359),
.Y(n_6625)
);

INVx2_ASAP7_75t_L g6626 ( 
.A(n_6359),
.Y(n_6626)
);

INVx2_ASAP7_75t_L g6627 ( 
.A(n_6391),
.Y(n_6627)
);

INVx3_ASAP7_75t_L g6628 ( 
.A(n_6028),
.Y(n_6628)
);

AND2x2_ASAP7_75t_L g6629 ( 
.A(n_6241),
.B(n_5827),
.Y(n_6629)
);

OAI21x1_ASAP7_75t_SL g6630 ( 
.A1(n_6153),
.A2(n_5704),
.B(n_5664),
.Y(n_6630)
);

INVx2_ASAP7_75t_L g6631 ( 
.A(n_6391),
.Y(n_6631)
);

NAND2xp5_ASAP7_75t_L g6632 ( 
.A(n_6043),
.B(n_5974),
.Y(n_6632)
);

AND2x2_ASAP7_75t_L g6633 ( 
.A(n_6241),
.B(n_5827),
.Y(n_6633)
);

INVx1_ASAP7_75t_L g6634 ( 
.A(n_6120),
.Y(n_6634)
);

INVx1_ASAP7_75t_L g6635 ( 
.A(n_6120),
.Y(n_6635)
);

AND2x2_ASAP7_75t_L g6636 ( 
.A(n_6145),
.B(n_6151),
.Y(n_6636)
);

INVx1_ASAP7_75t_L g6637 ( 
.A(n_6126),
.Y(n_6637)
);

NAND2xp5_ASAP7_75t_L g6638 ( 
.A(n_6043),
.B(n_5773),
.Y(n_6638)
);

AND2x4_ASAP7_75t_SL g6639 ( 
.A(n_6320),
.B(n_5654),
.Y(n_6639)
);

AND2x2_ASAP7_75t_L g6640 ( 
.A(n_6145),
.B(n_5960),
.Y(n_6640)
);

NOR4xp25_ASAP7_75t_SL g6641 ( 
.A(n_6254),
.B(n_5718),
.C(n_6014),
.D(n_5621),
.Y(n_6641)
);

INVx2_ASAP7_75t_L g6642 ( 
.A(n_6167),
.Y(n_6642)
);

NAND2xp5_ASAP7_75t_L g6643 ( 
.A(n_6048),
.B(n_5723),
.Y(n_6643)
);

AO21x2_ASAP7_75t_L g6644 ( 
.A1(n_6116),
.A2(n_5586),
.B(n_5596),
.Y(n_6644)
);

NAND2xp5_ASAP7_75t_L g6645 ( 
.A(n_6048),
.B(n_5983),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6126),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_6167),
.Y(n_6647)
);

OR2x2_ASAP7_75t_L g6648 ( 
.A(n_6160),
.B(n_5931),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_6128),
.Y(n_6649)
);

AND2x2_ASAP7_75t_L g6650 ( 
.A(n_6151),
.B(n_5960),
.Y(n_6650)
);

INVx1_ASAP7_75t_L g6651 ( 
.A(n_6128),
.Y(n_6651)
);

INVx5_ASAP7_75t_L g6652 ( 
.A(n_6089),
.Y(n_6652)
);

AND2x2_ASAP7_75t_L g6653 ( 
.A(n_6159),
.B(n_5960),
.Y(n_6653)
);

NAND2x1_ASAP7_75t_L g6654 ( 
.A(n_6284),
.B(n_5990),
.Y(n_6654)
);

BUFx3_ASAP7_75t_L g6655 ( 
.A(n_6316),
.Y(n_6655)
);

INVx2_ASAP7_75t_L g6656 ( 
.A(n_6079),
.Y(n_6656)
);

OAI31xp33_ASAP7_75t_L g6657 ( 
.A1(n_6032),
.A2(n_5938),
.A3(n_5815),
.B(n_5796),
.Y(n_6657)
);

OR2x2_ASAP7_75t_L g6658 ( 
.A(n_6160),
.B(n_5932),
.Y(n_6658)
);

AND2x2_ASAP7_75t_L g6659 ( 
.A(n_6159),
.B(n_5960),
.Y(n_6659)
);

NAND2xp5_ASAP7_75t_L g6660 ( 
.A(n_6079),
.B(n_5885),
.Y(n_6660)
);

INVx2_ASAP7_75t_L g6661 ( 
.A(n_6112),
.Y(n_6661)
);

OR2x2_ASAP7_75t_L g6662 ( 
.A(n_6164),
.B(n_6173),
.Y(n_6662)
);

AOI22xp33_ASAP7_75t_L g6663 ( 
.A1(n_6131),
.A2(n_5866),
.B1(n_5981),
.B2(n_5734),
.Y(n_6663)
);

AND2x2_ASAP7_75t_L g6664 ( 
.A(n_6180),
.B(n_5960),
.Y(n_6664)
);

AND2x2_ASAP7_75t_L g6665 ( 
.A(n_6180),
.B(n_5960),
.Y(n_6665)
);

AND2x2_ASAP7_75t_L g6666 ( 
.A(n_6190),
.B(n_5960),
.Y(n_6666)
);

AOI22xp33_ASAP7_75t_L g6667 ( 
.A1(n_6215),
.A2(n_5789),
.B1(n_5711),
.B2(n_5777),
.Y(n_6667)
);

NAND2xp5_ASAP7_75t_L g6668 ( 
.A(n_6112),
.B(n_6104),
.Y(n_6668)
);

AND2x2_ASAP7_75t_L g6669 ( 
.A(n_6190),
.B(n_5960),
.Y(n_6669)
);

AND2x4_ASAP7_75t_L g6670 ( 
.A(n_6040),
.B(n_5943),
.Y(n_6670)
);

NAND2x1p5_ASAP7_75t_L g6671 ( 
.A(n_6306),
.B(n_5643),
.Y(n_6671)
);

BUFx3_ASAP7_75t_L g6672 ( 
.A(n_6341),
.Y(n_6672)
);

INVx1_ASAP7_75t_L g6673 ( 
.A(n_6139),
.Y(n_6673)
);

AND2x2_ASAP7_75t_L g6674 ( 
.A(n_6227),
.B(n_5622),
.Y(n_6674)
);

AND2x2_ASAP7_75t_L g6675 ( 
.A(n_6227),
.B(n_5623),
.Y(n_6675)
);

HB1xp67_ASAP7_75t_L g6676 ( 
.A(n_6295),
.Y(n_6676)
);

INVx2_ASAP7_75t_L g6677 ( 
.A(n_6153),
.Y(n_6677)
);

INVx2_ASAP7_75t_SL g6678 ( 
.A(n_6028),
.Y(n_6678)
);

BUFx3_ASAP7_75t_L g6679 ( 
.A(n_6341),
.Y(n_6679)
);

OR2x2_ASAP7_75t_L g6680 ( 
.A(n_6164),
.B(n_5996),
.Y(n_6680)
);

BUFx3_ASAP7_75t_L g6681 ( 
.A(n_6341),
.Y(n_6681)
);

INVx2_ASAP7_75t_L g6682 ( 
.A(n_6181),
.Y(n_6682)
);

AND2x2_ASAP7_75t_L g6683 ( 
.A(n_6033),
.B(n_5624),
.Y(n_6683)
);

HB1xp67_ASAP7_75t_L g6684 ( 
.A(n_6298),
.Y(n_6684)
);

INVx2_ASAP7_75t_L g6685 ( 
.A(n_6181),
.Y(n_6685)
);

AND2x2_ASAP7_75t_L g6686 ( 
.A(n_6028),
.B(n_5678),
.Y(n_6686)
);

AND2x2_ASAP7_75t_L g6687 ( 
.A(n_6254),
.B(n_5680),
.Y(n_6687)
);

NAND2xp5_ASAP7_75t_L g6688 ( 
.A(n_6104),
.B(n_6113),
.Y(n_6688)
);

INVx1_ASAP7_75t_L g6689 ( 
.A(n_6139),
.Y(n_6689)
);

AND2x2_ASAP7_75t_L g6690 ( 
.A(n_6361),
.B(n_5957),
.Y(n_6690)
);

AND2x2_ASAP7_75t_L g6691 ( 
.A(n_6040),
.B(n_5656),
.Y(n_6691)
);

INVx1_ASAP7_75t_L g6692 ( 
.A(n_6142),
.Y(n_6692)
);

AO21x2_ASAP7_75t_L g6693 ( 
.A1(n_6284),
.A2(n_5620),
.B(n_5600),
.Y(n_6693)
);

BUFx2_ASAP7_75t_L g6694 ( 
.A(n_6280),
.Y(n_6694)
);

BUFx2_ASAP7_75t_L g6695 ( 
.A(n_6280),
.Y(n_6695)
);

INVx2_ASAP7_75t_L g6696 ( 
.A(n_6181),
.Y(n_6696)
);

BUFx3_ASAP7_75t_L g6697 ( 
.A(n_6280),
.Y(n_6697)
);

INVx1_ASAP7_75t_L g6698 ( 
.A(n_6142),
.Y(n_6698)
);

NAND2xp5_ASAP7_75t_L g6699 ( 
.A(n_6113),
.B(n_6335),
.Y(n_6699)
);

INVx1_ASAP7_75t_L g6700 ( 
.A(n_6144),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_6291),
.Y(n_6701)
);

AND2x2_ASAP7_75t_L g6702 ( 
.A(n_6392),
.B(n_5935),
.Y(n_6702)
);

INVx2_ASAP7_75t_L g6703 ( 
.A(n_6291),
.Y(n_6703)
);

NOR2xp33_ASAP7_75t_L g6704 ( 
.A(n_6089),
.B(n_5647),
.Y(n_6704)
);

AND2x2_ASAP7_75t_L g6705 ( 
.A(n_6392),
.B(n_5816),
.Y(n_6705)
);

INVx1_ASAP7_75t_L g6706 ( 
.A(n_6144),
.Y(n_6706)
);

AND2x2_ASAP7_75t_L g6707 ( 
.A(n_6173),
.B(n_5657),
.Y(n_6707)
);

AND2x2_ASAP7_75t_L g6708 ( 
.A(n_6215),
.B(n_5661),
.Y(n_6708)
);

AND2x2_ASAP7_75t_L g6709 ( 
.A(n_6292),
.B(n_5824),
.Y(n_6709)
);

BUFx6f_ASAP7_75t_L g6710 ( 
.A(n_6138),
.Y(n_6710)
);

AND2x2_ASAP7_75t_L g6711 ( 
.A(n_6292),
.B(n_5922),
.Y(n_6711)
);

OR2x2_ASAP7_75t_L g6712 ( 
.A(n_6017),
.B(n_6006),
.Y(n_6712)
);

AND2x2_ASAP7_75t_L g6713 ( 
.A(n_6292),
.B(n_5728),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_6147),
.Y(n_6714)
);

NAND3xp33_ASAP7_75t_SL g6715 ( 
.A(n_6256),
.B(n_5908),
.C(n_5858),
.Y(n_6715)
);

INVx1_ASAP7_75t_L g6716 ( 
.A(n_6147),
.Y(n_6716)
);

AND2x2_ASAP7_75t_L g6717 ( 
.A(n_6292),
.B(n_5944),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_6154),
.Y(n_6718)
);

OR2x6_ASAP7_75t_L g6719 ( 
.A(n_6312),
.B(n_5915),
.Y(n_6719)
);

INVx2_ASAP7_75t_L g6720 ( 
.A(n_6291),
.Y(n_6720)
);

AND2x2_ASAP7_75t_L g6721 ( 
.A(n_6176),
.B(n_5945),
.Y(n_6721)
);

INVx6_ASAP7_75t_L g6722 ( 
.A(n_6281),
.Y(n_6722)
);

AND2x4_ASAP7_75t_L g6723 ( 
.A(n_6176),
.B(n_5990),
.Y(n_6723)
);

NAND2xp5_ASAP7_75t_L g6724 ( 
.A(n_6188),
.B(n_5718),
.Y(n_6724)
);

INVxp67_ASAP7_75t_L g6725 ( 
.A(n_6291),
.Y(n_6725)
);

BUFx3_ASAP7_75t_L g6726 ( 
.A(n_6312),
.Y(n_6726)
);

INVx1_ASAP7_75t_L g6727 ( 
.A(n_6154),
.Y(n_6727)
);

HB1xp67_ASAP7_75t_L g6728 ( 
.A(n_6323),
.Y(n_6728)
);

AND2x2_ASAP7_75t_L g6729 ( 
.A(n_6177),
.B(n_5745),
.Y(n_6729)
);

AND2x2_ASAP7_75t_L g6730 ( 
.A(n_6177),
.B(n_5820),
.Y(n_6730)
);

INVxp67_ASAP7_75t_L g6731 ( 
.A(n_6291),
.Y(n_6731)
);

INVx1_ASAP7_75t_L g6732 ( 
.A(n_6157),
.Y(n_6732)
);

HB1xp67_ASAP7_75t_L g6733 ( 
.A(n_6218),
.Y(n_6733)
);

INVx1_ASAP7_75t_SL g6734 ( 
.A(n_6219),
.Y(n_6734)
);

BUFx3_ASAP7_75t_L g6735 ( 
.A(n_6312),
.Y(n_6735)
);

AND2x2_ASAP7_75t_L g6736 ( 
.A(n_6179),
.B(n_5766),
.Y(n_6736)
);

INVx2_ASAP7_75t_SL g6737 ( 
.A(n_6314),
.Y(n_6737)
);

INVx1_ASAP7_75t_L g6738 ( 
.A(n_6157),
.Y(n_6738)
);

BUFx2_ASAP7_75t_L g6739 ( 
.A(n_6178),
.Y(n_6739)
);

INVx1_ASAP7_75t_L g6740 ( 
.A(n_6158),
.Y(n_6740)
);

INVx1_ASAP7_75t_L g6741 ( 
.A(n_6158),
.Y(n_6741)
);

INVx1_ASAP7_75t_L g6742 ( 
.A(n_6161),
.Y(n_6742)
);

BUFx6f_ASAP7_75t_L g6743 ( 
.A(n_6138),
.Y(n_6743)
);

HB1xp67_ASAP7_75t_L g6744 ( 
.A(n_6220),
.Y(n_6744)
);

AND2x2_ASAP7_75t_L g6745 ( 
.A(n_6179),
.B(n_5767),
.Y(n_6745)
);

OR2x6_ASAP7_75t_L g6746 ( 
.A(n_6089),
.B(n_5691),
.Y(n_6746)
);

INVx2_ASAP7_75t_L g6747 ( 
.A(n_6314),
.Y(n_6747)
);

NAND2xp5_ASAP7_75t_L g6748 ( 
.A(n_6222),
.B(n_5867),
.Y(n_6748)
);

INVx1_ASAP7_75t_L g6749 ( 
.A(n_6161),
.Y(n_6749)
);

INVx2_ASAP7_75t_SL g6750 ( 
.A(n_6314),
.Y(n_6750)
);

INVx2_ASAP7_75t_L g6751 ( 
.A(n_6314),
.Y(n_6751)
);

AND2x4_ASAP7_75t_L g6752 ( 
.A(n_6187),
.B(n_5990),
.Y(n_6752)
);

HB1xp67_ASAP7_75t_L g6753 ( 
.A(n_6228),
.Y(n_6753)
);

INVx1_ASAP7_75t_L g6754 ( 
.A(n_6169),
.Y(n_6754)
);

BUFx3_ASAP7_75t_L g6755 ( 
.A(n_6058),
.Y(n_6755)
);

INVx2_ASAP7_75t_L g6756 ( 
.A(n_6314),
.Y(n_6756)
);

AO31x2_ASAP7_75t_L g6757 ( 
.A1(n_6195),
.A2(n_6204),
.A3(n_6217),
.B(n_6208),
.Y(n_6757)
);

BUFx3_ASAP7_75t_L g6758 ( 
.A(n_6058),
.Y(n_6758)
);

BUFx2_ASAP7_75t_L g6759 ( 
.A(n_6288),
.Y(n_6759)
);

INVx2_ASAP7_75t_L g6760 ( 
.A(n_6165),
.Y(n_6760)
);

INVx1_ASAP7_75t_L g6761 ( 
.A(n_6169),
.Y(n_6761)
);

OR2x2_ASAP7_75t_L g6762 ( 
.A(n_6237),
.B(n_5621),
.Y(n_6762)
);

INVx1_ASAP7_75t_L g6763 ( 
.A(n_6171),
.Y(n_6763)
);

HB1xp67_ASAP7_75t_L g6764 ( 
.A(n_6250),
.Y(n_6764)
);

HB1xp67_ASAP7_75t_L g6765 ( 
.A(n_6268),
.Y(n_6765)
);

INVx2_ASAP7_75t_L g6766 ( 
.A(n_6165),
.Y(n_6766)
);

INVx2_ASAP7_75t_L g6767 ( 
.A(n_6165),
.Y(n_6767)
);

OR2x2_ASAP7_75t_L g6768 ( 
.A(n_6255),
.B(n_5835),
.Y(n_6768)
);

INVx1_ASAP7_75t_L g6769 ( 
.A(n_6171),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6172),
.Y(n_6770)
);

AND2x4_ASAP7_75t_L g6771 ( 
.A(n_6492),
.B(n_6281),
.Y(n_6771)
);

INVxp67_ASAP7_75t_SL g6772 ( 
.A(n_6403),
.Y(n_6772)
);

NAND2xp5_ASAP7_75t_L g6773 ( 
.A(n_6492),
.B(n_6499),
.Y(n_6773)
);

INVx1_ASAP7_75t_L g6774 ( 
.A(n_6398),
.Y(n_6774)
);

INVx1_ASAP7_75t_L g6775 ( 
.A(n_6459),
.Y(n_6775)
);

BUFx3_ASAP7_75t_L g6776 ( 
.A(n_6412),
.Y(n_6776)
);

INVx2_ASAP7_75t_L g6777 ( 
.A(n_6682),
.Y(n_6777)
);

INVx1_ASAP7_75t_L g6778 ( 
.A(n_6733),
.Y(n_6778)
);

INVx1_ASAP7_75t_L g6779 ( 
.A(n_6744),
.Y(n_6779)
);

AND2x4_ASAP7_75t_L g6780 ( 
.A(n_6602),
.B(n_6281),
.Y(n_6780)
);

AND2x2_ASAP7_75t_L g6781 ( 
.A(n_6605),
.B(n_6080),
.Y(n_6781)
);

NAND2xp5_ASAP7_75t_L g6782 ( 
.A(n_6420),
.B(n_6034),
.Y(n_6782)
);

INVx1_ASAP7_75t_L g6783 ( 
.A(n_6753),
.Y(n_6783)
);

INVx1_ASAP7_75t_L g6784 ( 
.A(n_6764),
.Y(n_6784)
);

BUFx6f_ASAP7_75t_L g6785 ( 
.A(n_6403),
.Y(n_6785)
);

INVx2_ASAP7_75t_L g6786 ( 
.A(n_6682),
.Y(n_6786)
);

INVx3_ASAP7_75t_L g6787 ( 
.A(n_6412),
.Y(n_6787)
);

INVx1_ASAP7_75t_L g6788 ( 
.A(n_6765),
.Y(n_6788)
);

INVx2_ASAP7_75t_L g6789 ( 
.A(n_6685),
.Y(n_6789)
);

AND2x4_ASAP7_75t_L g6790 ( 
.A(n_6602),
.B(n_6281),
.Y(n_6790)
);

INVx2_ASAP7_75t_L g6791 ( 
.A(n_6685),
.Y(n_6791)
);

HB1xp67_ASAP7_75t_L g6792 ( 
.A(n_6655),
.Y(n_6792)
);

NAND2xp5_ASAP7_75t_L g6793 ( 
.A(n_6655),
.B(n_6124),
.Y(n_6793)
);

INVx3_ASAP7_75t_L g6794 ( 
.A(n_6536),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_6461),
.Y(n_6795)
);

AND2x2_ASAP7_75t_L g6796 ( 
.A(n_6605),
.B(n_6080),
.Y(n_6796)
);

AND2x2_ASAP7_75t_L g6797 ( 
.A(n_6426),
.B(n_6080),
.Y(n_6797)
);

INVx1_ASAP7_75t_L g6798 ( 
.A(n_6529),
.Y(n_6798)
);

INVx3_ASAP7_75t_L g6799 ( 
.A(n_6536),
.Y(n_6799)
);

AND2x2_ASAP7_75t_L g6800 ( 
.A(n_6426),
.B(n_6080),
.Y(n_6800)
);

INVx2_ASAP7_75t_L g6801 ( 
.A(n_6696),
.Y(n_6801)
);

NOR2xp67_ASAP7_75t_L g6802 ( 
.A(n_6527),
.B(n_6089),
.Y(n_6802)
);

AND2x4_ASAP7_75t_L g6803 ( 
.A(n_6678),
.B(n_6058),
.Y(n_6803)
);

BUFx2_ASAP7_75t_L g6804 ( 
.A(n_6455),
.Y(n_6804)
);

INVx1_ASAP7_75t_L g6805 ( 
.A(n_6549),
.Y(n_6805)
);

OR2x2_ASAP7_75t_L g6806 ( 
.A(n_6437),
.B(n_6132),
.Y(n_6806)
);

HB1xp67_ASAP7_75t_L g6807 ( 
.A(n_6525),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_6612),
.Y(n_6808)
);

NOR2xp33_ASAP7_75t_L g6809 ( 
.A(n_6455),
.B(n_6138),
.Y(n_6809)
);

INVx2_ASAP7_75t_L g6810 ( 
.A(n_6696),
.Y(n_6810)
);

OR2x2_ASAP7_75t_L g6811 ( 
.A(n_6643),
.B(n_6246),
.Y(n_6811)
);

INVxp67_ASAP7_75t_L g6812 ( 
.A(n_6759),
.Y(n_6812)
);

AND2x2_ASAP7_75t_L g6813 ( 
.A(n_6427),
.B(n_6288),
.Y(n_6813)
);

AO21x2_ASAP7_75t_L g6814 ( 
.A1(n_6642),
.A2(n_6091),
.B(n_6271),
.Y(n_6814)
);

NAND2xp5_ASAP7_75t_L g6815 ( 
.A(n_6725),
.B(n_6386),
.Y(n_6815)
);

INVx2_ASAP7_75t_L g6816 ( 
.A(n_6496),
.Y(n_6816)
);

BUFx2_ASAP7_75t_SL g6817 ( 
.A(n_6527),
.Y(n_6817)
);

AND2x2_ASAP7_75t_L g6818 ( 
.A(n_6427),
.B(n_6125),
.Y(n_6818)
);

NAND2xp5_ASAP7_75t_L g6819 ( 
.A(n_6731),
.B(n_6185),
.Y(n_6819)
);

BUFx2_ASAP7_75t_L g6820 ( 
.A(n_6759),
.Y(n_6820)
);

AND2x2_ASAP7_75t_L g6821 ( 
.A(n_6629),
.B(n_6125),
.Y(n_6821)
);

AND2x2_ASAP7_75t_L g6822 ( 
.A(n_6629),
.B(n_6125),
.Y(n_6822)
);

INVx3_ASAP7_75t_L g6823 ( 
.A(n_6536),
.Y(n_6823)
);

INVx2_ASAP7_75t_L g6824 ( 
.A(n_6496),
.Y(n_6824)
);

INVxp67_ASAP7_75t_SL g6825 ( 
.A(n_6403),
.Y(n_6825)
);

INVx2_ASAP7_75t_L g6826 ( 
.A(n_6408),
.Y(n_6826)
);

INVx2_ASAP7_75t_L g6827 ( 
.A(n_6408),
.Y(n_6827)
);

INVx1_ASAP7_75t_L g6828 ( 
.A(n_6482),
.Y(n_6828)
);

AND2x2_ASAP7_75t_L g6829 ( 
.A(n_6633),
.B(n_6137),
.Y(n_6829)
);

INVx1_ASAP7_75t_L g6830 ( 
.A(n_6676),
.Y(n_6830)
);

INVx2_ASAP7_75t_L g6831 ( 
.A(n_6432),
.Y(n_6831)
);

AND2x2_ASAP7_75t_L g6832 ( 
.A(n_6633),
.B(n_6137),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_6684),
.Y(n_6833)
);

INVx2_ASAP7_75t_L g6834 ( 
.A(n_6432),
.Y(n_6834)
);

INVx2_ASAP7_75t_L g6835 ( 
.A(n_6501),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6501),
.Y(n_6836)
);

INVx4_ASAP7_75t_L g6837 ( 
.A(n_6527),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6560),
.B(n_6187),
.Y(n_6838)
);

INVx2_ASAP7_75t_L g6839 ( 
.A(n_6526),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6435),
.B(n_6137),
.Y(n_6840)
);

AND2x2_ASAP7_75t_L g6841 ( 
.A(n_6435),
.B(n_6183),
.Y(n_6841)
);

INVx2_ASAP7_75t_L g6842 ( 
.A(n_6526),
.Y(n_6842)
);

NAND2xp5_ASAP7_75t_SL g6843 ( 
.A(n_6552),
.B(n_6509),
.Y(n_6843)
);

AND2x2_ASAP7_75t_L g6844 ( 
.A(n_6429),
.B(n_6183),
.Y(n_6844)
);

NOR2xp33_ASAP7_75t_L g6845 ( 
.A(n_6527),
.B(n_6183),
.Y(n_6845)
);

INVx4_ASAP7_75t_R g6846 ( 
.A(n_6550),
.Y(n_6846)
);

INVx2_ASAP7_75t_L g6847 ( 
.A(n_6403),
.Y(n_6847)
);

INVxp67_ASAP7_75t_L g6848 ( 
.A(n_6694),
.Y(n_6848)
);

INVx2_ASAP7_75t_L g6849 ( 
.A(n_6539),
.Y(n_6849)
);

NAND2x1p5_ASAP7_75t_L g6850 ( 
.A(n_6527),
.B(n_6183),
.Y(n_6850)
);

INVx2_ASAP7_75t_L g6851 ( 
.A(n_6539),
.Y(n_6851)
);

AND2x2_ASAP7_75t_L g6852 ( 
.A(n_6429),
.B(n_6182),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_6728),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6522),
.Y(n_6854)
);

AND2x4_ASAP7_75t_L g6855 ( 
.A(n_6678),
.B(n_6195),
.Y(n_6855)
);

AND2x2_ASAP7_75t_L g6856 ( 
.A(n_6563),
.B(n_6519),
.Y(n_6856)
);

BUFx3_ASAP7_75t_L g6857 ( 
.A(n_6613),
.Y(n_6857)
);

INVx1_ASAP7_75t_L g6858 ( 
.A(n_6522),
.Y(n_6858)
);

INVx3_ASAP7_75t_L g6859 ( 
.A(n_6654),
.Y(n_6859)
);

NAND2xp5_ASAP7_75t_SL g6860 ( 
.A(n_6474),
.B(n_6118),
.Y(n_6860)
);

AND2x2_ASAP7_75t_L g6861 ( 
.A(n_6563),
.B(n_6182),
.Y(n_6861)
);

OR2x2_ASAP7_75t_L g6862 ( 
.A(n_6466),
.B(n_6133),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6470),
.Y(n_6863)
);

AND2x2_ASAP7_75t_L g6864 ( 
.A(n_6519),
.B(n_6204),
.Y(n_6864)
);

OR2x2_ASAP7_75t_L g6865 ( 
.A(n_6688),
.B(n_6163),
.Y(n_6865)
);

BUFx3_ASAP7_75t_L g6866 ( 
.A(n_6613),
.Y(n_6866)
);

NAND2xp5_ASAP7_75t_L g6867 ( 
.A(n_6571),
.B(n_6208),
.Y(n_6867)
);

INVx3_ASAP7_75t_L g6868 ( 
.A(n_6539),
.Y(n_6868)
);

OR2x2_ASAP7_75t_L g6869 ( 
.A(n_6454),
.B(n_6174),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_6470),
.Y(n_6870)
);

INVx1_ASAP7_75t_L g6871 ( 
.A(n_6480),
.Y(n_6871)
);

INVxp67_ASAP7_75t_L g6872 ( 
.A(n_6694),
.Y(n_6872)
);

INVx1_ASAP7_75t_SL g6873 ( 
.A(n_6547),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6480),
.Y(n_6874)
);

NAND2xp5_ASAP7_75t_SL g6875 ( 
.A(n_6564),
.B(n_6166),
.Y(n_6875)
);

INVx2_ASAP7_75t_L g6876 ( 
.A(n_6565),
.Y(n_6876)
);

AND2x2_ASAP7_75t_L g6877 ( 
.A(n_6450),
.B(n_6217),
.Y(n_6877)
);

INVx2_ASAP7_75t_L g6878 ( 
.A(n_6565),
.Y(n_6878)
);

AND2x2_ASAP7_75t_L g6879 ( 
.A(n_6450),
.B(n_6221),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_6662),
.Y(n_6880)
);

NAND2xp5_ASAP7_75t_L g6881 ( 
.A(n_6695),
.B(n_6221),
.Y(n_6881)
);

AND2x2_ASAP7_75t_L g6882 ( 
.A(n_6584),
.B(n_6223),
.Y(n_6882)
);

INVx1_ASAP7_75t_L g6883 ( 
.A(n_6662),
.Y(n_6883)
);

INVx1_ASAP7_75t_L g6884 ( 
.A(n_6462),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6584),
.B(n_6223),
.Y(n_6885)
);

INVx1_ASAP7_75t_L g6886 ( 
.A(n_6462),
.Y(n_6886)
);

INVx1_ASAP7_75t_L g6887 ( 
.A(n_6463),
.Y(n_6887)
);

NAND2xp5_ASAP7_75t_L g6888 ( 
.A(n_6695),
.B(n_6279),
.Y(n_6888)
);

AND2x2_ASAP7_75t_L g6889 ( 
.A(n_6411),
.B(n_6279),
.Y(n_6889)
);

INVx1_ASAP7_75t_L g6890 ( 
.A(n_6463),
.Y(n_6890)
);

INVx1_ASAP7_75t_L g6891 ( 
.A(n_6505),
.Y(n_6891)
);

OR2x2_ASAP7_75t_SL g6892 ( 
.A(n_6500),
.B(n_6085),
.Y(n_6892)
);

INVx1_ASAP7_75t_L g6893 ( 
.A(n_6505),
.Y(n_6893)
);

AND2x2_ASAP7_75t_L g6894 ( 
.A(n_6411),
.B(n_6416),
.Y(n_6894)
);

AND2x2_ASAP7_75t_L g6895 ( 
.A(n_6416),
.B(n_6296),
.Y(n_6895)
);

NAND2xp5_ASAP7_75t_L g6896 ( 
.A(n_6490),
.B(n_6296),
.Y(n_6896)
);

AND2x2_ASAP7_75t_L g6897 ( 
.A(n_6425),
.B(n_6299),
.Y(n_6897)
);

AND2x2_ASAP7_75t_L g6898 ( 
.A(n_6425),
.B(n_6299),
.Y(n_6898)
);

INVx1_ASAP7_75t_L g6899 ( 
.A(n_6417),
.Y(n_6899)
);

INVx1_ASAP7_75t_L g6900 ( 
.A(n_6417),
.Y(n_6900)
);

INVx3_ASAP7_75t_L g6901 ( 
.A(n_6592),
.Y(n_6901)
);

INVx1_ASAP7_75t_L g6902 ( 
.A(n_6418),
.Y(n_6902)
);

AND2x2_ASAP7_75t_L g6903 ( 
.A(n_6636),
.B(n_6304),
.Y(n_6903)
);

INVx2_ASAP7_75t_L g6904 ( 
.A(n_6565),
.Y(n_6904)
);

OR2x2_ASAP7_75t_L g6905 ( 
.A(n_6418),
.B(n_6091),
.Y(n_6905)
);

INVx1_ASAP7_75t_L g6906 ( 
.A(n_6446),
.Y(n_6906)
);

INVx2_ASAP7_75t_L g6907 ( 
.A(n_6628),
.Y(n_6907)
);

INVx2_ASAP7_75t_L g6908 ( 
.A(n_6628),
.Y(n_6908)
);

AND2x2_ASAP7_75t_L g6909 ( 
.A(n_6636),
.B(n_6304),
.Y(n_6909)
);

AND2x2_ASAP7_75t_L g6910 ( 
.A(n_6404),
.B(n_6305),
.Y(n_6910)
);

HB1xp67_ASAP7_75t_L g6911 ( 
.A(n_6446),
.Y(n_6911)
);

INVx2_ASAP7_75t_L g6912 ( 
.A(n_6628),
.Y(n_6912)
);

HB1xp67_ASAP7_75t_L g6913 ( 
.A(n_6448),
.Y(n_6913)
);

AND2x2_ASAP7_75t_L g6914 ( 
.A(n_6404),
.B(n_6305),
.Y(n_6914)
);

AND2x2_ASAP7_75t_L g6915 ( 
.A(n_6479),
.B(n_6309),
.Y(n_6915)
);

AND2x2_ASAP7_75t_L g6916 ( 
.A(n_6479),
.B(n_6309),
.Y(n_6916)
);

OR2x2_ASAP7_75t_L g6917 ( 
.A(n_6405),
.B(n_6174),
.Y(n_6917)
);

BUFx3_ASAP7_75t_L g6918 ( 
.A(n_6550),
.Y(n_6918)
);

INVx1_ASAP7_75t_L g6919 ( 
.A(n_6448),
.Y(n_6919)
);

OR2x2_ASAP7_75t_L g6920 ( 
.A(n_6406),
.B(n_6174),
.Y(n_6920)
);

INVx1_ASAP7_75t_L g6921 ( 
.A(n_6609),
.Y(n_6921)
);

INVx2_ASAP7_75t_L g6922 ( 
.A(n_6693),
.Y(n_6922)
);

INVx1_ASAP7_75t_L g6923 ( 
.A(n_6609),
.Y(n_6923)
);

INVx2_ASAP7_75t_L g6924 ( 
.A(n_6693),
.Y(n_6924)
);

INVxp67_ASAP7_75t_L g6925 ( 
.A(n_6710),
.Y(n_6925)
);

HB1xp67_ASAP7_75t_L g6926 ( 
.A(n_6737),
.Y(n_6926)
);

INVx1_ASAP7_75t_L g6927 ( 
.A(n_6619),
.Y(n_6927)
);

NAND2x1_ASAP7_75t_L g6928 ( 
.A(n_6424),
.B(n_6434),
.Y(n_6928)
);

HB1xp67_ASAP7_75t_L g6929 ( 
.A(n_6737),
.Y(n_6929)
);

INVx4_ASAP7_75t_L g6930 ( 
.A(n_6652),
.Y(n_6930)
);

BUFx6f_ASAP7_75t_L g6931 ( 
.A(n_6710),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6619),
.Y(n_6932)
);

INVx2_ASAP7_75t_L g6933 ( 
.A(n_6693),
.Y(n_6933)
);

INVxp67_ASAP7_75t_SL g6934 ( 
.A(n_6523),
.Y(n_6934)
);

AND2x4_ASAP7_75t_L g6935 ( 
.A(n_6592),
.B(n_6311),
.Y(n_6935)
);

AND2x2_ASAP7_75t_L g6936 ( 
.A(n_6483),
.B(n_6311),
.Y(n_6936)
);

HB1xp67_ASAP7_75t_L g6937 ( 
.A(n_6750),
.Y(n_6937)
);

NAND2xp5_ASAP7_75t_L g6938 ( 
.A(n_6490),
.B(n_6200),
.Y(n_6938)
);

OAI22xp5_ASAP7_75t_L g6939 ( 
.A1(n_6444),
.A2(n_5858),
.B1(n_6166),
.B2(n_5887),
.Y(n_6939)
);

BUFx2_ASAP7_75t_L g6940 ( 
.A(n_6424),
.Y(n_6940)
);

INVx1_ASAP7_75t_SL g6941 ( 
.A(n_6547),
.Y(n_6941)
);

INVxp67_ASAP7_75t_L g6942 ( 
.A(n_6710),
.Y(n_6942)
);

INVx1_ASAP7_75t_L g6943 ( 
.A(n_6423),
.Y(n_6943)
);

HB1xp67_ASAP7_75t_L g6944 ( 
.A(n_6750),
.Y(n_6944)
);

AND2x2_ASAP7_75t_L g6945 ( 
.A(n_6483),
.B(n_6046),
.Y(n_6945)
);

BUFx3_ASAP7_75t_L g6946 ( 
.A(n_6672),
.Y(n_6946)
);

AND2x2_ASAP7_75t_L g6947 ( 
.A(n_6639),
.B(n_6046),
.Y(n_6947)
);

HB1xp67_ASAP7_75t_L g6948 ( 
.A(n_6511),
.Y(n_6948)
);

BUFx6f_ASAP7_75t_L g6949 ( 
.A(n_6710),
.Y(n_6949)
);

BUFx3_ASAP7_75t_L g6950 ( 
.A(n_6672),
.Y(n_6950)
);

AOI221xp5_ASAP7_75t_SL g6951 ( 
.A1(n_6443),
.A2(n_6192),
.B1(n_6303),
.B2(n_6261),
.C(n_6239),
.Y(n_6951)
);

INVx1_ASAP7_75t_L g6952 ( 
.A(n_6430),
.Y(n_6952)
);

AND2x2_ASAP7_75t_SL g6953 ( 
.A(n_6639),
.B(n_6085),
.Y(n_6953)
);

NAND2xp5_ASAP7_75t_L g6954 ( 
.A(n_6490),
.B(n_6200),
.Y(n_6954)
);

NAND2xp5_ASAP7_75t_L g6955 ( 
.A(n_6439),
.B(n_6200),
.Y(n_6955)
);

HB1xp67_ASAP7_75t_L g6956 ( 
.A(n_6511),
.Y(n_6956)
);

INVx2_ASAP7_75t_L g6957 ( 
.A(n_6424),
.Y(n_6957)
);

HB1xp67_ASAP7_75t_L g6958 ( 
.A(n_6521),
.Y(n_6958)
);

NAND2xp5_ASAP7_75t_L g6959 ( 
.A(n_6701),
.B(n_6255),
.Y(n_6959)
);

AO21x2_ASAP7_75t_L g6960 ( 
.A1(n_6642),
.A2(n_6647),
.B(n_6715),
.Y(n_6960)
);

AND2x2_ASAP7_75t_L g6961 ( 
.A(n_6618),
.B(n_6050),
.Y(n_6961)
);

AND2x2_ASAP7_75t_L g6962 ( 
.A(n_6618),
.B(n_6050),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_6433),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_6424),
.Y(n_6964)
);

INVx1_ASAP7_75t_L g6965 ( 
.A(n_6436),
.Y(n_6965)
);

AND2x2_ASAP7_75t_L g6966 ( 
.A(n_6545),
.B(n_6491),
.Y(n_6966)
);

INVx1_ASAP7_75t_L g6967 ( 
.A(n_6440),
.Y(n_6967)
);

AND2x2_ASAP7_75t_L g6968 ( 
.A(n_6545),
.B(n_6036),
.Y(n_6968)
);

NAND2xp5_ASAP7_75t_L g6969 ( 
.A(n_6701),
.B(n_6272),
.Y(n_6969)
);

AND2x2_ASAP7_75t_L g6970 ( 
.A(n_6491),
.B(n_6036),
.Y(n_6970)
);

INVx3_ASAP7_75t_L g6971 ( 
.A(n_6592),
.Y(n_6971)
);

AND2x2_ASAP7_75t_L g6972 ( 
.A(n_6590),
.B(n_6036),
.Y(n_6972)
);

INVx2_ASAP7_75t_L g6973 ( 
.A(n_6679),
.Y(n_6973)
);

OR2x2_ASAP7_75t_L g6974 ( 
.A(n_6575),
.B(n_6091),
.Y(n_6974)
);

OR2x2_ASAP7_75t_L g6975 ( 
.A(n_6638),
.B(n_6174),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6590),
.B(n_6036),
.Y(n_6976)
);

INVx2_ASAP7_75t_L g6977 ( 
.A(n_6679),
.Y(n_6977)
);

INVx2_ASAP7_75t_L g6978 ( 
.A(n_6681),
.Y(n_6978)
);

INVx2_ASAP7_75t_L g6979 ( 
.A(n_6681),
.Y(n_6979)
);

INVx1_ASAP7_75t_L g6980 ( 
.A(n_6441),
.Y(n_6980)
);

OR2x2_ASAP7_75t_L g6981 ( 
.A(n_6575),
.B(n_6272),
.Y(n_6981)
);

OR2x2_ASAP7_75t_L g6982 ( 
.A(n_6762),
.B(n_6277),
.Y(n_6982)
);

AND2x2_ASAP7_75t_L g6983 ( 
.A(n_6478),
.B(n_6506),
.Y(n_6983)
);

INVx2_ASAP7_75t_L g6984 ( 
.A(n_6521),
.Y(n_6984)
);

HB1xp67_ASAP7_75t_L g6985 ( 
.A(n_6621),
.Y(n_6985)
);

INVx2_ASAP7_75t_L g6986 ( 
.A(n_6621),
.Y(n_6986)
);

INVx1_ASAP7_75t_L g6987 ( 
.A(n_6447),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6451),
.Y(n_6988)
);

INVx2_ASAP7_75t_SL g6989 ( 
.A(n_6722),
.Y(n_6989)
);

INVx2_ASAP7_75t_SL g6990 ( 
.A(n_6722),
.Y(n_6990)
);

INVx2_ASAP7_75t_L g6991 ( 
.A(n_6488),
.Y(n_6991)
);

OR2x2_ASAP7_75t_L g6992 ( 
.A(n_6557),
.B(n_6174),
.Y(n_6992)
);

OR2x2_ASAP7_75t_SL g6993 ( 
.A(n_6647),
.B(n_6724),
.Y(n_6993)
);

OR2x2_ASAP7_75t_L g6994 ( 
.A(n_6457),
.B(n_6396),
.Y(n_6994)
);

OR2x2_ASAP7_75t_L g6995 ( 
.A(n_6668),
.B(n_6396),
.Y(n_6995)
);

INVx1_ASAP7_75t_L g6996 ( 
.A(n_6452),
.Y(n_6996)
);

INVx1_ASAP7_75t_L g6997 ( 
.A(n_6453),
.Y(n_6997)
);

AOI22xp33_ASAP7_75t_L g6998 ( 
.A1(n_6528),
.A2(n_6231),
.B1(n_6189),
.B2(n_6110),
.Y(n_6998)
);

AND2x2_ASAP7_75t_L g6999 ( 
.A(n_6478),
.B(n_6099),
.Y(n_6999)
);

AND2x4_ASAP7_75t_L g7000 ( 
.A(n_6488),
.B(n_6266),
.Y(n_7000)
);

INVx6_ASAP7_75t_L g7001 ( 
.A(n_6652),
.Y(n_7001)
);

INVx1_ASAP7_75t_L g7002 ( 
.A(n_6456),
.Y(n_7002)
);

AND2x2_ASAP7_75t_L g7003 ( 
.A(n_6506),
.B(n_6099),
.Y(n_7003)
);

AND2x4_ASAP7_75t_L g7004 ( 
.A(n_6488),
.B(n_6266),
.Y(n_7004)
);

INVx2_ASAP7_75t_L g7005 ( 
.A(n_6498),
.Y(n_7005)
);

NAND2xp5_ASAP7_75t_L g7006 ( 
.A(n_6703),
.B(n_6277),
.Y(n_7006)
);

AND2x2_ASAP7_75t_L g7007 ( 
.A(n_6518),
.B(n_6099),
.Y(n_7007)
);

AND2x2_ASAP7_75t_L g7008 ( 
.A(n_6518),
.B(n_6099),
.Y(n_7008)
);

NAND2xp5_ASAP7_75t_L g7009 ( 
.A(n_6703),
.B(n_6278),
.Y(n_7009)
);

INVx2_ASAP7_75t_L g7010 ( 
.A(n_6498),
.Y(n_7010)
);

AOI22xp33_ASAP7_75t_L g7011 ( 
.A1(n_6683),
.A2(n_6231),
.B1(n_6189),
.B2(n_6110),
.Y(n_7011)
);

OR2x2_ASAP7_75t_L g7012 ( 
.A(n_6645),
.B(n_6209),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6458),
.Y(n_7013)
);

INVx2_ASAP7_75t_L g7014 ( 
.A(n_6498),
.Y(n_7014)
);

NAND2xp5_ASAP7_75t_L g7015 ( 
.A(n_6720),
.B(n_6278),
.Y(n_7015)
);

NAND2xp5_ASAP7_75t_L g7016 ( 
.A(n_6720),
.B(n_6155),
.Y(n_7016)
);

NAND2xp5_ASAP7_75t_SL g7017 ( 
.A(n_6657),
.B(n_6219),
.Y(n_7017)
);

NOR2xp33_ASAP7_75t_L g7018 ( 
.A(n_6722),
.B(n_5654),
.Y(n_7018)
);

INVx1_ASAP7_75t_SL g7019 ( 
.A(n_6722),
.Y(n_7019)
);

INVx2_ASAP7_75t_L g7020 ( 
.A(n_6434),
.Y(n_7020)
);

INVx2_ASAP7_75t_L g7021 ( 
.A(n_6434),
.Y(n_7021)
);

INVx2_ASAP7_75t_L g7022 ( 
.A(n_6476),
.Y(n_7022)
);

OR2x6_ASAP7_75t_L g7023 ( 
.A(n_6743),
.B(n_6300),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6460),
.Y(n_7024)
);

BUFx2_ASAP7_75t_L g7025 ( 
.A(n_6697),
.Y(n_7025)
);

NAND3xp33_ASAP7_75t_L g7026 ( 
.A(n_6559),
.B(n_5868),
.C(n_5874),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6464),
.Y(n_7027)
);

NAND2xp5_ASAP7_75t_L g7028 ( 
.A(n_6747),
.B(n_6393),
.Y(n_7028)
);

AND2x2_ASAP7_75t_L g7029 ( 
.A(n_6517),
.B(n_6384),
.Y(n_7029)
);

AND2x2_ASAP7_75t_L g7030 ( 
.A(n_6517),
.B(n_6384),
.Y(n_7030)
);

AOI22xp33_ASAP7_75t_L g7031 ( 
.A1(n_6683),
.A2(n_6231),
.B1(n_6189),
.B2(n_6110),
.Y(n_7031)
);

AND2x2_ASAP7_75t_L g7032 ( 
.A(n_6495),
.B(n_6301),
.Y(n_7032)
);

INVx2_ASAP7_75t_L g7033 ( 
.A(n_6476),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_6495),
.B(n_6301),
.Y(n_7034)
);

NAND2xp5_ASAP7_75t_L g7035 ( 
.A(n_6747),
.B(n_6393),
.Y(n_7035)
);

INVx2_ASAP7_75t_L g7036 ( 
.A(n_6476),
.Y(n_7036)
);

INVxp67_ASAP7_75t_L g7037 ( 
.A(n_6743),
.Y(n_7037)
);

INVx1_ASAP7_75t_L g7038 ( 
.A(n_6467),
.Y(n_7038)
);

INVx2_ASAP7_75t_L g7039 ( 
.A(n_6486),
.Y(n_7039)
);

AND2x2_ASAP7_75t_L g7040 ( 
.A(n_6739),
.B(n_6310),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6475),
.Y(n_7041)
);

INVxp67_ASAP7_75t_SL g7042 ( 
.A(n_6671),
.Y(n_7042)
);

INVx1_ASAP7_75t_L g7043 ( 
.A(n_6485),
.Y(n_7043)
);

AND2x2_ASAP7_75t_L g7044 ( 
.A(n_6739),
.B(n_6310),
.Y(n_7044)
);

AND2x2_ASAP7_75t_L g7045 ( 
.A(n_6555),
.B(n_6315),
.Y(n_7045)
);

OR2x2_ASAP7_75t_L g7046 ( 
.A(n_6620),
.B(n_6209),
.Y(n_7046)
);

NAND2xp5_ASAP7_75t_L g7047 ( 
.A(n_6751),
.B(n_6397),
.Y(n_7047)
);

INVx2_ASAP7_75t_L g7048 ( 
.A(n_6486),
.Y(n_7048)
);

INVx2_ASAP7_75t_L g7049 ( 
.A(n_6486),
.Y(n_7049)
);

OR2x2_ASAP7_75t_L g7050 ( 
.A(n_6410),
.B(n_6349),
.Y(n_7050)
);

NAND2xp33_ASAP7_75t_R g7051 ( 
.A(n_6568),
.B(n_6266),
.Y(n_7051)
);

INVx1_ASAP7_75t_SL g7052 ( 
.A(n_6414),
.Y(n_7052)
);

AND2x2_ASAP7_75t_L g7053 ( 
.A(n_6555),
.B(n_6315),
.Y(n_7053)
);

INVx1_ASAP7_75t_L g7054 ( 
.A(n_6494),
.Y(n_7054)
);

AOI221x1_ASAP7_75t_L g7055 ( 
.A1(n_6487),
.A2(n_6300),
.B1(n_6242),
.B2(n_6243),
.C(n_6236),
.Y(n_7055)
);

AND2x2_ASAP7_75t_L g7056 ( 
.A(n_6569),
.B(n_6146),
.Y(n_7056)
);

BUFx3_ASAP7_75t_L g7057 ( 
.A(n_6755),
.Y(n_7057)
);

NAND2x1_ASAP7_75t_L g7058 ( 
.A(n_6487),
.B(n_6266),
.Y(n_7058)
);

AND2x4_ASAP7_75t_L g7059 ( 
.A(n_6402),
.B(n_6210),
.Y(n_7059)
);

INVx2_ASAP7_75t_L g7060 ( 
.A(n_6487),
.Y(n_7060)
);

INVx1_ASAP7_75t_L g7061 ( 
.A(n_6503),
.Y(n_7061)
);

AND2x4_ASAP7_75t_L g7062 ( 
.A(n_6402),
.B(n_6210),
.Y(n_7062)
);

INVx2_ASAP7_75t_L g7063 ( 
.A(n_6755),
.Y(n_7063)
);

INVx2_ASAP7_75t_L g7064 ( 
.A(n_6758),
.Y(n_7064)
);

INVx2_ASAP7_75t_L g7065 ( 
.A(n_6758),
.Y(n_7065)
);

OR2x2_ASAP7_75t_L g7066 ( 
.A(n_6421),
.B(n_6264),
.Y(n_7066)
);

HB1xp67_ASAP7_75t_L g7067 ( 
.A(n_6751),
.Y(n_7067)
);

AND2x2_ASAP7_75t_L g7068 ( 
.A(n_6569),
.B(n_6146),
.Y(n_7068)
);

INVx2_ASAP7_75t_L g7069 ( 
.A(n_6409),
.Y(n_7069)
);

BUFx3_ASAP7_75t_L g7070 ( 
.A(n_6743),
.Y(n_7070)
);

HB1xp67_ASAP7_75t_L g7071 ( 
.A(n_6756),
.Y(n_7071)
);

INVx2_ASAP7_75t_L g7072 ( 
.A(n_6409),
.Y(n_7072)
);

INVx1_ASAP7_75t_L g7073 ( 
.A(n_6504),
.Y(n_7073)
);

AOI22xp33_ASAP7_75t_L g7074 ( 
.A1(n_6597),
.A2(n_6356),
.B1(n_6363),
.B2(n_6056),
.Y(n_7074)
);

BUFx2_ASAP7_75t_L g7075 ( 
.A(n_6697),
.Y(n_7075)
);

INVx1_ASAP7_75t_L g7076 ( 
.A(n_6508),
.Y(n_7076)
);

INVx2_ASAP7_75t_L g7077 ( 
.A(n_6726),
.Y(n_7077)
);

HB1xp67_ASAP7_75t_L g7078 ( 
.A(n_6756),
.Y(n_7078)
);

OR2x2_ASAP7_75t_L g7079 ( 
.A(n_6428),
.B(n_6108),
.Y(n_7079)
);

AND2x4_ASAP7_75t_L g7080 ( 
.A(n_6402),
.B(n_6210),
.Y(n_7080)
);

INVx1_ASAP7_75t_L g7081 ( 
.A(n_6510),
.Y(n_7081)
);

INVx2_ASAP7_75t_L g7082 ( 
.A(n_6726),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_6735),
.Y(n_7083)
);

NAND2xp5_ASAP7_75t_L g7084 ( 
.A(n_6656),
.B(n_6397),
.Y(n_7084)
);

INVx1_ASAP7_75t_L g7085 ( 
.A(n_6512),
.Y(n_7085)
);

INVx1_ASAP7_75t_L g7086 ( 
.A(n_6513),
.Y(n_7086)
);

NAND2xp5_ASAP7_75t_L g7087 ( 
.A(n_6656),
.B(n_6082),
.Y(n_7087)
);

NOR3xp33_ASAP7_75t_L g7088 ( 
.A(n_6843),
.B(n_6579),
.C(n_6497),
.Y(n_7088)
);

AND2x4_ASAP7_75t_L g7089 ( 
.A(n_6901),
.B(n_6652),
.Y(n_7089)
);

NAND2xp5_ASAP7_75t_L g7090 ( 
.A(n_6843),
.B(n_6399),
.Y(n_7090)
);

INVx1_ASAP7_75t_L g7091 ( 
.A(n_6911),
.Y(n_7091)
);

INVx1_ASAP7_75t_L g7092 ( 
.A(n_6913),
.Y(n_7092)
);

INVx2_ASAP7_75t_SL g7093 ( 
.A(n_6901),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6804),
.B(n_6598),
.Y(n_7094)
);

NOR2x1_ASAP7_75t_L g7095 ( 
.A(n_6837),
.B(n_6735),
.Y(n_7095)
);

AND2x2_ASAP7_75t_L g7096 ( 
.A(n_6818),
.B(n_6561),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_6948),
.Y(n_7097)
);

INVx1_ASAP7_75t_L g7098 ( 
.A(n_6956),
.Y(n_7098)
);

AND2x2_ASAP7_75t_L g7099 ( 
.A(n_6818),
.B(n_6734),
.Y(n_7099)
);

INVx1_ASAP7_75t_L g7100 ( 
.A(n_6958),
.Y(n_7100)
);

AND2x2_ASAP7_75t_L g7101 ( 
.A(n_6821),
.B(n_6593),
.Y(n_7101)
);

INVxp33_ASAP7_75t_L g7102 ( 
.A(n_6809),
.Y(n_7102)
);

NAND2xp5_ASAP7_75t_L g7103 ( 
.A(n_6848),
.B(n_6400),
.Y(n_7103)
);

BUFx3_ASAP7_75t_L g7104 ( 
.A(n_6771),
.Y(n_7104)
);

INVx1_ASAP7_75t_SL g7105 ( 
.A(n_6820),
.Y(n_7105)
);

AND2x2_ASAP7_75t_L g7106 ( 
.A(n_6821),
.B(n_6822),
.Y(n_7106)
);

OAI22xp33_ASAP7_75t_L g7107 ( 
.A1(n_7051),
.A2(n_6719),
.B1(n_6671),
.B2(n_6762),
.Y(n_7107)
);

INVx1_ASAP7_75t_L g7108 ( 
.A(n_6985),
.Y(n_7108)
);

INVx2_ASAP7_75t_L g7109 ( 
.A(n_6901),
.Y(n_7109)
);

OR2x2_ASAP7_75t_L g7110 ( 
.A(n_6773),
.B(n_6530),
.Y(n_7110)
);

AND2x2_ASAP7_75t_L g7111 ( 
.A(n_6822),
.B(n_6401),
.Y(n_7111)
);

NAND2xp5_ASAP7_75t_L g7112 ( 
.A(n_6872),
.B(n_6419),
.Y(n_7112)
);

AND2x2_ASAP7_75t_L g7113 ( 
.A(n_6829),
.B(n_6604),
.Y(n_7113)
);

INVx1_ASAP7_75t_L g7114 ( 
.A(n_6807),
.Y(n_7114)
);

INVx2_ASAP7_75t_L g7115 ( 
.A(n_6971),
.Y(n_7115)
);

NAND2xp5_ASAP7_75t_L g7116 ( 
.A(n_6983),
.B(n_6661),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_6983),
.B(n_6661),
.Y(n_7117)
);

INVx2_ASAP7_75t_L g7118 ( 
.A(n_6971),
.Y(n_7118)
);

CKINVDCx14_ASAP7_75t_R g7119 ( 
.A(n_6829),
.Y(n_7119)
);

INVxp67_ASAP7_75t_L g7120 ( 
.A(n_6792),
.Y(n_7120)
);

INVx2_ASAP7_75t_L g7121 ( 
.A(n_6971),
.Y(n_7121)
);

AND2x2_ASAP7_75t_L g7122 ( 
.A(n_6832),
.B(n_6573),
.Y(n_7122)
);

AND2x2_ASAP7_75t_L g7123 ( 
.A(n_6832),
.B(n_6573),
.Y(n_7123)
);

NAND2x1p5_ASAP7_75t_L g7124 ( 
.A(n_6802),
.B(n_6652),
.Y(n_7124)
);

INVx2_ASAP7_75t_L g7125 ( 
.A(n_6837),
.Y(n_7125)
);

AND2x2_ASAP7_75t_L g7126 ( 
.A(n_6813),
.B(n_6587),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6813),
.B(n_6587),
.Y(n_7127)
);

INVx1_ASAP7_75t_L g7128 ( 
.A(n_7067),
.Y(n_7128)
);

OR2x2_ASAP7_75t_L g7129 ( 
.A(n_7052),
.B(n_6493),
.Y(n_7129)
);

AND2x4_ASAP7_75t_L g7130 ( 
.A(n_6771),
.B(n_6652),
.Y(n_7130)
);

AND2x2_ASAP7_75t_L g7131 ( 
.A(n_6840),
.B(n_6704),
.Y(n_7131)
);

OR2x2_ASAP7_75t_L g7132 ( 
.A(n_6838),
.B(n_6632),
.Y(n_7132)
);

NAND2xp5_ASAP7_75t_L g7133 ( 
.A(n_6984),
.B(n_6622),
.Y(n_7133)
);

OR2x6_ASAP7_75t_L g7134 ( 
.A(n_6850),
.B(n_6743),
.Y(n_7134)
);

INVx1_ASAP7_75t_L g7135 ( 
.A(n_7071),
.Y(n_7135)
);

INVx1_ASAP7_75t_L g7136 ( 
.A(n_7078),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6984),
.Y(n_7137)
);

INVx1_ASAP7_75t_L g7138 ( 
.A(n_6986),
.Y(n_7138)
);

INVx2_ASAP7_75t_L g7139 ( 
.A(n_6837),
.Y(n_7139)
);

NAND2x1_ASAP7_75t_L g7140 ( 
.A(n_6859),
.B(n_6719),
.Y(n_7140)
);

INVx1_ASAP7_75t_L g7141 ( 
.A(n_6986),
.Y(n_7141)
);

BUFx2_ASAP7_75t_L g7142 ( 
.A(n_6771),
.Y(n_7142)
);

BUFx2_ASAP7_75t_L g7143 ( 
.A(n_6850),
.Y(n_7143)
);

NAND2xp5_ASAP7_75t_L g7144 ( 
.A(n_6966),
.B(n_6622),
.Y(n_7144)
);

AND2x2_ASAP7_75t_L g7145 ( 
.A(n_6840),
.B(n_6687),
.Y(n_7145)
);

AND2x2_ASAP7_75t_L g7146 ( 
.A(n_6841),
.B(n_6687),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6856),
.Y(n_7147)
);

AND2x2_ASAP7_75t_L g7148 ( 
.A(n_6841),
.B(n_6708),
.Y(n_7148)
);

AND2x2_ASAP7_75t_L g7149 ( 
.A(n_6844),
.B(n_6708),
.Y(n_7149)
);

AND2x4_ASAP7_75t_L g7150 ( 
.A(n_6803),
.B(n_6507),
.Y(n_7150)
);

AND2x4_ASAP7_75t_L g7151 ( 
.A(n_6803),
.B(n_6507),
.Y(n_7151)
);

OR2x2_ASAP7_75t_L g7152 ( 
.A(n_6955),
.B(n_6994),
.Y(n_7152)
);

NAND2xp5_ASAP7_75t_L g7153 ( 
.A(n_6966),
.B(n_6860),
.Y(n_7153)
);

INVxp67_ASAP7_75t_SL g7154 ( 
.A(n_6922),
.Y(n_7154)
);

OR2x2_ASAP7_75t_L g7155 ( 
.A(n_7077),
.B(n_6558),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6856),
.Y(n_7156)
);

INVxp67_ASAP7_75t_L g7157 ( 
.A(n_6817),
.Y(n_7157)
);

OR2x2_ASAP7_75t_L g7158 ( 
.A(n_7077),
.B(n_6712),
.Y(n_7158)
);

NAND2xp5_ASAP7_75t_L g7159 ( 
.A(n_6860),
.B(n_6625),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_6868),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_6998),
.B(n_6625),
.Y(n_7161)
);

NAND2xp5_ASAP7_75t_L g7162 ( 
.A(n_6998),
.B(n_6626),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_SL g7163 ( 
.A(n_6951),
.B(n_6667),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_L g7164 ( 
.A(n_6863),
.B(n_6626),
.Y(n_7164)
);

NAND2xp5_ASAP7_75t_L g7165 ( 
.A(n_6870),
.B(n_6627),
.Y(n_7165)
);

AND2x2_ASAP7_75t_L g7166 ( 
.A(n_6844),
.B(n_6686),
.Y(n_7166)
);

AND2x2_ASAP7_75t_L g7167 ( 
.A(n_6781),
.B(n_6686),
.Y(n_7167)
);

INVx1_ASAP7_75t_L g7168 ( 
.A(n_6926),
.Y(n_7168)
);

AND2x4_ASAP7_75t_L g7169 ( 
.A(n_6803),
.B(n_6616),
.Y(n_7169)
);

AND2x2_ASAP7_75t_L g7170 ( 
.A(n_6781),
.B(n_6442),
.Y(n_7170)
);

AND2x2_ASAP7_75t_L g7171 ( 
.A(n_6796),
.B(n_6730),
.Y(n_7171)
);

AND2x2_ASAP7_75t_L g7172 ( 
.A(n_6796),
.B(n_7003),
.Y(n_7172)
);

HB1xp67_ASAP7_75t_L g7173 ( 
.A(n_6922),
.Y(n_7173)
);

OA21x2_ASAP7_75t_L g7174 ( 
.A1(n_7055),
.A2(n_7031),
.B(n_7011),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_6929),
.Y(n_7175)
);

OR2x2_ASAP7_75t_L g7176 ( 
.A(n_7082),
.B(n_6712),
.Y(n_7176)
);

INVx1_ASAP7_75t_L g7177 ( 
.A(n_6937),
.Y(n_7177)
);

INVx1_ASAP7_75t_L g7178 ( 
.A(n_6944),
.Y(n_7178)
);

AND2x4_ASAP7_75t_L g7179 ( 
.A(n_6780),
.B(n_6616),
.Y(n_7179)
);

INVx1_ASAP7_75t_L g7180 ( 
.A(n_6982),
.Y(n_7180)
);

AND2x4_ASAP7_75t_SL g7181 ( 
.A(n_6780),
.B(n_6790),
.Y(n_7181)
);

INVx2_ASAP7_75t_L g7182 ( 
.A(n_6868),
.Y(n_7182)
);

AND2x4_ASAP7_75t_L g7183 ( 
.A(n_6780),
.B(n_6627),
.Y(n_7183)
);

INVx2_ASAP7_75t_L g7184 ( 
.A(n_6868),
.Y(n_7184)
);

AND2x4_ASAP7_75t_L g7185 ( 
.A(n_6790),
.B(n_6631),
.Y(n_7185)
);

NOR2xp33_ASAP7_75t_L g7186 ( 
.A(n_6812),
.B(n_6699),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_6982),
.Y(n_7187)
);

INVx2_ASAP7_75t_L g7188 ( 
.A(n_6785),
.Y(n_7188)
);

AND2x2_ASAP7_75t_L g7189 ( 
.A(n_7003),
.B(n_6730),
.Y(n_7189)
);

INVxp67_ASAP7_75t_SL g7190 ( 
.A(n_6924),
.Y(n_7190)
);

OR2x2_ASAP7_75t_L g7191 ( 
.A(n_7082),
.B(n_6660),
.Y(n_7191)
);

OR2x2_ASAP7_75t_L g7192 ( 
.A(n_7083),
.B(n_6538),
.Y(n_7192)
);

AND2x2_ASAP7_75t_L g7193 ( 
.A(n_6972),
.B(n_6532),
.Y(n_7193)
);

NAND2xp5_ASAP7_75t_L g7194 ( 
.A(n_6871),
.B(n_6631),
.Y(n_7194)
);

INVxp67_ASAP7_75t_SL g7195 ( 
.A(n_6924),
.Y(n_7195)
);

BUFx2_ASAP7_75t_SL g7196 ( 
.A(n_6790),
.Y(n_7196)
);

OR2x2_ASAP7_75t_L g7197 ( 
.A(n_7083),
.B(n_6551),
.Y(n_7197)
);

AND2x4_ASAP7_75t_L g7198 ( 
.A(n_6855),
.B(n_6524),
.Y(n_7198)
);

AND2x2_ASAP7_75t_L g7199 ( 
.A(n_6972),
.B(n_6532),
.Y(n_7199)
);

INVx1_ASAP7_75t_L g7200 ( 
.A(n_6874),
.Y(n_7200)
);

AND2x2_ASAP7_75t_L g7201 ( 
.A(n_6976),
.B(n_6534),
.Y(n_7201)
);

AND2x2_ASAP7_75t_L g7202 ( 
.A(n_6976),
.B(n_6534),
.Y(n_7202)
);

AND2x2_ASAP7_75t_L g7203 ( 
.A(n_6797),
.B(n_6691),
.Y(n_7203)
);

NOR2xp67_ASAP7_75t_L g7204 ( 
.A(n_6859),
.B(n_6489),
.Y(n_7204)
);

OR2x2_ASAP7_75t_L g7205 ( 
.A(n_6995),
.B(n_6748),
.Y(n_7205)
);

AND2x4_ASAP7_75t_L g7206 ( 
.A(n_6855),
.B(n_6524),
.Y(n_7206)
);

INVx2_ASAP7_75t_L g7207 ( 
.A(n_6785),
.Y(n_7207)
);

NAND2xp5_ASAP7_75t_L g7208 ( 
.A(n_6795),
.B(n_6524),
.Y(n_7208)
);

OR2x6_ASAP7_75t_L g7209 ( 
.A(n_6857),
.B(n_6719),
.Y(n_7209)
);

AND2x2_ASAP7_75t_L g7210 ( 
.A(n_6797),
.B(n_6691),
.Y(n_7210)
);

AND2x2_ASAP7_75t_L g7211 ( 
.A(n_6800),
.B(n_6719),
.Y(n_7211)
);

AND2x2_ASAP7_75t_L g7212 ( 
.A(n_6800),
.B(n_6541),
.Y(n_7212)
);

AND2x2_ASAP7_75t_L g7213 ( 
.A(n_6894),
.B(n_6541),
.Y(n_7213)
);

INVx2_ASAP7_75t_L g7214 ( 
.A(n_6785),
.Y(n_7214)
);

NOR2xp67_ASAP7_75t_L g7215 ( 
.A(n_6859),
.B(n_6489),
.Y(n_7215)
);

AND2x2_ASAP7_75t_L g7216 ( 
.A(n_6894),
.B(n_6533),
.Y(n_7216)
);

AND2x2_ASAP7_75t_L g7217 ( 
.A(n_7056),
.B(n_7068),
.Y(n_7217)
);

INVxp67_ASAP7_75t_L g7218 ( 
.A(n_7025),
.Y(n_7218)
);

INVx2_ASAP7_75t_L g7219 ( 
.A(n_6785),
.Y(n_7219)
);

INVx2_ASAP7_75t_L g7220 ( 
.A(n_6794),
.Y(n_7220)
);

NAND3xp33_ASAP7_75t_L g7221 ( 
.A(n_7074),
.B(n_7051),
.C(n_7026),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_6899),
.Y(n_7222)
);

HB1xp67_ASAP7_75t_L g7223 ( 
.A(n_6933),
.Y(n_7223)
);

AND2x2_ASAP7_75t_L g7224 ( 
.A(n_7056),
.B(n_6713),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_6900),
.Y(n_7225)
);

NAND2xp5_ASAP7_75t_L g7226 ( 
.A(n_6774),
.B(n_6502),
.Y(n_7226)
);

AND2x2_ASAP7_75t_L g7227 ( 
.A(n_7068),
.B(n_6713),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_6902),
.Y(n_7228)
);

AND2x2_ASAP7_75t_L g7229 ( 
.A(n_7007),
.B(n_7008),
.Y(n_7229)
);

INVx1_ASAP7_75t_L g7230 ( 
.A(n_6906),
.Y(n_7230)
);

NAND2xp5_ASAP7_75t_L g7231 ( 
.A(n_6775),
.B(n_6502),
.Y(n_7231)
);

NAND2xp5_ASAP7_75t_L g7232 ( 
.A(n_6830),
.B(n_6515),
.Y(n_7232)
);

AND2x2_ASAP7_75t_L g7233 ( 
.A(n_7007),
.B(n_6548),
.Y(n_7233)
);

INVx3_ASAP7_75t_L g7234 ( 
.A(n_6928),
.Y(n_7234)
);

AND2x4_ASAP7_75t_L g7235 ( 
.A(n_6855),
.B(n_6670),
.Y(n_7235)
);

NAND2xp5_ASAP7_75t_L g7236 ( 
.A(n_6833),
.B(n_6515),
.Y(n_7236)
);

AND2x2_ASAP7_75t_L g7237 ( 
.A(n_7008),
.B(n_6548),
.Y(n_7237)
);

AND2x2_ASAP7_75t_L g7238 ( 
.A(n_6999),
.B(n_6589),
.Y(n_7238)
);

INVx1_ASAP7_75t_SL g7239 ( 
.A(n_6857),
.Y(n_7239)
);

OR2x2_ASAP7_75t_L g7240 ( 
.A(n_6993),
.B(n_6585),
.Y(n_7240)
);

AND2x2_ASAP7_75t_SL g7241 ( 
.A(n_7075),
.B(n_6663),
.Y(n_7241)
);

NAND2xp5_ASAP7_75t_L g7242 ( 
.A(n_6853),
.B(n_6537),
.Y(n_7242)
);

HB1xp67_ASAP7_75t_L g7243 ( 
.A(n_6933),
.Y(n_7243)
);

AND2x2_ASAP7_75t_L g7244 ( 
.A(n_6999),
.B(n_6589),
.Y(n_7244)
);

AND2x2_ASAP7_75t_L g7245 ( 
.A(n_6968),
.B(n_6970),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6919),
.Y(n_7246)
);

NAND2xp5_ASAP7_75t_L g7247 ( 
.A(n_6921),
.B(n_6537),
.Y(n_7247)
);

INVx4_ASAP7_75t_L g7248 ( 
.A(n_6787),
.Y(n_7248)
);

AND2x4_ASAP7_75t_L g7249 ( 
.A(n_7070),
.B(n_6670),
.Y(n_7249)
);

AND2x2_ASAP7_75t_L g7250 ( 
.A(n_6968),
.B(n_6674),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_L g7251 ( 
.A(n_6923),
.B(n_6927),
.Y(n_7251)
);

INVx1_ASAP7_75t_L g7252 ( 
.A(n_6932),
.Y(n_7252)
);

OR2x2_ASAP7_75t_L g7253 ( 
.A(n_6782),
.B(n_6407),
.Y(n_7253)
);

OAI22xp5_ASAP7_75t_L g7254 ( 
.A1(n_7074),
.A2(n_6641),
.B1(n_6413),
.B2(n_6415),
.Y(n_7254)
);

INVx2_ASAP7_75t_SL g7255 ( 
.A(n_6846),
.Y(n_7255)
);

AND2x2_ASAP7_75t_L g7256 ( 
.A(n_6970),
.B(n_6674),
.Y(n_7256)
);

INVx1_ASAP7_75t_L g7257 ( 
.A(n_6876),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_6876),
.Y(n_7258)
);

AND2x4_ASAP7_75t_L g7259 ( 
.A(n_7070),
.B(n_6670),
.Y(n_7259)
);

AND2x2_ASAP7_75t_L g7260 ( 
.A(n_6961),
.B(n_6962),
.Y(n_7260)
);

HB1xp67_ASAP7_75t_L g7261 ( 
.A(n_6974),
.Y(n_7261)
);

AND2x2_ASAP7_75t_L g7262 ( 
.A(n_6961),
.B(n_6675),
.Y(n_7262)
);

INVx2_ASAP7_75t_L g7263 ( 
.A(n_6794),
.Y(n_7263)
);

AND2x2_ASAP7_75t_L g7264 ( 
.A(n_6962),
.B(n_6873),
.Y(n_7264)
);

OR2x2_ASAP7_75t_L g7265 ( 
.A(n_6867),
.B(n_6407),
.Y(n_7265)
);

OR2x2_ASAP7_75t_L g7266 ( 
.A(n_6973),
.B(n_6977),
.Y(n_7266)
);

AND2x4_ASAP7_75t_L g7267 ( 
.A(n_6991),
.B(n_6572),
.Y(n_7267)
);

BUFx2_ASAP7_75t_L g7268 ( 
.A(n_6866),
.Y(n_7268)
);

AND2x2_ASAP7_75t_L g7269 ( 
.A(n_6941),
.B(n_6675),
.Y(n_7269)
);

AND2x2_ASAP7_75t_L g7270 ( 
.A(n_6809),
.B(n_6918),
.Y(n_7270)
);

AOI22xp5_ASAP7_75t_L g7271 ( 
.A1(n_6875),
.A2(n_6644),
.B1(n_6468),
.B2(n_6690),
.Y(n_7271)
);

AND2x2_ASAP7_75t_L g7272 ( 
.A(n_6918),
.B(n_6468),
.Y(n_7272)
);

NAND2xp5_ASAP7_75t_L g7273 ( 
.A(n_6828),
.B(n_6854),
.Y(n_7273)
);

AND2x2_ASAP7_75t_L g7274 ( 
.A(n_6915),
.B(n_6711),
.Y(n_7274)
);

AND2x2_ASAP7_75t_L g7275 ( 
.A(n_6915),
.B(n_6711),
.Y(n_7275)
);

NAND2xp5_ASAP7_75t_L g7276 ( 
.A(n_6858),
.B(n_6540),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_6878),
.Y(n_7277)
);

AND2x2_ASAP7_75t_L g7278 ( 
.A(n_6916),
.B(n_6709),
.Y(n_7278)
);

INVx2_ASAP7_75t_SL g7279 ( 
.A(n_6935),
.Y(n_7279)
);

INVx2_ASAP7_75t_L g7280 ( 
.A(n_6794),
.Y(n_7280)
);

AND2x4_ASAP7_75t_L g7281 ( 
.A(n_6991),
.B(n_6572),
.Y(n_7281)
);

INVx2_ASAP7_75t_L g7282 ( 
.A(n_6974),
.Y(n_7282)
);

INVxp67_ASAP7_75t_L g7283 ( 
.A(n_6940),
.Y(n_7283)
);

AND2x2_ASAP7_75t_L g7284 ( 
.A(n_6916),
.B(n_6709),
.Y(n_7284)
);

NAND2xp5_ASAP7_75t_L g7285 ( 
.A(n_6880),
.B(n_6540),
.Y(n_7285)
);

NAND3xp33_ASAP7_75t_L g7286 ( 
.A(n_6875),
.B(n_6415),
.C(n_6413),
.Y(n_7286)
);

INVx1_ASAP7_75t_L g7287 ( 
.A(n_6878),
.Y(n_7287)
);

AND2x2_ASAP7_75t_L g7288 ( 
.A(n_6936),
.B(n_6729),
.Y(n_7288)
);

INVx1_ASAP7_75t_L g7289 ( 
.A(n_6904),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_L g7290 ( 
.A(n_6883),
.B(n_6544),
.Y(n_7290)
);

HB1xp67_ASAP7_75t_L g7291 ( 
.A(n_6814),
.Y(n_7291)
);

AND2x4_ASAP7_75t_L g7292 ( 
.A(n_7005),
.B(n_6581),
.Y(n_7292)
);

AND2x2_ASAP7_75t_L g7293 ( 
.A(n_6936),
.B(n_6729),
.Y(n_7293)
);

INVx2_ASAP7_75t_L g7294 ( 
.A(n_6799),
.Y(n_7294)
);

INVx1_ASAP7_75t_L g7295 ( 
.A(n_6904),
.Y(n_7295)
);

INVx2_ASAP7_75t_L g7296 ( 
.A(n_6799),
.Y(n_7296)
);

OAI21xp5_ASAP7_75t_SL g7297 ( 
.A1(n_7017),
.A2(n_6690),
.B(n_6717),
.Y(n_7297)
);

NAND2xp5_ASAP7_75t_L g7298 ( 
.A(n_6798),
.B(n_6544),
.Y(n_7298)
);

AND2x2_ASAP7_75t_L g7299 ( 
.A(n_7018),
.B(n_6594),
.Y(n_7299)
);

NOR2xp67_ASAP7_75t_L g7300 ( 
.A(n_6799),
.B(n_6556),
.Y(n_7300)
);

OR2x2_ASAP7_75t_L g7301 ( 
.A(n_6973),
.B(n_6422),
.Y(n_7301)
);

OAI22xp5_ASAP7_75t_L g7302 ( 
.A1(n_7011),
.A2(n_7031),
.B1(n_6939),
.B2(n_7017),
.Y(n_7302)
);

NOR2xp33_ASAP7_75t_L g7303 ( 
.A(n_6787),
.B(n_5590),
.Y(n_7303)
);

INVx3_ASAP7_75t_L g7304 ( 
.A(n_6935),
.Y(n_7304)
);

INVx2_ASAP7_75t_L g7305 ( 
.A(n_6823),
.Y(n_7305)
);

AND2x2_ASAP7_75t_L g7306 ( 
.A(n_7018),
.B(n_6594),
.Y(n_7306)
);

NAND2xp5_ASAP7_75t_L g7307 ( 
.A(n_6805),
.B(n_6556),
.Y(n_7307)
);

INVx1_ASAP7_75t_L g7308 ( 
.A(n_6907),
.Y(n_7308)
);

AND2x2_ASAP7_75t_L g7309 ( 
.A(n_6947),
.B(n_6717),
.Y(n_7309)
);

INVx2_ASAP7_75t_L g7310 ( 
.A(n_6823),
.Y(n_7310)
);

AND2x4_ASAP7_75t_L g7311 ( 
.A(n_7005),
.B(n_6581),
.Y(n_7311)
);

INVx1_ASAP7_75t_L g7312 ( 
.A(n_6907),
.Y(n_7312)
);

INVx1_ASAP7_75t_L g7313 ( 
.A(n_6908),
.Y(n_7313)
);

AND2x2_ASAP7_75t_L g7314 ( 
.A(n_6947),
.B(n_6746),
.Y(n_7314)
);

OAI22xp5_ASAP7_75t_L g7315 ( 
.A1(n_7042),
.A2(n_6056),
.B1(n_5859),
.B2(n_5840),
.Y(n_7315)
);

INVx1_ASAP7_75t_L g7316 ( 
.A(n_6908),
.Y(n_7316)
);

AND2x2_ASAP7_75t_L g7317 ( 
.A(n_6945),
.B(n_6746),
.Y(n_7317)
);

OR2x2_ASAP7_75t_L g7318 ( 
.A(n_6977),
.B(n_6978),
.Y(n_7318)
);

AND2x4_ASAP7_75t_L g7319 ( 
.A(n_7010),
.B(n_7014),
.Y(n_7319)
);

INVx2_ASAP7_75t_L g7320 ( 
.A(n_6823),
.Y(n_7320)
);

HB1xp67_ASAP7_75t_L g7321 ( 
.A(n_6814),
.Y(n_7321)
);

INVx2_ASAP7_75t_L g7322 ( 
.A(n_6931),
.Y(n_7322)
);

NAND2xp5_ASAP7_75t_L g7323 ( 
.A(n_6808),
.B(n_6566),
.Y(n_7323)
);

INVx2_ASAP7_75t_L g7324 ( 
.A(n_6931),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_L g7325 ( 
.A(n_6778),
.B(n_6779),
.Y(n_7325)
);

AND2x2_ASAP7_75t_L g7326 ( 
.A(n_6945),
.B(n_6746),
.Y(n_7326)
);

NOR2xp33_ASAP7_75t_L g7327 ( 
.A(n_6787),
.B(n_5590),
.Y(n_7327)
);

NAND2xp5_ASAP7_75t_L g7328 ( 
.A(n_6783),
.B(n_6566),
.Y(n_7328)
);

AOI22xp33_ASAP7_75t_SL g7329 ( 
.A1(n_6960),
.A2(n_6644),
.B1(n_6630),
.B2(n_6562),
.Y(n_7329)
);

NAND2xp5_ASAP7_75t_L g7330 ( 
.A(n_6784),
.B(n_6570),
.Y(n_7330)
);

NAND2xp5_ASAP7_75t_L g7331 ( 
.A(n_6788),
.B(n_6570),
.Y(n_7331)
);

AND2x2_ASAP7_75t_L g7332 ( 
.A(n_6864),
.B(n_6746),
.Y(n_7332)
);

INVx1_ASAP7_75t_L g7333 ( 
.A(n_6912),
.Y(n_7333)
);

OR2x2_ASAP7_75t_L g7334 ( 
.A(n_6978),
.B(n_6422),
.Y(n_7334)
);

AND2x2_ASAP7_75t_L g7335 ( 
.A(n_6864),
.B(n_6640),
.Y(n_7335)
);

INVx1_ASAP7_75t_L g7336 ( 
.A(n_6912),
.Y(n_7336)
);

INVx1_ASAP7_75t_L g7337 ( 
.A(n_6777),
.Y(n_7337)
);

INVx2_ASAP7_75t_L g7338 ( 
.A(n_6931),
.Y(n_7338)
);

INVx2_ASAP7_75t_L g7339 ( 
.A(n_6931),
.Y(n_7339)
);

INVx1_ASAP7_75t_L g7340 ( 
.A(n_6777),
.Y(n_7340)
);

INVx1_ASAP7_75t_L g7341 ( 
.A(n_6786),
.Y(n_7341)
);

AND2x2_ASAP7_75t_L g7342 ( 
.A(n_6882),
.B(n_6640),
.Y(n_7342)
);

NAND2xp5_ASAP7_75t_L g7343 ( 
.A(n_6826),
.B(n_6757),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_6786),
.Y(n_7344)
);

AND2x2_ASAP7_75t_L g7345 ( 
.A(n_6882),
.B(n_6885),
.Y(n_7345)
);

AND2x2_ASAP7_75t_L g7346 ( 
.A(n_6885),
.B(n_6650),
.Y(n_7346)
);

AND2x2_ASAP7_75t_L g7347 ( 
.A(n_6776),
.B(n_6650),
.Y(n_7347)
);

AND2x2_ASAP7_75t_L g7348 ( 
.A(n_6776),
.B(n_6653),
.Y(n_7348)
);

AND2x2_ASAP7_75t_L g7349 ( 
.A(n_6903),
.B(n_6653),
.Y(n_7349)
);

NAND3xp33_ASAP7_75t_L g7350 ( 
.A(n_6816),
.B(n_6677),
.C(n_6760),
.Y(n_7350)
);

NAND2xp5_ASAP7_75t_L g7351 ( 
.A(n_6826),
.B(n_6757),
.Y(n_7351)
);

HB1xp67_ASAP7_75t_L g7352 ( 
.A(n_6814),
.Y(n_7352)
);

AND2x2_ASAP7_75t_L g7353 ( 
.A(n_6903),
.B(n_6659),
.Y(n_7353)
);

AND2x2_ASAP7_75t_L g7354 ( 
.A(n_6909),
.B(n_6659),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_L g7355 ( 
.A(n_6827),
.B(n_6831),
.Y(n_7355)
);

INVx1_ASAP7_75t_L g7356 ( 
.A(n_6789),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_6827),
.B(n_6757),
.Y(n_7357)
);

INVx1_ASAP7_75t_L g7358 ( 
.A(n_6789),
.Y(n_7358)
);

OR2x2_ASAP7_75t_L g7359 ( 
.A(n_6979),
.B(n_6431),
.Y(n_7359)
);

NOR2xp33_ASAP7_75t_L g7360 ( 
.A(n_7119),
.B(n_6866),
.Y(n_7360)
);

BUFx3_ASAP7_75t_L g7361 ( 
.A(n_7142),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_7173),
.Y(n_7362)
);

AND2x4_ASAP7_75t_L g7363 ( 
.A(n_7235),
.B(n_7010),
.Y(n_7363)
);

NAND2xp5_ASAP7_75t_L g7364 ( 
.A(n_7122),
.B(n_7123),
.Y(n_7364)
);

AND2x2_ASAP7_75t_L g7365 ( 
.A(n_7106),
.B(n_6877),
.Y(n_7365)
);

INVx1_ASAP7_75t_L g7366 ( 
.A(n_7173),
.Y(n_7366)
);

HB1xp67_ASAP7_75t_L g7367 ( 
.A(n_7174),
.Y(n_7367)
);

AND2x2_ASAP7_75t_L g7368 ( 
.A(n_7245),
.B(n_6909),
.Y(n_7368)
);

AOI21xp5_ASAP7_75t_L g7369 ( 
.A1(n_7163),
.A2(n_6960),
.B(n_6934),
.Y(n_7369)
);

HB1xp67_ASAP7_75t_L g7370 ( 
.A(n_7174),
.Y(n_7370)
);

OR2x2_ASAP7_75t_L g7371 ( 
.A(n_7105),
.B(n_7063),
.Y(n_7371)
);

INVx3_ASAP7_75t_L g7372 ( 
.A(n_7235),
.Y(n_7372)
);

AND2x2_ASAP7_75t_L g7373 ( 
.A(n_7255),
.B(n_6877),
.Y(n_7373)
);

AND2x2_ASAP7_75t_L g7374 ( 
.A(n_7217),
.B(n_7229),
.Y(n_7374)
);

AND2x2_ASAP7_75t_L g7375 ( 
.A(n_7193),
.B(n_6879),
.Y(n_7375)
);

AND2x2_ASAP7_75t_L g7376 ( 
.A(n_7199),
.B(n_6879),
.Y(n_7376)
);

AND2x2_ASAP7_75t_L g7377 ( 
.A(n_7201),
.B(n_6910),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_7223),
.Y(n_7378)
);

AND2x2_ASAP7_75t_L g7379 ( 
.A(n_7202),
.B(n_6910),
.Y(n_7379)
);

INVx2_ASAP7_75t_L g7380 ( 
.A(n_7198),
.Y(n_7380)
);

CKINVDCx5p33_ASAP7_75t_R g7381 ( 
.A(n_7196),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_7189),
.B(n_7146),
.Y(n_7382)
);

AND2x2_ASAP7_75t_L g7383 ( 
.A(n_7145),
.B(n_6914),
.Y(n_7383)
);

NAND2xp5_ASAP7_75t_L g7384 ( 
.A(n_7250),
.B(n_6772),
.Y(n_7384)
);

AND2x2_ASAP7_75t_L g7385 ( 
.A(n_7233),
.B(n_7237),
.Y(n_7385)
);

HB1xp67_ASAP7_75t_L g7386 ( 
.A(n_7261),
.Y(n_7386)
);

AND2x2_ASAP7_75t_L g7387 ( 
.A(n_7166),
.B(n_7148),
.Y(n_7387)
);

AND2x2_ASAP7_75t_L g7388 ( 
.A(n_7119),
.B(n_6914),
.Y(n_7388)
);

OR2x2_ASAP7_75t_L g7389 ( 
.A(n_7105),
.B(n_7063),
.Y(n_7389)
);

AND2x2_ASAP7_75t_L g7390 ( 
.A(n_7238),
.B(n_6889),
.Y(n_7390)
);

NOR2xp33_ASAP7_75t_L g7391 ( 
.A(n_7102),
.B(n_7157),
.Y(n_7391)
);

INVxp67_ASAP7_75t_L g7392 ( 
.A(n_7095),
.Y(n_7392)
);

INVx2_ASAP7_75t_L g7393 ( 
.A(n_7198),
.Y(n_7393)
);

AND2x2_ASAP7_75t_L g7394 ( 
.A(n_7244),
.B(n_6831),
.Y(n_7394)
);

AND2x2_ASAP7_75t_L g7395 ( 
.A(n_7213),
.B(n_6834),
.Y(n_7395)
);

AND2x2_ASAP7_75t_L g7396 ( 
.A(n_7256),
.B(n_6834),
.Y(n_7396)
);

AND2x2_ASAP7_75t_L g7397 ( 
.A(n_7149),
.B(n_6835),
.Y(n_7397)
);

NOR2x1_ASAP7_75t_L g7398 ( 
.A(n_7134),
.B(n_7057),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_7223),
.Y(n_7399)
);

AND2x4_ASAP7_75t_SL g7400 ( 
.A(n_7150),
.B(n_6835),
.Y(n_7400)
);

INVx1_ASAP7_75t_L g7401 ( 
.A(n_7243),
.Y(n_7401)
);

NAND2xp5_ASAP7_75t_L g7402 ( 
.A(n_7224),
.B(n_6825),
.Y(n_7402)
);

INVx1_ASAP7_75t_L g7403 ( 
.A(n_7243),
.Y(n_7403)
);

BUFx3_ASAP7_75t_L g7404 ( 
.A(n_7104),
.Y(n_7404)
);

BUFx3_ASAP7_75t_L g7405 ( 
.A(n_7104),
.Y(n_7405)
);

INVx1_ASAP7_75t_L g7406 ( 
.A(n_7154),
.Y(n_7406)
);

AND2x2_ASAP7_75t_L g7407 ( 
.A(n_7227),
.B(n_6889),
.Y(n_7407)
);

NAND2xp5_ASAP7_75t_L g7408 ( 
.A(n_7239),
.B(n_6836),
.Y(n_7408)
);

AND2x2_ASAP7_75t_L g7409 ( 
.A(n_7111),
.B(n_6895),
.Y(n_7409)
);

INVx2_ASAP7_75t_L g7410 ( 
.A(n_7206),
.Y(n_7410)
);

INVx2_ASAP7_75t_L g7411 ( 
.A(n_7206),
.Y(n_7411)
);

OR2x2_ASAP7_75t_L g7412 ( 
.A(n_7144),
.B(n_7064),
.Y(n_7412)
);

NOR2xp33_ASAP7_75t_L g7413 ( 
.A(n_7102),
.B(n_6793),
.Y(n_7413)
);

INVx1_ASAP7_75t_SL g7414 ( 
.A(n_7181),
.Y(n_7414)
);

NOR2x1_ASAP7_75t_L g7415 ( 
.A(n_7134),
.B(n_7107),
.Y(n_7415)
);

AND2x2_ASAP7_75t_L g7416 ( 
.A(n_7126),
.B(n_7127),
.Y(n_7416)
);

AND2x2_ASAP7_75t_SL g7417 ( 
.A(n_7088),
.B(n_6845),
.Y(n_7417)
);

AND2x4_ASAP7_75t_SL g7418 ( 
.A(n_7150),
.B(n_6836),
.Y(n_7418)
);

INVx2_ASAP7_75t_L g7419 ( 
.A(n_7304),
.Y(n_7419)
);

OR2x2_ASAP7_75t_L g7420 ( 
.A(n_7144),
.B(n_7064),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_7154),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_7239),
.B(n_7272),
.Y(n_7422)
);

AND2x2_ASAP7_75t_L g7423 ( 
.A(n_7101),
.B(n_6839),
.Y(n_7423)
);

INVx1_ASAP7_75t_L g7424 ( 
.A(n_7190),
.Y(n_7424)
);

NAND2xp5_ASAP7_75t_L g7425 ( 
.A(n_7345),
.B(n_6839),
.Y(n_7425)
);

INVx1_ASAP7_75t_L g7426 ( 
.A(n_7190),
.Y(n_7426)
);

HB1xp67_ASAP7_75t_L g7427 ( 
.A(n_7261),
.Y(n_7427)
);

AND2x2_ASAP7_75t_L g7428 ( 
.A(n_7172),
.B(n_6895),
.Y(n_7428)
);

NAND2xp5_ASAP7_75t_L g7429 ( 
.A(n_7264),
.B(n_6842),
.Y(n_7429)
);

AND2x2_ASAP7_75t_L g7430 ( 
.A(n_7171),
.B(n_6897),
.Y(n_7430)
);

INVx2_ASAP7_75t_L g7431 ( 
.A(n_7304),
.Y(n_7431)
);

AND2x4_ASAP7_75t_L g7432 ( 
.A(n_7204),
.B(n_7215),
.Y(n_7432)
);

AND2x2_ASAP7_75t_L g7433 ( 
.A(n_7269),
.B(n_6897),
.Y(n_7433)
);

HB1xp67_ASAP7_75t_L g7434 ( 
.A(n_7291),
.Y(n_7434)
);

NOR2xp33_ASAP7_75t_L g7435 ( 
.A(n_7157),
.B(n_7057),
.Y(n_7435)
);

INVx1_ASAP7_75t_L g7436 ( 
.A(n_7195),
.Y(n_7436)
);

NAND2xp5_ASAP7_75t_L g7437 ( 
.A(n_7274),
.B(n_6842),
.Y(n_7437)
);

INVx1_ASAP7_75t_SL g7438 ( 
.A(n_7181),
.Y(n_7438)
);

OR2x2_ASAP7_75t_L g7439 ( 
.A(n_7116),
.B(n_7065),
.Y(n_7439)
);

AND2x2_ASAP7_75t_L g7440 ( 
.A(n_7275),
.B(n_7040),
.Y(n_7440)
);

AND2x2_ASAP7_75t_L g7441 ( 
.A(n_7262),
.B(n_7040),
.Y(n_7441)
);

INVx1_ASAP7_75t_L g7442 ( 
.A(n_7195),
.Y(n_7442)
);

INVx2_ASAP7_75t_L g7443 ( 
.A(n_7234),
.Y(n_7443)
);

AND2x2_ASAP7_75t_L g7444 ( 
.A(n_7278),
.B(n_7044),
.Y(n_7444)
);

NAND2xp5_ASAP7_75t_L g7445 ( 
.A(n_7284),
.B(n_7065),
.Y(n_7445)
);

INVx1_ASAP7_75t_L g7446 ( 
.A(n_7319),
.Y(n_7446)
);

INVx2_ASAP7_75t_L g7447 ( 
.A(n_7234),
.Y(n_7447)
);

AND2x2_ASAP7_75t_L g7448 ( 
.A(n_7212),
.B(n_7044),
.Y(n_7448)
);

CKINVDCx16_ASAP7_75t_R g7449 ( 
.A(n_7099),
.Y(n_7449)
);

AND2x2_ASAP7_75t_L g7450 ( 
.A(n_7113),
.B(n_6898),
.Y(n_7450)
);

OR2x2_ASAP7_75t_L g7451 ( 
.A(n_7116),
.B(n_6979),
.Y(n_7451)
);

AND2x2_ASAP7_75t_L g7452 ( 
.A(n_7096),
.B(n_6898),
.Y(n_7452)
);

NAND2xp5_ASAP7_75t_L g7453 ( 
.A(n_7309),
.B(n_6946),
.Y(n_7453)
);

AND2x2_ASAP7_75t_L g7454 ( 
.A(n_7170),
.B(n_6946),
.Y(n_7454)
);

INVx1_ASAP7_75t_L g7455 ( 
.A(n_7319),
.Y(n_7455)
);

INVx2_ASAP7_75t_L g7456 ( 
.A(n_7134),
.Y(n_7456)
);

INVx2_ASAP7_75t_L g7457 ( 
.A(n_7124),
.Y(n_7457)
);

INVx1_ASAP7_75t_L g7458 ( 
.A(n_7147),
.Y(n_7458)
);

AND2x2_ASAP7_75t_L g7459 ( 
.A(n_7203),
.B(n_6950),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7156),
.Y(n_7460)
);

INVx1_ASAP7_75t_SL g7461 ( 
.A(n_7268),
.Y(n_7461)
);

AND2x4_ASAP7_75t_L g7462 ( 
.A(n_7300),
.B(n_7279),
.Y(n_7462)
);

AND2x2_ASAP7_75t_L g7463 ( 
.A(n_7210),
.B(n_6950),
.Y(n_7463)
);

NAND2xp5_ASAP7_75t_L g7464 ( 
.A(n_7260),
.B(n_7014),
.Y(n_7464)
);

AND2x2_ASAP7_75t_L g7465 ( 
.A(n_7167),
.B(n_7019),
.Y(n_7465)
);

INVx1_ASAP7_75t_L g7466 ( 
.A(n_7117),
.Y(n_7466)
);

OR2x2_ASAP7_75t_L g7467 ( 
.A(n_7117),
.B(n_6892),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_7133),
.Y(n_7468)
);

AND2x2_ASAP7_75t_L g7469 ( 
.A(n_7094),
.B(n_6953),
.Y(n_7469)
);

INVx1_ASAP7_75t_L g7470 ( 
.A(n_7133),
.Y(n_7470)
);

INVx1_ASAP7_75t_L g7471 ( 
.A(n_7291),
.Y(n_7471)
);

AND2x2_ASAP7_75t_L g7472 ( 
.A(n_7270),
.B(n_6953),
.Y(n_7472)
);

INVxp67_ASAP7_75t_L g7473 ( 
.A(n_7143),
.Y(n_7473)
);

OR2x2_ASAP7_75t_L g7474 ( 
.A(n_7266),
.B(n_6881),
.Y(n_7474)
);

NAND2xp5_ASAP7_75t_L g7475 ( 
.A(n_7288),
.B(n_6816),
.Y(n_7475)
);

OR2x2_ASAP7_75t_L g7476 ( 
.A(n_7318),
.B(n_6806),
.Y(n_7476)
);

NAND2xp5_ASAP7_75t_L g7477 ( 
.A(n_7293),
.B(n_6824),
.Y(n_7477)
);

AND2x4_ASAP7_75t_SL g7478 ( 
.A(n_7151),
.B(n_6949),
.Y(n_7478)
);

INVx1_ASAP7_75t_L g7479 ( 
.A(n_7321),
.Y(n_7479)
);

HB1xp67_ASAP7_75t_L g7480 ( 
.A(n_7321),
.Y(n_7480)
);

AND2x2_ASAP7_75t_L g7481 ( 
.A(n_7211),
.B(n_6824),
.Y(n_7481)
);

AND2x2_ASAP7_75t_L g7482 ( 
.A(n_7216),
.B(n_6989),
.Y(n_7482)
);

INVx2_ASAP7_75t_L g7483 ( 
.A(n_7124),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_7352),
.Y(n_7484)
);

INVx1_ASAP7_75t_L g7485 ( 
.A(n_7352),
.Y(n_7485)
);

NAND2xp5_ASAP7_75t_L g7486 ( 
.A(n_7299),
.B(n_6925),
.Y(n_7486)
);

NAND2xp5_ASAP7_75t_L g7487 ( 
.A(n_7306),
.B(n_6942),
.Y(n_7487)
);

OR2x2_ASAP7_75t_L g7488 ( 
.A(n_7159),
.B(n_6865),
.Y(n_7488)
);

AND2x2_ASAP7_75t_L g7489 ( 
.A(n_7314),
.B(n_6989),
.Y(n_7489)
);

INVx4_ASAP7_75t_L g7490 ( 
.A(n_7248),
.Y(n_7490)
);

INVx1_ASAP7_75t_L g7491 ( 
.A(n_7355),
.Y(n_7491)
);

INVx2_ASAP7_75t_L g7492 ( 
.A(n_7249),
.Y(n_7492)
);

OR2x2_ASAP7_75t_L g7493 ( 
.A(n_7159),
.B(n_6992),
.Y(n_7493)
);

AND2x2_ASAP7_75t_L g7494 ( 
.A(n_7131),
.B(n_6990),
.Y(n_7494)
);

NAND2xp5_ASAP7_75t_L g7495 ( 
.A(n_7183),
.B(n_7037),
.Y(n_7495)
);

AND2x2_ASAP7_75t_L g7496 ( 
.A(n_7317),
.B(n_6990),
.Y(n_7496)
);

AND2x2_ASAP7_75t_L g7497 ( 
.A(n_7326),
.B(n_6847),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_7355),
.Y(n_7498)
);

INVx3_ASAP7_75t_L g7499 ( 
.A(n_7249),
.Y(n_7499)
);

INVxp67_ASAP7_75t_SL g7500 ( 
.A(n_7107),
.Y(n_7500)
);

INVx1_ASAP7_75t_SL g7501 ( 
.A(n_7140),
.Y(n_7501)
);

AND2x2_ASAP7_75t_L g7502 ( 
.A(n_7332),
.B(n_6847),
.Y(n_7502)
);

INVx2_ASAP7_75t_L g7503 ( 
.A(n_7259),
.Y(n_7503)
);

AND2x2_ASAP7_75t_L g7504 ( 
.A(n_7335),
.B(n_7020),
.Y(n_7504)
);

INVx5_ASAP7_75t_L g7505 ( 
.A(n_7248),
.Y(n_7505)
);

INVx2_ASAP7_75t_L g7506 ( 
.A(n_7259),
.Y(n_7506)
);

AND2x2_ASAP7_75t_L g7507 ( 
.A(n_7342),
.B(n_7346),
.Y(n_7507)
);

NOR2xp33_ASAP7_75t_L g7508 ( 
.A(n_7283),
.B(n_6845),
.Y(n_7508)
);

AND2x2_ASAP7_75t_L g7509 ( 
.A(n_7349),
.B(n_7020),
.Y(n_7509)
);

OR2x2_ASAP7_75t_L g7510 ( 
.A(n_7191),
.B(n_6888),
.Y(n_7510)
);

AND2x2_ASAP7_75t_L g7511 ( 
.A(n_7353),
.B(n_7021),
.Y(n_7511)
);

INVx1_ASAP7_75t_SL g7512 ( 
.A(n_7151),
.Y(n_7512)
);

AND2x2_ASAP7_75t_L g7513 ( 
.A(n_7354),
.B(n_7021),
.Y(n_7513)
);

AND2x2_ASAP7_75t_L g7514 ( 
.A(n_7303),
.B(n_7022),
.Y(n_7514)
);

NAND2xp5_ASAP7_75t_L g7515 ( 
.A(n_7183),
.B(n_7022),
.Y(n_7515)
);

INVx1_ASAP7_75t_L g7516 ( 
.A(n_7359),
.Y(n_7516)
);

INVx1_ASAP7_75t_L g7517 ( 
.A(n_7109),
.Y(n_7517)
);

AND2x2_ASAP7_75t_L g7518 ( 
.A(n_7303),
.B(n_7033),
.Y(n_7518)
);

NOR2xp33_ASAP7_75t_L g7519 ( 
.A(n_7283),
.B(n_6819),
.Y(n_7519)
);

AND2x2_ASAP7_75t_L g7520 ( 
.A(n_7327),
.B(n_7033),
.Y(n_7520)
);

AND2x4_ASAP7_75t_L g7521 ( 
.A(n_7093),
.B(n_6935),
.Y(n_7521)
);

AND2x2_ASAP7_75t_L g7522 ( 
.A(n_7327),
.B(n_7036),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7115),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_7118),
.Y(n_7524)
);

NAND2xp5_ASAP7_75t_L g7525 ( 
.A(n_7185),
.B(n_7036),
.Y(n_7525)
);

NAND2xp5_ASAP7_75t_L g7526 ( 
.A(n_7185),
.B(n_7039),
.Y(n_7526)
);

A2O1A1Ixp33_ASAP7_75t_SL g7527 ( 
.A1(n_7088),
.A2(n_7139),
.B(n_7125),
.C(n_7271),
.Y(n_7527)
);

AND2x4_ASAP7_75t_L g7528 ( 
.A(n_7089),
.B(n_6849),
.Y(n_7528)
);

AND2x4_ASAP7_75t_L g7529 ( 
.A(n_7089),
.B(n_6849),
.Y(n_7529)
);

INVx1_ASAP7_75t_SL g7530 ( 
.A(n_7169),
.Y(n_7530)
);

AND2x2_ASAP7_75t_L g7531 ( 
.A(n_7209),
.B(n_7000),
.Y(n_7531)
);

AND2x4_ASAP7_75t_L g7532 ( 
.A(n_7292),
.B(n_6851),
.Y(n_7532)
);

INVx1_ASAP7_75t_L g7533 ( 
.A(n_7121),
.Y(n_7533)
);

AND2x2_ASAP7_75t_L g7534 ( 
.A(n_7347),
.B(n_7039),
.Y(n_7534)
);

INVx2_ASAP7_75t_L g7535 ( 
.A(n_7292),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7180),
.Y(n_7536)
);

AND2x4_ASAP7_75t_L g7537 ( 
.A(n_7311),
.B(n_6851),
.Y(n_7537)
);

AND2x2_ASAP7_75t_L g7538 ( 
.A(n_7348),
.B(n_7048),
.Y(n_7538)
);

AND2x2_ASAP7_75t_L g7539 ( 
.A(n_7209),
.B(n_7048),
.Y(n_7539)
);

AND2x2_ASAP7_75t_L g7540 ( 
.A(n_7209),
.B(n_7169),
.Y(n_7540)
);

NAND2xp5_ASAP7_75t_L g7541 ( 
.A(n_7218),
.B(n_7049),
.Y(n_7541)
);

AND2x2_ASAP7_75t_L g7542 ( 
.A(n_7179),
.B(n_7241),
.Y(n_7542)
);

INVx1_ASAP7_75t_L g7543 ( 
.A(n_7187),
.Y(n_7543)
);

AND2x2_ASAP7_75t_L g7544 ( 
.A(n_7179),
.B(n_7049),
.Y(n_7544)
);

INVx2_ASAP7_75t_L g7545 ( 
.A(n_7311),
.Y(n_7545)
);

INVx1_ASAP7_75t_L g7546 ( 
.A(n_7137),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_7138),
.Y(n_7547)
);

INVx1_ASAP7_75t_L g7548 ( 
.A(n_7141),
.Y(n_7548)
);

NOR2xp67_ASAP7_75t_L g7549 ( 
.A(n_7218),
.B(n_6981),
.Y(n_7549)
);

INVx1_ASAP7_75t_L g7550 ( 
.A(n_7267),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7267),
.Y(n_7551)
);

INVx1_ASAP7_75t_SL g7552 ( 
.A(n_7301),
.Y(n_7552)
);

INVx2_ASAP7_75t_SL g7553 ( 
.A(n_7130),
.Y(n_7553)
);

INVx1_ASAP7_75t_L g7554 ( 
.A(n_7281),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_L g7555 ( 
.A(n_7120),
.B(n_7060),
.Y(n_7555)
);

HB1xp67_ASAP7_75t_L g7556 ( 
.A(n_7282),
.Y(n_7556)
);

OR2x6_ASAP7_75t_SL g7557 ( 
.A(n_7153),
.B(n_7060),
.Y(n_7557)
);

INVx2_ASAP7_75t_L g7558 ( 
.A(n_7130),
.Y(n_7558)
);

INVx1_ASAP7_75t_L g7559 ( 
.A(n_7281),
.Y(n_7559)
);

INVx2_ASAP7_75t_L g7560 ( 
.A(n_7160),
.Y(n_7560)
);

AND2x4_ASAP7_75t_L g7561 ( 
.A(n_7182),
.B(n_7000),
.Y(n_7561)
);

INVx2_ASAP7_75t_L g7562 ( 
.A(n_7184),
.Y(n_7562)
);

BUFx2_ASAP7_75t_L g7563 ( 
.A(n_7120),
.Y(n_7563)
);

INVx1_ASAP7_75t_L g7564 ( 
.A(n_7334),
.Y(n_7564)
);

INVx2_ASAP7_75t_L g7565 ( 
.A(n_7220),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7241),
.B(n_7032),
.Y(n_7566)
);

HB1xp67_ASAP7_75t_L g7567 ( 
.A(n_7282),
.Y(n_7567)
);

NOR2xp33_ASAP7_75t_L g7568 ( 
.A(n_7153),
.B(n_6815),
.Y(n_7568)
);

AND2x2_ASAP7_75t_L g7569 ( 
.A(n_7186),
.B(n_7032),
.Y(n_7569)
);

AND2x2_ASAP7_75t_SL g7570 ( 
.A(n_7240),
.B(n_7090),
.Y(n_7570)
);

INVx2_ASAP7_75t_L g7571 ( 
.A(n_7263),
.Y(n_7571)
);

INVx1_ASAP7_75t_L g7572 ( 
.A(n_7257),
.Y(n_7572)
);

INVx2_ASAP7_75t_L g7573 ( 
.A(n_7280),
.Y(n_7573)
);

AND2x2_ASAP7_75t_L g7574 ( 
.A(n_7186),
.B(n_7034),
.Y(n_7574)
);

OR2x2_ASAP7_75t_L g7575 ( 
.A(n_7192),
.B(n_6862),
.Y(n_7575)
);

INVx1_ASAP7_75t_L g7576 ( 
.A(n_7258),
.Y(n_7576)
);

AND2x2_ASAP7_75t_L g7577 ( 
.A(n_7168),
.B(n_7034),
.Y(n_7577)
);

HB1xp67_ASAP7_75t_L g7578 ( 
.A(n_7294),
.Y(n_7578)
);

AND2x2_ASAP7_75t_L g7579 ( 
.A(n_7175),
.B(n_7029),
.Y(n_7579)
);

HB1xp67_ASAP7_75t_L g7580 ( 
.A(n_7296),
.Y(n_7580)
);

AND2x2_ASAP7_75t_L g7581 ( 
.A(n_7177),
.B(n_7029),
.Y(n_7581)
);

OR2x2_ASAP7_75t_L g7582 ( 
.A(n_7197),
.B(n_6960),
.Y(n_7582)
);

AND2x2_ASAP7_75t_L g7583 ( 
.A(n_7178),
.B(n_7030),
.Y(n_7583)
);

AND2x2_ASAP7_75t_L g7584 ( 
.A(n_7114),
.B(n_7030),
.Y(n_7584)
);

AND2x2_ASAP7_75t_L g7585 ( 
.A(n_7129),
.B(n_6957),
.Y(n_7585)
);

NAND2xp5_ASAP7_75t_L g7586 ( 
.A(n_7297),
.B(n_6957),
.Y(n_7586)
);

OR2x2_ASAP7_75t_L g7587 ( 
.A(n_7155),
.B(n_7012),
.Y(n_7587)
);

NOR2xp33_ASAP7_75t_L g7588 ( 
.A(n_7221),
.B(n_7163),
.Y(n_7588)
);

INVx2_ASAP7_75t_L g7589 ( 
.A(n_7305),
.Y(n_7589)
);

OR2x2_ASAP7_75t_L g7590 ( 
.A(n_7090),
.B(n_7050),
.Y(n_7590)
);

INVxp67_ASAP7_75t_SL g7591 ( 
.A(n_7329),
.Y(n_7591)
);

INVx2_ASAP7_75t_SL g7592 ( 
.A(n_7310),
.Y(n_7592)
);

NOR2xp33_ASAP7_75t_L g7593 ( 
.A(n_7297),
.B(n_6930),
.Y(n_7593)
);

AND2x2_ASAP7_75t_L g7594 ( 
.A(n_7097),
.B(n_7000),
.Y(n_7594)
);

NAND2xp5_ASAP7_75t_L g7595 ( 
.A(n_7098),
.B(n_6964),
.Y(n_7595)
);

OR2x2_ASAP7_75t_L g7596 ( 
.A(n_7265),
.B(n_7046),
.Y(n_7596)
);

INVx2_ASAP7_75t_L g7597 ( 
.A(n_7320),
.Y(n_7597)
);

INVx2_ASAP7_75t_L g7598 ( 
.A(n_7158),
.Y(n_7598)
);

AND2x2_ASAP7_75t_L g7599 ( 
.A(n_7100),
.B(n_7004),
.Y(n_7599)
);

INVx2_ASAP7_75t_L g7600 ( 
.A(n_7176),
.Y(n_7600)
);

INVx2_ASAP7_75t_L g7601 ( 
.A(n_7188),
.Y(n_7601)
);

INVx1_ASAP7_75t_L g7602 ( 
.A(n_7277),
.Y(n_7602)
);

AND2x2_ASAP7_75t_L g7603 ( 
.A(n_7108),
.B(n_7004),
.Y(n_7603)
);

INVx2_ASAP7_75t_L g7604 ( 
.A(n_7207),
.Y(n_7604)
);

INVx2_ASAP7_75t_L g7605 ( 
.A(n_7214),
.Y(n_7605)
);

INVxp67_ASAP7_75t_SL g7606 ( 
.A(n_7329),
.Y(n_7606)
);

HB1xp67_ASAP7_75t_L g7607 ( 
.A(n_7549),
.Y(n_7607)
);

NOR2xp67_ASAP7_75t_L g7608 ( 
.A(n_7372),
.B(n_6981),
.Y(n_7608)
);

INVx1_ASAP7_75t_L g7609 ( 
.A(n_7386),
.Y(n_7609)
);

INVx1_ASAP7_75t_L g7610 ( 
.A(n_7386),
.Y(n_7610)
);

AND2x4_ASAP7_75t_L g7611 ( 
.A(n_7521),
.B(n_7091),
.Y(n_7611)
);

INVx2_ASAP7_75t_L g7612 ( 
.A(n_7432),
.Y(n_7612)
);

INVx1_ASAP7_75t_L g7613 ( 
.A(n_7427),
.Y(n_7613)
);

AND2x2_ASAP7_75t_L g7614 ( 
.A(n_7388),
.B(n_7092),
.Y(n_7614)
);

AND2x2_ASAP7_75t_L g7615 ( 
.A(n_7542),
.B(n_7128),
.Y(n_7615)
);

NAND2xp5_ASAP7_75t_L g7616 ( 
.A(n_7367),
.B(n_7135),
.Y(n_7616)
);

AND2x2_ASAP7_75t_L g7617 ( 
.A(n_7373),
.B(n_7136),
.Y(n_7617)
);

HB1xp67_ASAP7_75t_L g7618 ( 
.A(n_7432),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7427),
.Y(n_7619)
);

OR2x2_ASAP7_75t_L g7620 ( 
.A(n_7361),
.B(n_7208),
.Y(n_7620)
);

INVx2_ASAP7_75t_L g7621 ( 
.A(n_7432),
.Y(n_7621)
);

INVx1_ASAP7_75t_L g7622 ( 
.A(n_7556),
.Y(n_7622)
);

INVx1_ASAP7_75t_L g7623 ( 
.A(n_7556),
.Y(n_7623)
);

INVx1_ASAP7_75t_L g7624 ( 
.A(n_7567),
.Y(n_7624)
);

NAND2xp5_ASAP7_75t_L g7625 ( 
.A(n_7367),
.B(n_7287),
.Y(n_7625)
);

AND2x4_ASAP7_75t_L g7626 ( 
.A(n_7521),
.B(n_7219),
.Y(n_7626)
);

NAND2xp5_ASAP7_75t_L g7627 ( 
.A(n_7370),
.B(n_7289),
.Y(n_7627)
);

AND2x2_ASAP7_75t_L g7628 ( 
.A(n_7448),
.B(n_7253),
.Y(n_7628)
);

HB1xp67_ASAP7_75t_SL g7629 ( 
.A(n_7370),
.Y(n_7629)
);

HB1xp67_ASAP7_75t_L g7630 ( 
.A(n_7361),
.Y(n_7630)
);

AND2x2_ASAP7_75t_L g7631 ( 
.A(n_7448),
.B(n_7322),
.Y(n_7631)
);

INVx1_ASAP7_75t_L g7632 ( 
.A(n_7567),
.Y(n_7632)
);

AND2x2_ASAP7_75t_L g7633 ( 
.A(n_7452),
.B(n_7324),
.Y(n_7633)
);

INVx1_ASAP7_75t_SL g7634 ( 
.A(n_7557),
.Y(n_7634)
);

AND2x2_ASAP7_75t_L g7635 ( 
.A(n_7452),
.B(n_7338),
.Y(n_7635)
);

INVx2_ASAP7_75t_L g7636 ( 
.A(n_7372),
.Y(n_7636)
);

OR2x2_ASAP7_75t_L g7637 ( 
.A(n_7449),
.B(n_7208),
.Y(n_7637)
);

AND2x2_ASAP7_75t_L g7638 ( 
.A(n_7450),
.B(n_7339),
.Y(n_7638)
);

INVx2_ASAP7_75t_L g7639 ( 
.A(n_7372),
.Y(n_7639)
);

NAND2xp5_ASAP7_75t_L g7640 ( 
.A(n_7591),
.B(n_7295),
.Y(n_7640)
);

AND2x2_ASAP7_75t_L g7641 ( 
.A(n_7450),
.B(n_7368),
.Y(n_7641)
);

NAND2xp5_ASAP7_75t_L g7642 ( 
.A(n_7591),
.B(n_7606),
.Y(n_7642)
);

AND2x2_ASAP7_75t_L g7643 ( 
.A(n_7368),
.B(n_6964),
.Y(n_7643)
);

HB1xp67_ASAP7_75t_L g7644 ( 
.A(n_7505),
.Y(n_7644)
);

INVx1_ASAP7_75t_L g7645 ( 
.A(n_7578),
.Y(n_7645)
);

OR2x2_ASAP7_75t_L g7646 ( 
.A(n_7512),
.B(n_7110),
.Y(n_7646)
);

INVx2_ASAP7_75t_SL g7647 ( 
.A(n_7400),
.Y(n_7647)
);

OR2x2_ASAP7_75t_L g7648 ( 
.A(n_7530),
.B(n_7132),
.Y(n_7648)
);

AND2x2_ASAP7_75t_L g7649 ( 
.A(n_7416),
.B(n_7069),
.Y(n_7649)
);

INVx1_ASAP7_75t_L g7650 ( 
.A(n_7578),
.Y(n_7650)
);

AND2x2_ASAP7_75t_L g7651 ( 
.A(n_7382),
.B(n_7069),
.Y(n_7651)
);

NAND2xp5_ASAP7_75t_L g7652 ( 
.A(n_7606),
.B(n_7557),
.Y(n_7652)
);

OR2x2_ASAP7_75t_L g7653 ( 
.A(n_7422),
.B(n_7152),
.Y(n_7653)
);

NAND2xp5_ASAP7_75t_L g7654 ( 
.A(n_7588),
.B(n_7308),
.Y(n_7654)
);

AND2x2_ASAP7_75t_L g7655 ( 
.A(n_7382),
.B(n_7072),
.Y(n_7655)
);

OR2x2_ASAP7_75t_L g7656 ( 
.A(n_7371),
.B(n_7103),
.Y(n_7656)
);

OR2x2_ASAP7_75t_L g7657 ( 
.A(n_7389),
.B(n_7103),
.Y(n_7657)
);

INVx1_ASAP7_75t_L g7658 ( 
.A(n_7580),
.Y(n_7658)
);

INVxp67_ASAP7_75t_L g7659 ( 
.A(n_7360),
.Y(n_7659)
);

OR2x2_ASAP7_75t_L g7660 ( 
.A(n_7408),
.B(n_7112),
.Y(n_7660)
);

AND2x2_ASAP7_75t_SL g7661 ( 
.A(n_7570),
.B(n_7205),
.Y(n_7661)
);

AND2x2_ASAP7_75t_L g7662 ( 
.A(n_7454),
.B(n_7072),
.Y(n_7662)
);

INVx1_ASAP7_75t_L g7663 ( 
.A(n_7580),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7419),
.Y(n_7664)
);

NAND2xp5_ASAP7_75t_L g7665 ( 
.A(n_7588),
.B(n_7312),
.Y(n_7665)
);

AND2x2_ASAP7_75t_L g7666 ( 
.A(n_7454),
.B(n_6896),
.Y(n_7666)
);

INVx2_ASAP7_75t_L g7667 ( 
.A(n_7499),
.Y(n_7667)
);

OR2x2_ASAP7_75t_L g7668 ( 
.A(n_7461),
.B(n_7112),
.Y(n_7668)
);

NOR2x1_ASAP7_75t_L g7669 ( 
.A(n_7499),
.B(n_6930),
.Y(n_7669)
);

NAND2xp5_ASAP7_75t_L g7670 ( 
.A(n_7570),
.B(n_7369),
.Y(n_7670)
);

INVx1_ASAP7_75t_L g7671 ( 
.A(n_7419),
.Y(n_7671)
);

INVx1_ASAP7_75t_L g7672 ( 
.A(n_7431),
.Y(n_7672)
);

HB1xp67_ASAP7_75t_L g7673 ( 
.A(n_7505),
.Y(n_7673)
);

NAND2xp5_ASAP7_75t_L g7674 ( 
.A(n_7527),
.B(n_7313),
.Y(n_7674)
);

OR2x2_ASAP7_75t_L g7675 ( 
.A(n_7437),
.B(n_7325),
.Y(n_7675)
);

INVx1_ASAP7_75t_L g7676 ( 
.A(n_7431),
.Y(n_7676)
);

AND2x4_ASAP7_75t_L g7677 ( 
.A(n_7521),
.B(n_7499),
.Y(n_7677)
);

INVx2_ASAP7_75t_L g7678 ( 
.A(n_7505),
.Y(n_7678)
);

INVx2_ASAP7_75t_L g7679 ( 
.A(n_7505),
.Y(n_7679)
);

AND2x2_ASAP7_75t_L g7680 ( 
.A(n_7440),
.B(n_7200),
.Y(n_7680)
);

AND2x2_ASAP7_75t_L g7681 ( 
.A(n_7440),
.B(n_7316),
.Y(n_7681)
);

NAND2xp5_ASAP7_75t_L g7682 ( 
.A(n_7527),
.B(n_7333),
.Y(n_7682)
);

INVxp67_ASAP7_75t_SL g7683 ( 
.A(n_7582),
.Y(n_7683)
);

NAND2xp5_ASAP7_75t_L g7684 ( 
.A(n_7444),
.B(n_7336),
.Y(n_7684)
);

INVxp67_ASAP7_75t_L g7685 ( 
.A(n_7360),
.Y(n_7685)
);

INVxp33_ASAP7_75t_L g7686 ( 
.A(n_7413),
.Y(n_7686)
);

NAND2xp5_ASAP7_75t_L g7687 ( 
.A(n_7444),
.B(n_7161),
.Y(n_7687)
);

AND2x2_ASAP7_75t_L g7688 ( 
.A(n_7459),
.B(n_6949),
.Y(n_7688)
);

AND2x2_ASAP7_75t_L g7689 ( 
.A(n_7463),
.B(n_6949),
.Y(n_7689)
);

AND2x4_ASAP7_75t_L g7690 ( 
.A(n_7400),
.B(n_6949),
.Y(n_7690)
);

INVx2_ASAP7_75t_L g7691 ( 
.A(n_7418),
.Y(n_7691)
);

INVxp67_ASAP7_75t_L g7692 ( 
.A(n_7398),
.Y(n_7692)
);

AND2x2_ASAP7_75t_L g7693 ( 
.A(n_7441),
.B(n_6884),
.Y(n_7693)
);

INVx1_ASAP7_75t_L g7694 ( 
.A(n_7446),
.Y(n_7694)
);

INVx2_ASAP7_75t_L g7695 ( 
.A(n_7418),
.Y(n_7695)
);

AND2x2_ASAP7_75t_L g7696 ( 
.A(n_7441),
.B(n_6886),
.Y(n_7696)
);

OR2x2_ASAP7_75t_L g7697 ( 
.A(n_7445),
.B(n_7325),
.Y(n_7697)
);

INVx1_ASAP7_75t_L g7698 ( 
.A(n_7455),
.Y(n_7698)
);

OR2x2_ASAP7_75t_L g7699 ( 
.A(n_7586),
.B(n_7364),
.Y(n_7699)
);

AND2x4_ASAP7_75t_L g7700 ( 
.A(n_7462),
.B(n_7004),
.Y(n_7700)
);

AND2x4_ASAP7_75t_SL g7701 ( 
.A(n_7494),
.B(n_6930),
.Y(n_7701)
);

OR2x2_ASAP7_75t_L g7702 ( 
.A(n_7429),
.B(n_7425),
.Y(n_7702)
);

INVx3_ASAP7_75t_L g7703 ( 
.A(n_7462),
.Y(n_7703)
);

AND2x4_ASAP7_75t_L g7704 ( 
.A(n_7462),
.B(n_7059),
.Y(n_7704)
);

INVx2_ASAP7_75t_L g7705 ( 
.A(n_7478),
.Y(n_7705)
);

AND2x2_ASAP7_75t_L g7706 ( 
.A(n_7387),
.B(n_6887),
.Y(n_7706)
);

OR2x2_ASAP7_75t_L g7707 ( 
.A(n_7412),
.B(n_7164),
.Y(n_7707)
);

INVx1_ASAP7_75t_SL g7708 ( 
.A(n_7478),
.Y(n_7708)
);

INVx1_ASAP7_75t_L g7709 ( 
.A(n_7550),
.Y(n_7709)
);

INVx2_ASAP7_75t_L g7710 ( 
.A(n_7363),
.Y(n_7710)
);

NAND2xp67_ASAP7_75t_L g7711 ( 
.A(n_7540),
.B(n_7251),
.Y(n_7711)
);

AO22x1_ASAP7_75t_L g7712 ( 
.A1(n_7500),
.A2(n_7254),
.B1(n_7302),
.B2(n_7162),
.Y(n_7712)
);

INVx2_ASAP7_75t_L g7713 ( 
.A(n_7363),
.Y(n_7713)
);

INVx2_ASAP7_75t_L g7714 ( 
.A(n_7363),
.Y(n_7714)
);

INVx1_ASAP7_75t_L g7715 ( 
.A(n_7551),
.Y(n_7715)
);

AND2x2_ASAP7_75t_L g7716 ( 
.A(n_7428),
.B(n_6890),
.Y(n_7716)
);

INVx2_ASAP7_75t_L g7717 ( 
.A(n_7532),
.Y(n_7717)
);

NAND2xp5_ASAP7_75t_L g7718 ( 
.A(n_7500),
.B(n_7161),
.Y(n_7718)
);

AND2x4_ASAP7_75t_L g7719 ( 
.A(n_7532),
.B(n_7537),
.Y(n_7719)
);

OR2x2_ASAP7_75t_L g7720 ( 
.A(n_7420),
.B(n_7164),
.Y(n_7720)
);

AOI22xp33_ASAP7_75t_SL g7721 ( 
.A1(n_7566),
.A2(n_7302),
.B1(n_7254),
.B2(n_7315),
.Y(n_7721)
);

AOI22xp33_ASAP7_75t_L g7722 ( 
.A1(n_7417),
.A2(n_7315),
.B1(n_6644),
.B2(n_6562),
.Y(n_7722)
);

NAND2xp5_ASAP7_75t_L g7723 ( 
.A(n_7395),
.B(n_7162),
.Y(n_7723)
);

INVx1_ASAP7_75t_L g7724 ( 
.A(n_7554),
.Y(n_7724)
);

AND2x2_ASAP7_75t_L g7725 ( 
.A(n_7423),
.B(n_6893),
.Y(n_7725)
);

INVx2_ASAP7_75t_L g7726 ( 
.A(n_7532),
.Y(n_7726)
);

NAND2xp5_ASAP7_75t_L g7727 ( 
.A(n_7395),
.B(n_6891),
.Y(n_7727)
);

INVx1_ASAP7_75t_L g7728 ( 
.A(n_7559),
.Y(n_7728)
);

OR2x2_ASAP7_75t_L g7729 ( 
.A(n_7439),
.B(n_7451),
.Y(n_7729)
);

NAND2xp5_ASAP7_75t_L g7730 ( 
.A(n_7397),
.B(n_7222),
.Y(n_7730)
);

NAND2x1p5_ASAP7_75t_L g7731 ( 
.A(n_7490),
.B(n_7058),
.Y(n_7731)
);

HB1xp67_ASAP7_75t_L g7732 ( 
.A(n_7434),
.Y(n_7732)
);

INVx1_ASAP7_75t_L g7733 ( 
.A(n_7406),
.Y(n_7733)
);

HB1xp67_ASAP7_75t_L g7734 ( 
.A(n_7381),
.Y(n_7734)
);

NAND2xp5_ASAP7_75t_L g7735 ( 
.A(n_7397),
.B(n_7225),
.Y(n_7735)
);

NOR2xp33_ASAP7_75t_L g7736 ( 
.A(n_7501),
.B(n_7273),
.Y(n_7736)
);

HB1xp67_ASAP7_75t_L g7737 ( 
.A(n_7381),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_7421),
.Y(n_7738)
);

INVx1_ASAP7_75t_L g7739 ( 
.A(n_7424),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_7426),
.Y(n_7740)
);

AND2x2_ASAP7_75t_SL g7741 ( 
.A(n_7417),
.B(n_7469),
.Y(n_7741)
);

INVx2_ASAP7_75t_L g7742 ( 
.A(n_7537),
.Y(n_7742)
);

AND2x2_ASAP7_75t_L g7743 ( 
.A(n_7423),
.B(n_7228),
.Y(n_7743)
);

INVx4_ASAP7_75t_L g7744 ( 
.A(n_7490),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7436),
.Y(n_7745)
);

OR2x2_ASAP7_75t_L g7746 ( 
.A(n_7402),
.B(n_7165),
.Y(n_7746)
);

AND2x2_ASAP7_75t_L g7747 ( 
.A(n_7365),
.B(n_7230),
.Y(n_7747)
);

AND2x2_ASAP7_75t_L g7748 ( 
.A(n_7465),
.B(n_7246),
.Y(n_7748)
);

AND2x2_ASAP7_75t_L g7749 ( 
.A(n_7433),
.B(n_7252),
.Y(n_7749)
);

INVx1_ASAP7_75t_L g7750 ( 
.A(n_7442),
.Y(n_7750)
);

AND2x2_ASAP7_75t_L g7751 ( 
.A(n_7394),
.B(n_6623),
.Y(n_7751)
);

INVx1_ASAP7_75t_SL g7752 ( 
.A(n_7472),
.Y(n_7752)
);

AND2x2_ASAP7_75t_L g7753 ( 
.A(n_7394),
.B(n_6623),
.Y(n_7753)
);

INVx1_ASAP7_75t_SL g7754 ( 
.A(n_7414),
.Y(n_7754)
);

INVx1_ASAP7_75t_L g7755 ( 
.A(n_7535),
.Y(n_7755)
);

INVx1_ASAP7_75t_L g7756 ( 
.A(n_7535),
.Y(n_7756)
);

HB1xp67_ASAP7_75t_L g7757 ( 
.A(n_7404),
.Y(n_7757)
);

INVx1_ASAP7_75t_L g7758 ( 
.A(n_7545),
.Y(n_7758)
);

AND2x2_ASAP7_75t_L g7759 ( 
.A(n_7396),
.B(n_7165),
.Y(n_7759)
);

AND2x2_ASAP7_75t_L g7760 ( 
.A(n_7396),
.B(n_7194),
.Y(n_7760)
);

AND2x2_ASAP7_75t_L g7761 ( 
.A(n_7375),
.B(n_7194),
.Y(n_7761)
);

INVx2_ASAP7_75t_L g7762 ( 
.A(n_7537),
.Y(n_7762)
);

INVx1_ASAP7_75t_SL g7763 ( 
.A(n_7438),
.Y(n_7763)
);

OR2x2_ASAP7_75t_L g7764 ( 
.A(n_7475),
.B(n_7226),
.Y(n_7764)
);

INVx6_ASAP7_75t_L g7765 ( 
.A(n_7490),
.Y(n_7765)
);

INVx1_ASAP7_75t_L g7766 ( 
.A(n_7545),
.Y(n_7766)
);

INVx1_ASAP7_75t_L g7767 ( 
.A(n_7362),
.Y(n_7767)
);

INVx2_ASAP7_75t_L g7768 ( 
.A(n_7404),
.Y(n_7768)
);

INVx1_ASAP7_75t_L g7769 ( 
.A(n_7366),
.Y(n_7769)
);

INVx1_ASAP7_75t_SL g7770 ( 
.A(n_7563),
.Y(n_7770)
);

INVx1_ASAP7_75t_L g7771 ( 
.A(n_7378),
.Y(n_7771)
);

OR2x2_ASAP7_75t_L g7772 ( 
.A(n_7477),
.B(n_7226),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_7399),
.Y(n_7773)
);

AND2x2_ASAP7_75t_L g7774 ( 
.A(n_7376),
.B(n_7231),
.Y(n_7774)
);

INVx1_ASAP7_75t_L g7775 ( 
.A(n_7401),
.Y(n_7775)
);

AND2x2_ASAP7_75t_L g7776 ( 
.A(n_7374),
.B(n_7231),
.Y(n_7776)
);

OR2x2_ASAP7_75t_L g7777 ( 
.A(n_7515),
.B(n_7232),
.Y(n_7777)
);

INVx2_ASAP7_75t_L g7778 ( 
.A(n_7405),
.Y(n_7778)
);

AND2x2_ASAP7_75t_L g7779 ( 
.A(n_7409),
.B(n_7232),
.Y(n_7779)
);

INVxp67_ASAP7_75t_SL g7780 ( 
.A(n_7415),
.Y(n_7780)
);

OR2x2_ASAP7_75t_L g7781 ( 
.A(n_7525),
.B(n_7236),
.Y(n_7781)
);

NAND2xp5_ASAP7_75t_L g7782 ( 
.A(n_7592),
.B(n_7337),
.Y(n_7782)
);

INVx1_ASAP7_75t_L g7783 ( 
.A(n_7403),
.Y(n_7783)
);

OR2x2_ASAP7_75t_L g7784 ( 
.A(n_7526),
.B(n_7236),
.Y(n_7784)
);

OR2x2_ASAP7_75t_L g7785 ( 
.A(n_7552),
.B(n_7242),
.Y(n_7785)
);

NOR2xp33_ASAP7_75t_L g7786 ( 
.A(n_7453),
.B(n_7273),
.Y(n_7786)
);

AND2x2_ASAP7_75t_L g7787 ( 
.A(n_7407),
.B(n_7242),
.Y(n_7787)
);

AND2x2_ASAP7_75t_L g7788 ( 
.A(n_7383),
.B(n_7328),
.Y(n_7788)
);

INVx1_ASAP7_75t_L g7789 ( 
.A(n_7579),
.Y(n_7789)
);

AND2x4_ASAP7_75t_L g7790 ( 
.A(n_7561),
.B(n_7059),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_7581),
.Y(n_7791)
);

NAND2xp5_ASAP7_75t_L g7792 ( 
.A(n_7592),
.B(n_7340),
.Y(n_7792)
);

AND2x2_ASAP7_75t_L g7793 ( 
.A(n_7430),
.B(n_7328),
.Y(n_7793)
);

INVx1_ASAP7_75t_L g7794 ( 
.A(n_7583),
.Y(n_7794)
);

INVx2_ASAP7_75t_L g7795 ( 
.A(n_7405),
.Y(n_7795)
);

AOI221xp5_ASAP7_75t_L g7796 ( 
.A1(n_7568),
.A2(n_7286),
.B1(n_7350),
.B2(n_7251),
.C(n_7331),
.Y(n_7796)
);

INVx1_ASAP7_75t_L g7797 ( 
.A(n_7434),
.Y(n_7797)
);

AND2x6_ASAP7_75t_SL g7798 ( 
.A(n_7391),
.B(n_7330),
.Y(n_7798)
);

INVx1_ASAP7_75t_L g7799 ( 
.A(n_7480),
.Y(n_7799)
);

AND2x2_ASAP7_75t_L g7800 ( 
.A(n_7377),
.B(n_7330),
.Y(n_7800)
);

INVxp67_ASAP7_75t_L g7801 ( 
.A(n_7593),
.Y(n_7801)
);

NAND2xp5_ASAP7_75t_L g7802 ( 
.A(n_7577),
.B(n_7341),
.Y(n_7802)
);

AND2x2_ASAP7_75t_L g7803 ( 
.A(n_7379),
.B(n_7331),
.Y(n_7803)
);

OR2x2_ASAP7_75t_L g7804 ( 
.A(n_7384),
.B(n_7298),
.Y(n_7804)
);

AND2x2_ASAP7_75t_L g7805 ( 
.A(n_7390),
.B(n_6608),
.Y(n_7805)
);

AND2x2_ASAP7_75t_L g7806 ( 
.A(n_7385),
.B(n_6608),
.Y(n_7806)
);

AND2x2_ASAP7_75t_L g7807 ( 
.A(n_7482),
.B(n_6702),
.Y(n_7807)
);

NAND2xp5_ASAP7_75t_L g7808 ( 
.A(n_7391),
.B(n_7584),
.Y(n_7808)
);

INVx1_ASAP7_75t_L g7809 ( 
.A(n_7480),
.Y(n_7809)
);

INVx2_ASAP7_75t_L g7810 ( 
.A(n_7561),
.Y(n_7810)
);

NAND2xp5_ASAP7_75t_L g7811 ( 
.A(n_7568),
.B(n_7344),
.Y(n_7811)
);

INVx1_ASAP7_75t_L g7812 ( 
.A(n_7541),
.Y(n_7812)
);

AND2x2_ASAP7_75t_L g7813 ( 
.A(n_7489),
.B(n_6702),
.Y(n_7813)
);

INVx1_ASAP7_75t_L g7814 ( 
.A(n_7555),
.Y(n_7814)
);

AND2x2_ASAP7_75t_L g7815 ( 
.A(n_7751),
.B(n_7481),
.Y(n_7815)
);

AND2x2_ASAP7_75t_L g7816 ( 
.A(n_7753),
.B(n_7496),
.Y(n_7816)
);

INVx1_ASAP7_75t_L g7817 ( 
.A(n_7732),
.Y(n_7817)
);

OR2x2_ASAP7_75t_L g7818 ( 
.A(n_7754),
.B(n_7763),
.Y(n_7818)
);

OR2x2_ASAP7_75t_L g7819 ( 
.A(n_7754),
.B(n_7474),
.Y(n_7819)
);

INVx2_ASAP7_75t_L g7820 ( 
.A(n_7677),
.Y(n_7820)
);

INVx2_ASAP7_75t_L g7821 ( 
.A(n_7677),
.Y(n_7821)
);

INVx2_ASAP7_75t_L g7822 ( 
.A(n_7719),
.Y(n_7822)
);

INVx1_ASAP7_75t_L g7823 ( 
.A(n_7732),
.Y(n_7823)
);

INVx1_ASAP7_75t_L g7824 ( 
.A(n_7629),
.Y(n_7824)
);

AND2x2_ASAP7_75t_L g7825 ( 
.A(n_7813),
.B(n_7514),
.Y(n_7825)
);

INVx2_ASAP7_75t_L g7826 ( 
.A(n_7719),
.Y(n_7826)
);

INVxp67_ASAP7_75t_SL g7827 ( 
.A(n_7629),
.Y(n_7827)
);

NAND2xp5_ASAP7_75t_L g7828 ( 
.A(n_7634),
.B(n_7585),
.Y(n_7828)
);

AND2x2_ASAP7_75t_L g7829 ( 
.A(n_7807),
.B(n_7518),
.Y(n_7829)
);

NAND2xp5_ASAP7_75t_L g7830 ( 
.A(n_7634),
.B(n_7569),
.Y(n_7830)
);

NAND2xp5_ASAP7_75t_L g7831 ( 
.A(n_7712),
.B(n_7574),
.Y(n_7831)
);

INVx2_ASAP7_75t_L g7832 ( 
.A(n_7703),
.Y(n_7832)
);

NAND2xp5_ASAP7_75t_L g7833 ( 
.A(n_7608),
.B(n_7598),
.Y(n_7833)
);

NOR2xp33_ASAP7_75t_SL g7834 ( 
.A(n_7780),
.B(n_7473),
.Y(n_7834)
);

AND2x2_ASAP7_75t_L g7835 ( 
.A(n_7641),
.B(n_7520),
.Y(n_7835)
);

INVx1_ASAP7_75t_L g7836 ( 
.A(n_7607),
.Y(n_7836)
);

INVx1_ASAP7_75t_L g7837 ( 
.A(n_7618),
.Y(n_7837)
);

BUFx2_ASAP7_75t_L g7838 ( 
.A(n_7690),
.Y(n_7838)
);

OR2x2_ASAP7_75t_L g7839 ( 
.A(n_7763),
.B(n_7467),
.Y(n_7839)
);

INVx1_ASAP7_75t_L g7840 ( 
.A(n_7644),
.Y(n_7840)
);

OR2x2_ASAP7_75t_L g7841 ( 
.A(n_7770),
.B(n_7464),
.Y(n_7841)
);

OR2x2_ASAP7_75t_L g7842 ( 
.A(n_7770),
.B(n_7598),
.Y(n_7842)
);

INVx1_ASAP7_75t_SL g7843 ( 
.A(n_7661),
.Y(n_7843)
);

AND2x2_ASAP7_75t_L g7844 ( 
.A(n_7806),
.B(n_7522),
.Y(n_7844)
);

NAND2xp5_ASAP7_75t_L g7845 ( 
.A(n_7652),
.B(n_7642),
.Y(n_7845)
);

OR2x2_ASAP7_75t_L g7846 ( 
.A(n_7752),
.B(n_7600),
.Y(n_7846)
);

INVx2_ASAP7_75t_L g7847 ( 
.A(n_7703),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_7673),
.Y(n_7848)
);

NAND2xp5_ASAP7_75t_SL g7849 ( 
.A(n_7690),
.B(n_7413),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_7710),
.Y(n_7850)
);

INVx2_ASAP7_75t_L g7851 ( 
.A(n_7731),
.Y(n_7851)
);

INVx1_ASAP7_75t_L g7852 ( 
.A(n_7713),
.Y(n_7852)
);

OAI21xp5_ASAP7_75t_L g7853 ( 
.A1(n_7670),
.A2(n_7593),
.B(n_7392),
.Y(n_7853)
);

OR2x2_ASAP7_75t_L g7854 ( 
.A(n_7752),
.B(n_7600),
.Y(n_7854)
);

INVx2_ASAP7_75t_L g7855 ( 
.A(n_7731),
.Y(n_7855)
);

NAND2xp5_ASAP7_75t_L g7856 ( 
.A(n_7652),
.B(n_7473),
.Y(n_7856)
);

OR2x2_ASAP7_75t_L g7857 ( 
.A(n_7687),
.B(n_7476),
.Y(n_7857)
);

INVx1_ASAP7_75t_L g7858 ( 
.A(n_7714),
.Y(n_7858)
);

NAND2xp5_ASAP7_75t_L g7859 ( 
.A(n_7647),
.B(n_7544),
.Y(n_7859)
);

NAND2x1p5_ASAP7_75t_L g7860 ( 
.A(n_7669),
.B(n_7553),
.Y(n_7860)
);

INVx1_ASAP7_75t_L g7861 ( 
.A(n_7717),
.Y(n_7861)
);

INVx1_ASAP7_75t_SL g7862 ( 
.A(n_7670),
.Y(n_7862)
);

NAND2xp5_ASAP7_75t_L g7863 ( 
.A(n_7642),
.B(n_7519),
.Y(n_7863)
);

NAND2xp5_ASAP7_75t_L g7864 ( 
.A(n_7721),
.B(n_7519),
.Y(n_7864)
);

INVx1_ASAP7_75t_L g7865 ( 
.A(n_7726),
.Y(n_7865)
);

AND2x2_ASAP7_75t_L g7866 ( 
.A(n_7631),
.B(n_7649),
.Y(n_7866)
);

AND2x2_ASAP7_75t_SL g7867 ( 
.A(n_7741),
.B(n_7587),
.Y(n_7867)
);

BUFx2_ASAP7_75t_L g7868 ( 
.A(n_7790),
.Y(n_7868)
);

AND3x2_ASAP7_75t_L g7869 ( 
.A(n_7630),
.B(n_7392),
.C(n_7443),
.Y(n_7869)
);

INVx1_ASAP7_75t_L g7870 ( 
.A(n_7742),
.Y(n_7870)
);

AND2x2_ASAP7_75t_L g7871 ( 
.A(n_7805),
.B(n_7504),
.Y(n_7871)
);

AND2x2_ASAP7_75t_L g7872 ( 
.A(n_7633),
.B(n_7509),
.Y(n_7872)
);

AND2x2_ASAP7_75t_L g7873 ( 
.A(n_7635),
.B(n_7511),
.Y(n_7873)
);

INVx2_ASAP7_75t_SL g7874 ( 
.A(n_7790),
.Y(n_7874)
);

INVx1_ASAP7_75t_L g7875 ( 
.A(n_7762),
.Y(n_7875)
);

NAND2xp5_ASAP7_75t_L g7876 ( 
.A(n_7721),
.B(n_7508),
.Y(n_7876)
);

OR2x2_ASAP7_75t_L g7877 ( 
.A(n_7687),
.B(n_7492),
.Y(n_7877)
);

INVx1_ASAP7_75t_L g7878 ( 
.A(n_7810),
.Y(n_7878)
);

NOR2xp33_ASAP7_75t_L g7879 ( 
.A(n_7686),
.B(n_7486),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_7622),
.Y(n_7880)
);

AND2x2_ASAP7_75t_L g7881 ( 
.A(n_7638),
.B(n_7513),
.Y(n_7881)
);

AND2x2_ASAP7_75t_L g7882 ( 
.A(n_7666),
.B(n_7534),
.Y(n_7882)
);

INVxp67_ASAP7_75t_L g7883 ( 
.A(n_7757),
.Y(n_7883)
);

INVx2_ASAP7_75t_L g7884 ( 
.A(n_7700),
.Y(n_7884)
);

AND2x4_ASAP7_75t_L g7885 ( 
.A(n_7700),
.B(n_7561),
.Y(n_7885)
);

NAND2xp5_ASAP7_75t_L g7886 ( 
.A(n_7718),
.B(n_7508),
.Y(n_7886)
);

AND2x2_ASAP7_75t_L g7887 ( 
.A(n_7688),
.B(n_7538),
.Y(n_7887)
);

NAND2xp5_ASAP7_75t_L g7888 ( 
.A(n_7718),
.B(n_7492),
.Y(n_7888)
);

INVx2_ASAP7_75t_L g7889 ( 
.A(n_7704),
.Y(n_7889)
);

NOR2x1p5_ASAP7_75t_L g7890 ( 
.A(n_7780),
.B(n_7487),
.Y(n_7890)
);

AND2x2_ASAP7_75t_L g7891 ( 
.A(n_7689),
.B(n_7497),
.Y(n_7891)
);

AND2x2_ASAP7_75t_L g7892 ( 
.A(n_7628),
.B(n_7502),
.Y(n_7892)
);

INVx1_ASAP7_75t_L g7893 ( 
.A(n_7623),
.Y(n_7893)
);

AND2x2_ASAP7_75t_L g7894 ( 
.A(n_7615),
.B(n_7507),
.Y(n_7894)
);

NAND2xp5_ASAP7_75t_L g7895 ( 
.A(n_7624),
.B(n_7503),
.Y(n_7895)
);

NAND4xp25_ASAP7_75t_L g7896 ( 
.A(n_7796),
.B(n_7435),
.C(n_7495),
.D(n_7595),
.Y(n_7896)
);

AND2x4_ASAP7_75t_L g7897 ( 
.A(n_7704),
.B(n_7503),
.Y(n_7897)
);

INVx1_ASAP7_75t_L g7898 ( 
.A(n_7632),
.Y(n_7898)
);

NAND2xp33_ASAP7_75t_SL g7899 ( 
.A(n_7722),
.B(n_7488),
.Y(n_7899)
);

OR2x2_ASAP7_75t_L g7900 ( 
.A(n_7723),
.B(n_7506),
.Y(n_7900)
);

INVx1_ASAP7_75t_L g7901 ( 
.A(n_7667),
.Y(n_7901)
);

AND2x2_ASAP7_75t_L g7902 ( 
.A(n_7651),
.B(n_7539),
.Y(n_7902)
);

AND2x2_ASAP7_75t_L g7903 ( 
.A(n_7655),
.B(n_7531),
.Y(n_7903)
);

INVx1_ASAP7_75t_L g7904 ( 
.A(n_7636),
.Y(n_7904)
);

INVx1_ASAP7_75t_L g7905 ( 
.A(n_7639),
.Y(n_7905)
);

INVx1_ASAP7_75t_L g7906 ( 
.A(n_7611),
.Y(n_7906)
);

AND2x2_ASAP7_75t_L g7907 ( 
.A(n_7643),
.B(n_7531),
.Y(n_7907)
);

AND2x2_ASAP7_75t_L g7908 ( 
.A(n_7691),
.B(n_7594),
.Y(n_7908)
);

OR2x2_ASAP7_75t_L g7909 ( 
.A(n_7723),
.B(n_7506),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_7611),
.Y(n_7910)
);

AND2x2_ASAP7_75t_L g7911 ( 
.A(n_7695),
.B(n_7594),
.Y(n_7911)
);

INVx1_ASAP7_75t_L g7912 ( 
.A(n_7681),
.Y(n_7912)
);

AND2x2_ASAP7_75t_L g7913 ( 
.A(n_7662),
.B(n_7599),
.Y(n_7913)
);

NAND2xp5_ASAP7_75t_L g7914 ( 
.A(n_7796),
.B(n_7601),
.Y(n_7914)
);

NAND2xp5_ASAP7_75t_L g7915 ( 
.A(n_7609),
.B(n_7601),
.Y(n_7915)
);

AND2x2_ASAP7_75t_L g7916 ( 
.A(n_7776),
.B(n_7599),
.Y(n_7916)
);

OR2x2_ASAP7_75t_L g7917 ( 
.A(n_7620),
.B(n_7510),
.Y(n_7917)
);

INVx1_ASAP7_75t_L g7918 ( 
.A(n_7725),
.Y(n_7918)
);

AND2x2_ASAP7_75t_L g7919 ( 
.A(n_7614),
.B(n_7603),
.Y(n_7919)
);

NAND2xp5_ASAP7_75t_L g7920 ( 
.A(n_7610),
.B(n_7604),
.Y(n_7920)
);

AND3x1_ASAP7_75t_L g7921 ( 
.A(n_7674),
.B(n_7435),
.C(n_7393),
.Y(n_7921)
);

AND2x2_ASAP7_75t_L g7922 ( 
.A(n_7706),
.B(n_7603),
.Y(n_7922)
);

OR2x2_ASAP7_75t_L g7923 ( 
.A(n_7637),
.B(n_7575),
.Y(n_7923)
);

AND2x2_ASAP7_75t_L g7924 ( 
.A(n_7617),
.B(n_7380),
.Y(n_7924)
);

INVx1_ASAP7_75t_L g7925 ( 
.A(n_7626),
.Y(n_7925)
);

OR2x2_ASAP7_75t_L g7926 ( 
.A(n_7727),
.B(n_7380),
.Y(n_7926)
);

HB1xp67_ASAP7_75t_L g7927 ( 
.A(n_7626),
.Y(n_7927)
);

INVx1_ASAP7_75t_L g7928 ( 
.A(n_7693),
.Y(n_7928)
);

AND2x2_ASAP7_75t_L g7929 ( 
.A(n_7761),
.B(n_7779),
.Y(n_7929)
);

NAND2xp5_ASAP7_75t_L g7930 ( 
.A(n_7613),
.B(n_7604),
.Y(n_7930)
);

NAND2xp5_ASAP7_75t_L g7931 ( 
.A(n_7619),
.B(n_7605),
.Y(n_7931)
);

NAND2xp5_ASAP7_75t_L g7932 ( 
.A(n_7759),
.B(n_7605),
.Y(n_7932)
);

NAND2xp5_ASAP7_75t_L g7933 ( 
.A(n_7760),
.B(n_7516),
.Y(n_7933)
);

AND2x4_ASAP7_75t_L g7934 ( 
.A(n_7612),
.B(n_7393),
.Y(n_7934)
);

AND2x2_ASAP7_75t_L g7935 ( 
.A(n_7734),
.B(n_7410),
.Y(n_7935)
);

NAND2xp5_ASAP7_75t_L g7936 ( 
.A(n_7696),
.B(n_7565),
.Y(n_7936)
);

NAND2xp5_ASAP7_75t_L g7937 ( 
.A(n_7680),
.B(n_7565),
.Y(n_7937)
);

INVx1_ASAP7_75t_L g7938 ( 
.A(n_7727),
.Y(n_7938)
);

BUFx2_ASAP7_75t_L g7939 ( 
.A(n_7692),
.Y(n_7939)
);

AND2x2_ASAP7_75t_L g7940 ( 
.A(n_7737),
.B(n_7410),
.Y(n_7940)
);

OR2x2_ASAP7_75t_L g7941 ( 
.A(n_7708),
.B(n_7411),
.Y(n_7941)
);

INVx1_ASAP7_75t_L g7942 ( 
.A(n_7684),
.Y(n_7942)
);

OR2x2_ASAP7_75t_L g7943 ( 
.A(n_7708),
.B(n_7411),
.Y(n_7943)
);

AND2x2_ASAP7_75t_L g7944 ( 
.A(n_7774),
.B(n_7564),
.Y(n_7944)
);

OR2x2_ASAP7_75t_L g7945 ( 
.A(n_7684),
.B(n_7596),
.Y(n_7945)
);

AND2x2_ASAP7_75t_L g7946 ( 
.A(n_7787),
.B(n_7443),
.Y(n_7946)
);

AND2x2_ASAP7_75t_L g7947 ( 
.A(n_7788),
.B(n_7447),
.Y(n_7947)
);

NAND2xp5_ASAP7_75t_L g7948 ( 
.A(n_7798),
.B(n_7571),
.Y(n_7948)
);

AOI22xp33_ASAP7_75t_L g7949 ( 
.A1(n_7674),
.A2(n_6562),
.B1(n_6811),
.B2(n_6707),
.Y(n_7949)
);

INVxp67_ASAP7_75t_L g7950 ( 
.A(n_7736),
.Y(n_7950)
);

INVx1_ASAP7_75t_L g7951 ( 
.A(n_7743),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_7646),
.Y(n_7952)
);

INVx3_ASAP7_75t_L g7953 ( 
.A(n_7765),
.Y(n_7953)
);

INVx1_ASAP7_75t_L g7954 ( 
.A(n_7797),
.Y(n_7954)
);

INVx2_ASAP7_75t_L g7955 ( 
.A(n_7765),
.Y(n_7955)
);

OR2x2_ASAP7_75t_L g7956 ( 
.A(n_7808),
.B(n_7590),
.Y(n_7956)
);

INVx1_ASAP7_75t_L g7957 ( 
.A(n_7799),
.Y(n_7957)
);

INVx1_ASAP7_75t_L g7958 ( 
.A(n_7809),
.Y(n_7958)
);

OAI21xp33_ASAP7_75t_L g7959 ( 
.A1(n_7682),
.A2(n_7493),
.B(n_7553),
.Y(n_7959)
);

AND2x2_ASAP7_75t_L g7960 ( 
.A(n_7793),
.B(n_7447),
.Y(n_7960)
);

BUFx2_ASAP7_75t_L g7961 ( 
.A(n_7692),
.Y(n_7961)
);

INVx1_ASAP7_75t_L g7962 ( 
.A(n_7716),
.Y(n_7962)
);

OAI21xp5_ASAP7_75t_L g7963 ( 
.A1(n_7682),
.A2(n_7470),
.B(n_7468),
.Y(n_7963)
);

AND2x2_ASAP7_75t_L g7964 ( 
.A(n_7800),
.B(n_7558),
.Y(n_7964)
);

INVx2_ASAP7_75t_L g7965 ( 
.A(n_7744),
.Y(n_7965)
);

INVx2_ASAP7_75t_L g7966 ( 
.A(n_7744),
.Y(n_7966)
);

INVxp67_ASAP7_75t_SL g7967 ( 
.A(n_7625),
.Y(n_7967)
);

AND2x2_ASAP7_75t_L g7968 ( 
.A(n_7803),
.B(n_7558),
.Y(n_7968)
);

AND2x2_ASAP7_75t_L g7969 ( 
.A(n_7748),
.B(n_7456),
.Y(n_7969)
);

INVx1_ASAP7_75t_L g7970 ( 
.A(n_7648),
.Y(n_7970)
);

AND2x2_ASAP7_75t_L g7971 ( 
.A(n_7705),
.B(n_7456),
.Y(n_7971)
);

INVx1_ASAP7_75t_L g7972 ( 
.A(n_7656),
.Y(n_7972)
);

INVx1_ASAP7_75t_L g7973 ( 
.A(n_7657),
.Y(n_7973)
);

AND2x2_ASAP7_75t_L g7974 ( 
.A(n_7789),
.B(n_7517),
.Y(n_7974)
);

NOR2xp33_ASAP7_75t_L g7975 ( 
.A(n_7659),
.B(n_7466),
.Y(n_7975)
);

AND2x2_ASAP7_75t_L g7976 ( 
.A(n_7791),
.B(n_7523),
.Y(n_7976)
);

AND2x2_ASAP7_75t_L g7977 ( 
.A(n_7794),
.B(n_7524),
.Y(n_7977)
);

OR2x2_ASAP7_75t_L g7978 ( 
.A(n_7808),
.B(n_7533),
.Y(n_7978)
);

INVxp33_ASAP7_75t_L g7979 ( 
.A(n_7786),
.Y(n_7979)
);

OR2x2_ASAP7_75t_L g7980 ( 
.A(n_7729),
.B(n_7298),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_L g7981 ( 
.A(n_7798),
.B(n_7571),
.Y(n_7981)
);

OR2x2_ASAP7_75t_L g7982 ( 
.A(n_7699),
.B(n_7307),
.Y(n_7982)
);

NAND2xp5_ASAP7_75t_L g7983 ( 
.A(n_7645),
.B(n_7573),
.Y(n_7983)
);

INVx1_ASAP7_75t_L g7984 ( 
.A(n_7650),
.Y(n_7984)
);

INVx2_ASAP7_75t_L g7985 ( 
.A(n_7621),
.Y(n_7985)
);

NAND2xp5_ASAP7_75t_L g7986 ( 
.A(n_7658),
.B(n_7573),
.Y(n_7986)
);

HB1xp67_ASAP7_75t_L g7987 ( 
.A(n_7711),
.Y(n_7987)
);

OR2x2_ASAP7_75t_L g7988 ( 
.A(n_7785),
.B(n_7307),
.Y(n_7988)
);

AND2x2_ASAP7_75t_L g7989 ( 
.A(n_7768),
.B(n_7589),
.Y(n_7989)
);

AND2x2_ASAP7_75t_L g7990 ( 
.A(n_7778),
.B(n_7589),
.Y(n_7990)
);

AND2x2_ASAP7_75t_L g7991 ( 
.A(n_7795),
.B(n_7597),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_7663),
.Y(n_7992)
);

INVx1_ASAP7_75t_L g7993 ( 
.A(n_7730),
.Y(n_7993)
);

OR2x2_ASAP7_75t_L g7994 ( 
.A(n_7668),
.B(n_7323),
.Y(n_7994)
);

OR2x2_ASAP7_75t_L g7995 ( 
.A(n_7660),
.B(n_7323),
.Y(n_7995)
);

INVx1_ASAP7_75t_SL g7996 ( 
.A(n_7616),
.Y(n_7996)
);

INVx2_ASAP7_75t_L g7997 ( 
.A(n_7701),
.Y(n_7997)
);

INVx1_ASAP7_75t_L g7998 ( 
.A(n_7730),
.Y(n_7998)
);

AND2x2_ASAP7_75t_L g7999 ( 
.A(n_7749),
.B(n_7597),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_7735),
.Y(n_8000)
);

AND2x2_ASAP7_75t_L g8001 ( 
.A(n_7747),
.B(n_7528),
.Y(n_8001)
);

OR2x2_ASAP7_75t_L g8002 ( 
.A(n_7764),
.B(n_7276),
.Y(n_8002)
);

NAND2xp5_ASAP7_75t_L g8003 ( 
.A(n_7755),
.B(n_7528),
.Y(n_8003)
);

HB1xp67_ASAP7_75t_L g8004 ( 
.A(n_7625),
.Y(n_8004)
);

INVx1_ASAP7_75t_L g8005 ( 
.A(n_7735),
.Y(n_8005)
);

AND2x2_ASAP7_75t_L g8006 ( 
.A(n_7659),
.B(n_7528),
.Y(n_8006)
);

INVx1_ASAP7_75t_L g8007 ( 
.A(n_7927),
.Y(n_8007)
);

OAI211xp5_ASAP7_75t_L g8008 ( 
.A1(n_7949),
.A2(n_7616),
.B(n_7640),
.C(n_7654),
.Y(n_8008)
);

INVx2_ASAP7_75t_L g8009 ( 
.A(n_7885),
.Y(n_8009)
);

AND2x2_ASAP7_75t_L g8010 ( 
.A(n_7913),
.B(n_7685),
.Y(n_8010)
);

NAND2xp5_ASAP7_75t_SL g8011 ( 
.A(n_7885),
.B(n_7529),
.Y(n_8011)
);

INVx1_ASAP7_75t_L g8012 ( 
.A(n_7868),
.Y(n_8012)
);

INVx1_ASAP7_75t_L g8013 ( 
.A(n_7838),
.Y(n_8013)
);

OAI22xp33_ASAP7_75t_SL g8014 ( 
.A1(n_7864),
.A2(n_7627),
.B1(n_7001),
.B2(n_7683),
.Y(n_8014)
);

NAND2xp5_ASAP7_75t_L g8015 ( 
.A(n_7897),
.B(n_7529),
.Y(n_8015)
);

INVx1_ASAP7_75t_L g8016 ( 
.A(n_7833),
.Y(n_8016)
);

OR2x2_ASAP7_75t_L g8017 ( 
.A(n_7906),
.B(n_7707),
.Y(n_8017)
);

AND2x4_ASAP7_75t_L g8018 ( 
.A(n_7897),
.B(n_7874),
.Y(n_8018)
);

INVx1_ASAP7_75t_L g8019 ( 
.A(n_7833),
.Y(n_8019)
);

AND2x2_ASAP7_75t_L g8020 ( 
.A(n_7892),
.B(n_7685),
.Y(n_8020)
);

NAND2xp5_ASAP7_75t_L g8021 ( 
.A(n_7919),
.B(n_7529),
.Y(n_8021)
);

OR2x2_ASAP7_75t_L g8022 ( 
.A(n_7910),
.B(n_7720),
.Y(n_8022)
);

NAND2xp5_ASAP7_75t_L g8023 ( 
.A(n_7922),
.B(n_7756),
.Y(n_8023)
);

INVx1_ASAP7_75t_L g8024 ( 
.A(n_7827),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_7818),
.Y(n_8025)
);

OR2x2_ASAP7_75t_L g8026 ( 
.A(n_7843),
.B(n_7802),
.Y(n_8026)
);

AND2x2_ASAP7_75t_L g8027 ( 
.A(n_7907),
.B(n_7758),
.Y(n_8027)
);

OR2x2_ASAP7_75t_L g8028 ( 
.A(n_7843),
.B(n_7802),
.Y(n_8028)
);

AND3x2_ASAP7_75t_L g8029 ( 
.A(n_7834),
.B(n_7683),
.C(n_7801),
.Y(n_8029)
);

INVxp67_ASAP7_75t_L g8030 ( 
.A(n_7834),
.Y(n_8030)
);

OR2x2_ASAP7_75t_L g8031 ( 
.A(n_7846),
.B(n_7772),
.Y(n_8031)
);

AND2x2_ASAP7_75t_L g8032 ( 
.A(n_7902),
.B(n_7766),
.Y(n_8032)
);

NAND2xp5_ASAP7_75t_L g8033 ( 
.A(n_7866),
.B(n_7664),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_7924),
.Y(n_8034)
);

INVx2_ASAP7_75t_SL g8035 ( 
.A(n_8001),
.Y(n_8035)
);

HB1xp67_ASAP7_75t_L g8036 ( 
.A(n_7860),
.Y(n_8036)
);

NAND2xp5_ASAP7_75t_L g8037 ( 
.A(n_7872),
.B(n_7671),
.Y(n_8037)
);

INVx1_ASAP7_75t_L g8038 ( 
.A(n_7941),
.Y(n_8038)
);

AND2x2_ASAP7_75t_L g8039 ( 
.A(n_7873),
.B(n_7881),
.Y(n_8039)
);

INVx1_ASAP7_75t_L g8040 ( 
.A(n_7943),
.Y(n_8040)
);

INVxp33_ASAP7_75t_L g8041 ( 
.A(n_7916),
.Y(n_8041)
);

NAND2xp5_ASAP7_75t_L g8042 ( 
.A(n_7894),
.B(n_7672),
.Y(n_8042)
);

INVx2_ASAP7_75t_L g8043 ( 
.A(n_7860),
.Y(n_8043)
);

AND2x2_ASAP7_75t_L g8044 ( 
.A(n_7835),
.B(n_7694),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_7925),
.Y(n_8045)
);

AND2x2_ASAP7_75t_L g8046 ( 
.A(n_7816),
.B(n_7698),
.Y(n_8046)
);

AND2x2_ASAP7_75t_L g8047 ( 
.A(n_7903),
.B(n_7709),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_8006),
.Y(n_8048)
);

OR2x2_ASAP7_75t_L g8049 ( 
.A(n_7854),
.B(n_7653),
.Y(n_8049)
);

AND2x2_ASAP7_75t_L g8050 ( 
.A(n_7891),
.B(n_7715),
.Y(n_8050)
);

AND2x2_ASAP7_75t_L g8051 ( 
.A(n_7815),
.B(n_7724),
.Y(n_8051)
);

INVx1_ASAP7_75t_L g8052 ( 
.A(n_7820),
.Y(n_8052)
);

AND2x2_ASAP7_75t_L g8053 ( 
.A(n_7871),
.B(n_7728),
.Y(n_8053)
);

INVx1_ASAP7_75t_L g8054 ( 
.A(n_7821),
.Y(n_8054)
);

INVx1_ASAP7_75t_L g8055 ( 
.A(n_7908),
.Y(n_8055)
);

OAI21xp5_ASAP7_75t_L g8056 ( 
.A1(n_7864),
.A2(n_7640),
.B(n_7627),
.Y(n_8056)
);

INVx2_ASAP7_75t_L g8057 ( 
.A(n_7869),
.Y(n_8057)
);

INVx1_ASAP7_75t_L g8058 ( 
.A(n_7911),
.Y(n_8058)
);

AOI22xp5_ASAP7_75t_L g8059 ( 
.A1(n_7876),
.A2(n_7921),
.B1(n_7899),
.B2(n_7867),
.Y(n_8059)
);

OR2x2_ASAP7_75t_L g8060 ( 
.A(n_7828),
.B(n_7777),
.Y(n_8060)
);

AOI22xp5_ASAP7_75t_L g8061 ( 
.A1(n_7876),
.A2(n_7665),
.B1(n_7654),
.B2(n_7801),
.Y(n_8061)
);

INVx1_ASAP7_75t_L g8062 ( 
.A(n_7934),
.Y(n_8062)
);

NAND2xp5_ASAP7_75t_L g8063 ( 
.A(n_7934),
.B(n_7676),
.Y(n_8063)
);

INVx2_ASAP7_75t_SL g8064 ( 
.A(n_7842),
.Y(n_8064)
);

NOR2x1_ASAP7_75t_L g8065 ( 
.A(n_7948),
.B(n_7471),
.Y(n_8065)
);

INVx1_ASAP7_75t_L g8066 ( 
.A(n_7888),
.Y(n_8066)
);

INVx2_ASAP7_75t_L g8067 ( 
.A(n_7887),
.Y(n_8067)
);

INVx2_ASAP7_75t_L g8068 ( 
.A(n_7844),
.Y(n_8068)
);

INVx3_ASAP7_75t_L g8069 ( 
.A(n_7953),
.Y(n_8069)
);

INVx1_ASAP7_75t_L g8070 ( 
.A(n_7888),
.Y(n_8070)
);

INVx2_ASAP7_75t_SL g8071 ( 
.A(n_7953),
.Y(n_8071)
);

INVx1_ASAP7_75t_L g8072 ( 
.A(n_7964),
.Y(n_8072)
);

NAND2xp5_ASAP7_75t_L g8073 ( 
.A(n_7825),
.B(n_7560),
.Y(n_8073)
);

BUFx3_ASAP7_75t_L g8074 ( 
.A(n_7884),
.Y(n_8074)
);

OR2x2_ASAP7_75t_L g8075 ( 
.A(n_7828),
.B(n_7781),
.Y(n_8075)
);

NAND2xp5_ASAP7_75t_L g8076 ( 
.A(n_7829),
.B(n_7560),
.Y(n_8076)
);

NAND2xp5_ASAP7_75t_L g8077 ( 
.A(n_7837),
.B(n_7562),
.Y(n_8077)
);

INVx1_ASAP7_75t_L g8078 ( 
.A(n_7968),
.Y(n_8078)
);

INVx1_ASAP7_75t_L g8079 ( 
.A(n_7936),
.Y(n_8079)
);

NAND2xp5_ASAP7_75t_L g8080 ( 
.A(n_7882),
.B(n_7832),
.Y(n_8080)
);

O2A1O1Ixp33_ASAP7_75t_L g8081 ( 
.A1(n_7914),
.A2(n_7665),
.B(n_7811),
.C(n_7498),
.Y(n_8081)
);

INVx2_ASAP7_75t_L g8082 ( 
.A(n_7889),
.Y(n_8082)
);

INVx2_ASAP7_75t_L g8083 ( 
.A(n_7877),
.Y(n_8083)
);

INVx2_ASAP7_75t_SL g8084 ( 
.A(n_7847),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_7936),
.Y(n_8085)
);

INVx2_ASAP7_75t_L g8086 ( 
.A(n_7822),
.Y(n_8086)
);

AOI21xp33_ASAP7_75t_L g8087 ( 
.A1(n_7819),
.A2(n_7702),
.B(n_7746),
.Y(n_8087)
);

INVx1_ASAP7_75t_L g8088 ( 
.A(n_7839),
.Y(n_8088)
);

NAND2xp5_ASAP7_75t_L g8089 ( 
.A(n_7826),
.B(n_7562),
.Y(n_8089)
);

INVx1_ASAP7_75t_L g8090 ( 
.A(n_7969),
.Y(n_8090)
);

INVx1_ASAP7_75t_L g8091 ( 
.A(n_8003),
.Y(n_8091)
);

NAND2xp5_ASAP7_75t_L g8092 ( 
.A(n_7946),
.B(n_7491),
.Y(n_8092)
);

NOR2xp33_ASAP7_75t_L g8093 ( 
.A(n_7896),
.B(n_7784),
.Y(n_8093)
);

OR2x2_ASAP7_75t_L g8094 ( 
.A(n_7830),
.B(n_7804),
.Y(n_8094)
);

A2O1A1Ixp33_ASAP7_75t_L g8095 ( 
.A1(n_7914),
.A2(n_6917),
.B(n_7811),
.C(n_6861),
.Y(n_8095)
);

AND2x2_ASAP7_75t_L g8096 ( 
.A(n_7935),
.B(n_7812),
.Y(n_8096)
);

AND2x2_ASAP7_75t_L g8097 ( 
.A(n_7940),
.B(n_7814),
.Y(n_8097)
);

NAND2x2_ASAP7_75t_L g8098 ( 
.A(n_7890),
.B(n_7675),
.Y(n_8098)
);

INVx2_ASAP7_75t_L g8099 ( 
.A(n_7900),
.Y(n_8099)
);

NAND2xp5_ASAP7_75t_L g8100 ( 
.A(n_7947),
.B(n_7536),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_7960),
.Y(n_8101)
);

INVx1_ASAP7_75t_L g8102 ( 
.A(n_7909),
.Y(n_8102)
);

INVx2_ASAP7_75t_L g8103 ( 
.A(n_7926),
.Y(n_8103)
);

INVx1_ASAP7_75t_L g8104 ( 
.A(n_7999),
.Y(n_8104)
);

NAND2xp5_ASAP7_75t_L g8105 ( 
.A(n_7928),
.B(n_7543),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_7830),
.Y(n_8106)
);

AND2x4_ASAP7_75t_SL g8107 ( 
.A(n_7997),
.B(n_7457),
.Y(n_8107)
);

OAI21xp33_ASAP7_75t_L g8108 ( 
.A1(n_7896),
.A2(n_7697),
.B(n_7460),
.Y(n_8108)
);

AND2x2_ASAP7_75t_L g8109 ( 
.A(n_7971),
.B(n_7458),
.Y(n_8109)
);

AND2x2_ASAP7_75t_L g8110 ( 
.A(n_7929),
.B(n_7944),
.Y(n_8110)
);

BUFx2_ASAP7_75t_L g8111 ( 
.A(n_7824),
.Y(n_8111)
);

INVx1_ASAP7_75t_L g8112 ( 
.A(n_7937),
.Y(n_8112)
);

INVx1_ASAP7_75t_L g8113 ( 
.A(n_7937),
.Y(n_8113)
);

AND2x2_ASAP7_75t_L g8114 ( 
.A(n_7962),
.B(n_7457),
.Y(n_8114)
);

AND2x2_ASAP7_75t_L g8115 ( 
.A(n_7912),
.B(n_7483),
.Y(n_8115)
);

OR2x2_ASAP7_75t_L g8116 ( 
.A(n_7831),
.B(n_7276),
.Y(n_8116)
);

AND2x4_ASAP7_75t_L g8117 ( 
.A(n_7851),
.B(n_7483),
.Y(n_8117)
);

INVx1_ASAP7_75t_SL g8118 ( 
.A(n_7996),
.Y(n_8118)
);

INVx1_ASAP7_75t_L g8119 ( 
.A(n_7859),
.Y(n_8119)
);

OAI21xp33_ASAP7_75t_L g8120 ( 
.A1(n_7831),
.A2(n_7290),
.B(n_7285),
.Y(n_8120)
);

AND2x2_ASAP7_75t_SL g8121 ( 
.A(n_7921),
.B(n_7857),
.Y(n_8121)
);

OR2x2_ASAP7_75t_L g8122 ( 
.A(n_7886),
.B(n_7285),
.Y(n_8122)
);

INVx1_ASAP7_75t_L g8123 ( 
.A(n_7895),
.Y(n_8123)
);

NAND2xp5_ASAP7_75t_L g8124 ( 
.A(n_7918),
.B(n_7767),
.Y(n_8124)
);

OR2x2_ASAP7_75t_L g8125 ( 
.A(n_7886),
.B(n_7290),
.Y(n_8125)
);

NAND2xp5_ASAP7_75t_L g8126 ( 
.A(n_7985),
.B(n_7769),
.Y(n_8126)
);

AND2x2_ASAP7_75t_L g8127 ( 
.A(n_7951),
.B(n_7771),
.Y(n_8127)
);

AOI22xp5_ASAP7_75t_L g8128 ( 
.A1(n_7862),
.A2(n_7023),
.B1(n_7001),
.B2(n_7773),
.Y(n_8128)
);

INVx1_ASAP7_75t_L g8129 ( 
.A(n_7895),
.Y(n_8129)
);

AND2x2_ASAP7_75t_L g8130 ( 
.A(n_7952),
.B(n_7775),
.Y(n_8130)
);

OR2x2_ASAP7_75t_L g8131 ( 
.A(n_7923),
.B(n_7247),
.Y(n_8131)
);

AND2x2_ASAP7_75t_L g8132 ( 
.A(n_7970),
.B(n_7783),
.Y(n_8132)
);

OR2x2_ASAP7_75t_L g8133 ( 
.A(n_7945),
.B(n_7247),
.Y(n_8133)
);

INVx1_ASAP7_75t_L g8134 ( 
.A(n_7817),
.Y(n_8134)
);

NAND4xp25_ASAP7_75t_L g8135 ( 
.A(n_7879),
.B(n_7738),
.C(n_7739),
.D(n_7733),
.Y(n_8135)
);

OAI21xp33_ASAP7_75t_L g8136 ( 
.A1(n_7863),
.A2(n_7792),
.B(n_7782),
.Y(n_8136)
);

NAND2xp5_ASAP7_75t_L g8137 ( 
.A(n_7939),
.B(n_7546),
.Y(n_8137)
);

INVx1_ASAP7_75t_L g8138 ( 
.A(n_7823),
.Y(n_8138)
);

NAND2x2_ASAP7_75t_L g8139 ( 
.A(n_7841),
.B(n_7782),
.Y(n_8139)
);

OAI22xp33_ASAP7_75t_SL g8140 ( 
.A1(n_7948),
.A2(n_7001),
.B1(n_7023),
.B2(n_7479),
.Y(n_8140)
);

INVx1_ASAP7_75t_L g8141 ( 
.A(n_7856),
.Y(n_8141)
);

OAI21xp33_ASAP7_75t_L g8142 ( 
.A1(n_7863),
.A2(n_7792),
.B(n_7023),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7856),
.Y(n_8143)
);

AND2x2_ASAP7_75t_L g8144 ( 
.A(n_7989),
.B(n_7547),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7932),
.Y(n_8145)
);

AND2x2_ASAP7_75t_L g8146 ( 
.A(n_7990),
.B(n_7548),
.Y(n_8146)
);

AND2x2_ASAP7_75t_L g8147 ( 
.A(n_7991),
.B(n_7740),
.Y(n_8147)
);

INVx2_ASAP7_75t_L g8148 ( 
.A(n_7917),
.Y(n_8148)
);

INVx2_ASAP7_75t_L g8149 ( 
.A(n_7961),
.Y(n_8149)
);

INVx3_ASAP7_75t_L g8150 ( 
.A(n_7855),
.Y(n_8150)
);

INVx1_ASAP7_75t_L g8151 ( 
.A(n_7932),
.Y(n_8151)
);

AND2x2_ASAP7_75t_L g8152 ( 
.A(n_7955),
.B(n_7745),
.Y(n_8152)
);

AOI31xp33_ASAP7_75t_L g8153 ( 
.A1(n_7981),
.A2(n_7750),
.A3(n_7679),
.B(n_7678),
.Y(n_8153)
);

AND2x2_ASAP7_75t_L g8154 ( 
.A(n_7974),
.B(n_7572),
.Y(n_8154)
);

INVxp67_ASAP7_75t_SL g8155 ( 
.A(n_7849),
.Y(n_8155)
);

NAND2xp5_ASAP7_75t_L g8156 ( 
.A(n_7836),
.B(n_7576),
.Y(n_8156)
);

INVx1_ASAP7_75t_L g8157 ( 
.A(n_7980),
.Y(n_8157)
);

AOI22xp5_ASAP7_75t_L g8158 ( 
.A1(n_7862),
.A2(n_7023),
.B1(n_6801),
.B2(n_6810),
.Y(n_8158)
);

INVx1_ASAP7_75t_L g8159 ( 
.A(n_7915),
.Y(n_8159)
);

NAND2xp5_ASAP7_75t_L g8160 ( 
.A(n_7987),
.B(n_7602),
.Y(n_8160)
);

AOI21xp33_ASAP7_75t_L g8161 ( 
.A1(n_7981),
.A2(n_7485),
.B(n_7484),
.Y(n_8161)
);

INVx1_ASAP7_75t_L g8162 ( 
.A(n_7915),
.Y(n_8162)
);

INVx2_ASAP7_75t_L g8163 ( 
.A(n_7965),
.Y(n_8163)
);

INVx4_ASAP7_75t_L g8164 ( 
.A(n_7966),
.Y(n_8164)
);

AND2x2_ASAP7_75t_L g8165 ( 
.A(n_7976),
.B(n_7356),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7959),
.B(n_7358),
.Y(n_8166)
);

INVx1_ASAP7_75t_L g8167 ( 
.A(n_8018),
.Y(n_8167)
);

AND2x2_ASAP7_75t_L g8168 ( 
.A(n_8039),
.B(n_7977),
.Y(n_8168)
);

NOR2xp33_ASAP7_75t_SL g8169 ( 
.A(n_8121),
.B(n_7996),
.Y(n_8169)
);

INVx1_ASAP7_75t_L g8170 ( 
.A(n_8018),
.Y(n_8170)
);

INVx1_ASAP7_75t_L g8171 ( 
.A(n_8015),
.Y(n_8171)
);

OAI22xp5_ASAP7_75t_L g8172 ( 
.A1(n_8059),
.A2(n_7883),
.B1(n_7950),
.B2(n_7979),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_8011),
.Y(n_8173)
);

AND2x2_ASAP7_75t_L g8174 ( 
.A(n_8110),
.B(n_7878),
.Y(n_8174)
);

NAND2xp5_ASAP7_75t_L g8175 ( 
.A(n_8012),
.B(n_7959),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_8021),
.Y(n_8176)
);

INVx1_ASAP7_75t_L g8177 ( 
.A(n_8027),
.Y(n_8177)
);

INVx2_ASAP7_75t_L g8178 ( 
.A(n_8029),
.Y(n_8178)
);

OAI21xp33_ASAP7_75t_L g8179 ( 
.A1(n_8059),
.A2(n_8093),
.B(n_8041),
.Y(n_8179)
);

AND2x2_ASAP7_75t_L g8180 ( 
.A(n_8032),
.B(n_7972),
.Y(n_8180)
);

AND2x4_ASAP7_75t_L g8181 ( 
.A(n_8062),
.B(n_7850),
.Y(n_8181)
);

OAI21xp5_ASAP7_75t_L g8182 ( 
.A1(n_8030),
.A2(n_7845),
.B(n_7853),
.Y(n_8182)
);

INVx1_ASAP7_75t_L g8183 ( 
.A(n_8013),
.Y(n_8183)
);

NAND2xp5_ASAP7_75t_L g8184 ( 
.A(n_8069),
.B(n_7840),
.Y(n_8184)
);

NAND2x1_ASAP7_75t_L g8185 ( 
.A(n_8069),
.B(n_7059),
.Y(n_8185)
);

NAND2xp5_ASAP7_75t_L g8186 ( 
.A(n_8035),
.B(n_7848),
.Y(n_8186)
);

NAND2xp5_ASAP7_75t_L g8187 ( 
.A(n_8009),
.B(n_7852),
.Y(n_8187)
);

INVx1_ASAP7_75t_SL g8188 ( 
.A(n_8118),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_8020),
.Y(n_8189)
);

INVx1_ASAP7_75t_SL g8190 ( 
.A(n_8118),
.Y(n_8190)
);

NAND2xp5_ASAP7_75t_L g8191 ( 
.A(n_8107),
.B(n_7858),
.Y(n_8191)
);

NAND2xp5_ASAP7_75t_L g8192 ( 
.A(n_8071),
.B(n_8117),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_8010),
.Y(n_8193)
);

NOR2x1p5_ASAP7_75t_L g8194 ( 
.A(n_8155),
.B(n_7933),
.Y(n_8194)
);

AND2x2_ASAP7_75t_L g8195 ( 
.A(n_8050),
.B(n_7973),
.Y(n_8195)
);

NAND2xp5_ASAP7_75t_L g8196 ( 
.A(n_8117),
.B(n_7861),
.Y(n_8196)
);

AND2x4_ASAP7_75t_L g8197 ( 
.A(n_8064),
.B(n_7865),
.Y(n_8197)
);

OAI21xp5_ASAP7_75t_L g8198 ( 
.A1(n_8056),
.A2(n_7845),
.B(n_7853),
.Y(n_8198)
);

AND2x2_ASAP7_75t_L g8199 ( 
.A(n_8046),
.B(n_7870),
.Y(n_8199)
);

HB1xp67_ASAP7_75t_L g8200 ( 
.A(n_8036),
.Y(n_8200)
);

AND2x4_ASAP7_75t_SL g8201 ( 
.A(n_8148),
.B(n_7901),
.Y(n_8201)
);

NAND3xp33_ASAP7_75t_L g8202 ( 
.A(n_8056),
.B(n_7963),
.C(n_8004),
.Y(n_8202)
);

NAND2xp5_ASAP7_75t_L g8203 ( 
.A(n_8007),
.B(n_7875),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_8047),
.Y(n_8204)
);

INVx1_ASAP7_75t_L g8205 ( 
.A(n_8063),
.Y(n_8205)
);

INVx1_ASAP7_75t_L g8206 ( 
.A(n_8109),
.Y(n_8206)
);

AND2x2_ASAP7_75t_L g8207 ( 
.A(n_8044),
.B(n_7904),
.Y(n_8207)
);

INVx1_ASAP7_75t_L g8208 ( 
.A(n_8073),
.Y(n_8208)
);

AND2x2_ASAP7_75t_L g8209 ( 
.A(n_8053),
.B(n_7905),
.Y(n_8209)
);

NAND2xp5_ASAP7_75t_L g8210 ( 
.A(n_8067),
.B(n_7967),
.Y(n_8210)
);

OR2x2_ASAP7_75t_L g8211 ( 
.A(n_8049),
.B(n_7994),
.Y(n_8211)
);

INVx1_ASAP7_75t_L g8212 ( 
.A(n_8076),
.Y(n_8212)
);

NOR2xp33_ASAP7_75t_L g8213 ( 
.A(n_8074),
.B(n_7988),
.Y(n_8213)
);

HB1xp67_ASAP7_75t_L g8214 ( 
.A(n_8043),
.Y(n_8214)
);

INVx1_ASAP7_75t_L g8215 ( 
.A(n_8051),
.Y(n_8215)
);

BUFx2_ASAP7_75t_L g8216 ( 
.A(n_8164),
.Y(n_8216)
);

NAND2xp5_ASAP7_75t_L g8217 ( 
.A(n_8090),
.B(n_7880),
.Y(n_8217)
);

AND2x2_ASAP7_75t_L g8218 ( 
.A(n_8068),
.B(n_7933),
.Y(n_8218)
);

O2A1O1Ixp33_ASAP7_75t_SL g8219 ( 
.A1(n_8095),
.A2(n_7351),
.B(n_7357),
.C(n_7343),
.Y(n_8219)
);

OR2x2_ASAP7_75t_L g8220 ( 
.A(n_8131),
.B(n_7982),
.Y(n_8220)
);

HB1xp67_ASAP7_75t_L g8221 ( 
.A(n_8065),
.Y(n_8221)
);

OAI22xp5_ASAP7_75t_L g8222 ( 
.A1(n_8098),
.A2(n_7956),
.B1(n_7978),
.B2(n_7079),
.Y(n_8222)
);

INVx1_ASAP7_75t_L g8223 ( 
.A(n_8114),
.Y(n_8223)
);

INVx1_ASAP7_75t_L g8224 ( 
.A(n_8115),
.Y(n_8224)
);

INVx2_ASAP7_75t_L g8225 ( 
.A(n_8017),
.Y(n_8225)
);

INVx1_ASAP7_75t_L g8226 ( 
.A(n_8023),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_8089),
.Y(n_8227)
);

AOI211xp5_ASAP7_75t_L g8228 ( 
.A1(n_8014),
.A2(n_7963),
.B(n_7975),
.C(n_7938),
.Y(n_8228)
);

INVx3_ASAP7_75t_L g8229 ( 
.A(n_8164),
.Y(n_8229)
);

OR2x2_ASAP7_75t_L g8230 ( 
.A(n_8116),
.B(n_7995),
.Y(n_8230)
);

NAND2xp5_ASAP7_75t_L g8231 ( 
.A(n_8038),
.B(n_7893),
.Y(n_8231)
);

NAND2xp5_ASAP7_75t_L g8232 ( 
.A(n_8040),
.B(n_8034),
.Y(n_8232)
);

AND2x2_ASAP7_75t_L g8233 ( 
.A(n_8082),
.B(n_7942),
.Y(n_8233)
);

AOI21xp33_ASAP7_75t_SL g8234 ( 
.A1(n_8153),
.A2(n_7930),
.B(n_7920),
.Y(n_8234)
);

INVx1_ASAP7_75t_L g8235 ( 
.A(n_8026),
.Y(n_8235)
);

AND2x2_ASAP7_75t_L g8236 ( 
.A(n_8086),
.B(n_7984),
.Y(n_8236)
);

A2O1A1Ixp33_ASAP7_75t_L g8237 ( 
.A1(n_8081),
.A2(n_6938),
.B(n_6954),
.C(n_7954),
.Y(n_8237)
);

INVx2_ASAP7_75t_L g8238 ( 
.A(n_8022),
.Y(n_8238)
);

OR2x2_ASAP7_75t_L g8239 ( 
.A(n_8031),
.B(n_8002),
.Y(n_8239)
);

INVx1_ASAP7_75t_L g8240 ( 
.A(n_8028),
.Y(n_8240)
);

AOI21xp33_ASAP7_75t_SL g8241 ( 
.A1(n_8153),
.A2(n_7930),
.B(n_7920),
.Y(n_8241)
);

AND2x2_ASAP7_75t_L g8242 ( 
.A(n_8072),
.B(n_7992),
.Y(n_8242)
);

NAND4xp25_ASAP7_75t_L g8243 ( 
.A(n_8087),
.B(n_7931),
.C(n_7986),
.D(n_7983),
.Y(n_8243)
);

INVx2_ASAP7_75t_L g8244 ( 
.A(n_8150),
.Y(n_8244)
);

NAND2xp5_ASAP7_75t_L g8245 ( 
.A(n_8078),
.B(n_7898),
.Y(n_8245)
);

INVx1_ASAP7_75t_L g8246 ( 
.A(n_8080),
.Y(n_8246)
);

AND2x2_ASAP7_75t_L g8247 ( 
.A(n_8055),
.B(n_7957),
.Y(n_8247)
);

INVx1_ASAP7_75t_L g8248 ( 
.A(n_8111),
.Y(n_8248)
);

AND2x2_ASAP7_75t_L g8249 ( 
.A(n_8058),
.B(n_7958),
.Y(n_8249)
);

NAND2xp5_ASAP7_75t_L g8250 ( 
.A(n_8150),
.B(n_7993),
.Y(n_8250)
);

AND2x2_ASAP7_75t_SL g8251 ( 
.A(n_8094),
.B(n_7931),
.Y(n_8251)
);

INVx1_ASAP7_75t_L g8252 ( 
.A(n_8065),
.Y(n_8252)
);

NOR2x1p5_ASAP7_75t_L g8253 ( 
.A(n_8042),
.B(n_8033),
.Y(n_8253)
);

AND2x2_ASAP7_75t_L g8254 ( 
.A(n_8096),
.B(n_7998),
.Y(n_8254)
);

INVx1_ASAP7_75t_L g8255 ( 
.A(n_8060),
.Y(n_8255)
);

O2A1O1Ixp5_ASAP7_75t_R g8256 ( 
.A1(n_8037),
.A2(n_7986),
.B(n_7983),
.C(n_7343),
.Y(n_8256)
);

INVx2_ASAP7_75t_L g8257 ( 
.A(n_8057),
.Y(n_8257)
);

OAI22xp33_ASAP7_75t_L g8258 ( 
.A1(n_8061),
.A2(n_6905),
.B1(n_6677),
.B2(n_6975),
.Y(n_8258)
);

NAND2xp5_ASAP7_75t_L g8259 ( 
.A(n_8052),
.B(n_8000),
.Y(n_8259)
);

INVx2_ASAP7_75t_L g8260 ( 
.A(n_8149),
.Y(n_8260)
);

INVx1_ASAP7_75t_L g8261 ( 
.A(n_8075),
.Y(n_8261)
);

INVx1_ASAP7_75t_SL g8262 ( 
.A(n_8133),
.Y(n_8262)
);

NOR2xp33_ASAP7_75t_L g8263 ( 
.A(n_8120),
.B(n_8005),
.Y(n_8263)
);

INVx1_ASAP7_75t_L g8264 ( 
.A(n_8165),
.Y(n_8264)
);

OAI21xp5_ASAP7_75t_SL g8265 ( 
.A1(n_8061),
.A2(n_6801),
.B(n_6791),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_8147),
.Y(n_8266)
);

AOI21xp33_ASAP7_75t_SL g8267 ( 
.A1(n_8161),
.A2(n_7357),
.B(n_7351),
.Y(n_8267)
);

INVx1_ASAP7_75t_L g8268 ( 
.A(n_8166),
.Y(n_8268)
);

INVxp67_ASAP7_75t_L g8269 ( 
.A(n_8077),
.Y(n_8269)
);

NAND2xp5_ASAP7_75t_L g8270 ( 
.A(n_8054),
.B(n_6943),
.Y(n_8270)
);

OR2x2_ASAP7_75t_L g8271 ( 
.A(n_8101),
.B(n_7084),
.Y(n_8271)
);

NAND2xp5_ASAP7_75t_L g8272 ( 
.A(n_8120),
.B(n_6952),
.Y(n_8272)
);

INVx2_ASAP7_75t_L g8273 ( 
.A(n_8084),
.Y(n_8273)
);

OR2x2_ASAP7_75t_L g8274 ( 
.A(n_8106),
.B(n_7028),
.Y(n_8274)
);

INVx1_ASAP7_75t_L g8275 ( 
.A(n_8048),
.Y(n_8275)
);

INVx2_ASAP7_75t_L g8276 ( 
.A(n_8088),
.Y(n_8276)
);

A2O1A1Ixp33_ASAP7_75t_L g8277 ( 
.A1(n_8108),
.A2(n_6810),
.B(n_6791),
.C(n_6905),
.Y(n_8277)
);

INVxp33_ASAP7_75t_L g8278 ( 
.A(n_8097),
.Y(n_8278)
);

NOR2xp33_ASAP7_75t_L g8279 ( 
.A(n_8024),
.B(n_7085),
.Y(n_8279)
);

INVx1_ASAP7_75t_L g8280 ( 
.A(n_8100),
.Y(n_8280)
);

AND2x2_ASAP7_75t_L g8281 ( 
.A(n_8104),
.B(n_7062),
.Y(n_8281)
);

INVx1_ASAP7_75t_SL g8282 ( 
.A(n_8122),
.Y(n_8282)
);

AND2x2_ASAP7_75t_L g8283 ( 
.A(n_8025),
.B(n_7062),
.Y(n_8283)
);

INVxp67_ASAP7_75t_L g8284 ( 
.A(n_8144),
.Y(n_8284)
);

AND2x4_ASAP7_75t_L g8285 ( 
.A(n_8083),
.B(n_7062),
.Y(n_8285)
);

NAND2xp5_ASAP7_75t_L g8286 ( 
.A(n_8146),
.B(n_6963),
.Y(n_8286)
);

INVx1_ASAP7_75t_L g8287 ( 
.A(n_8154),
.Y(n_8287)
);

INVx3_ASAP7_75t_L g8288 ( 
.A(n_8099),
.Y(n_8288)
);

INVx2_ASAP7_75t_L g8289 ( 
.A(n_8103),
.Y(n_8289)
);

BUFx2_ASAP7_75t_SL g8290 ( 
.A(n_8130),
.Y(n_8290)
);

INVx2_ASAP7_75t_SL g8291 ( 
.A(n_8132),
.Y(n_8291)
);

INVx1_ASAP7_75t_L g8292 ( 
.A(n_8092),
.Y(n_8292)
);

NAND2xp5_ASAP7_75t_L g8293 ( 
.A(n_8045),
.B(n_8102),
.Y(n_8293)
);

INVx1_ASAP7_75t_L g8294 ( 
.A(n_8125),
.Y(n_8294)
);

INVx1_ASAP7_75t_L g8295 ( 
.A(n_8139),
.Y(n_8295)
);

NAND2xp5_ASAP7_75t_L g8296 ( 
.A(n_8136),
.B(n_6965),
.Y(n_8296)
);

OR2x2_ASAP7_75t_L g8297 ( 
.A(n_8135),
.B(n_8137),
.Y(n_8297)
);

AND2x2_ASAP7_75t_L g8298 ( 
.A(n_8152),
.B(n_7080),
.Y(n_8298)
);

OAI21xp33_ASAP7_75t_L g8299 ( 
.A1(n_8108),
.A2(n_6969),
.B(n_6959),
.Y(n_8299)
);

NAND2xp5_ASAP7_75t_L g8300 ( 
.A(n_8136),
.B(n_6967),
.Y(n_8300)
);

AND2x2_ASAP7_75t_L g8301 ( 
.A(n_8163),
.B(n_7080),
.Y(n_8301)
);

NAND2x1_ASAP7_75t_SL g8302 ( 
.A(n_8128),
.B(n_7080),
.Y(n_8302)
);

AND2x2_ASAP7_75t_L g8303 ( 
.A(n_8127),
.B(n_6707),
.Y(n_8303)
);

INVx2_ASAP7_75t_L g8304 ( 
.A(n_8016),
.Y(n_8304)
);

AND2x4_ASAP7_75t_L g8305 ( 
.A(n_8157),
.B(n_6581),
.Y(n_8305)
);

AND2x4_ASAP7_75t_L g8306 ( 
.A(n_8134),
.B(n_6586),
.Y(n_8306)
);

NOR2xp33_ASAP7_75t_L g8307 ( 
.A(n_8135),
.B(n_7054),
.Y(n_8307)
);

INVxp67_ASAP7_75t_SL g8308 ( 
.A(n_8014),
.Y(n_8308)
);

AND2x2_ASAP7_75t_SL g8309 ( 
.A(n_8141),
.B(n_7035),
.Y(n_8309)
);

AND2x2_ASAP7_75t_L g8310 ( 
.A(n_8119),
.B(n_6664),
.Y(n_8310)
);

NAND2xp5_ASAP7_75t_L g8311 ( 
.A(n_8167),
.B(n_8019),
.Y(n_8311)
);

NAND2xp5_ASAP7_75t_L g8312 ( 
.A(n_8170),
.B(n_8066),
.Y(n_8312)
);

AOI21xp33_ASAP7_75t_SL g8313 ( 
.A1(n_8211),
.A2(n_8251),
.B(n_8239),
.Y(n_8313)
);

AOI22xp33_ASAP7_75t_SL g8314 ( 
.A1(n_8169),
.A2(n_8008),
.B1(n_8143),
.B2(n_8140),
.Y(n_8314)
);

INVx1_ASAP7_75t_L g8315 ( 
.A(n_8221),
.Y(n_8315)
);

INVx2_ASAP7_75t_L g8316 ( 
.A(n_8185),
.Y(n_8316)
);

OAI322xp33_ASAP7_75t_L g8317 ( 
.A1(n_8169),
.A2(n_8158),
.A3(n_8070),
.B1(n_8159),
.B2(n_8162),
.C1(n_8123),
.C2(n_8129),
.Y(n_8317)
);

NAND2xp5_ASAP7_75t_SL g8318 ( 
.A(n_8197),
.B(n_8140),
.Y(n_8318)
);

OR2x2_ASAP7_75t_L g8319 ( 
.A(n_8190),
.B(n_8126),
.Y(n_8319)
);

INVx1_ASAP7_75t_L g8320 ( 
.A(n_8252),
.Y(n_8320)
);

OAI221xp5_ASAP7_75t_L g8321 ( 
.A1(n_8198),
.A2(n_8202),
.B1(n_8179),
.B2(n_8302),
.C(n_8308),
.Y(n_8321)
);

NAND2x1_ASAP7_75t_SL g8322 ( 
.A(n_8229),
.B(n_8128),
.Y(n_8322)
);

AOI22xp5_ASAP7_75t_L g8323 ( 
.A1(n_8202),
.A2(n_8142),
.B1(n_8091),
.B2(n_8145),
.Y(n_8323)
);

INVx1_ASAP7_75t_L g8324 ( 
.A(n_8168),
.Y(n_8324)
);

INVx1_ASAP7_75t_L g8325 ( 
.A(n_8303),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_8216),
.Y(n_8326)
);

INVx1_ASAP7_75t_L g8327 ( 
.A(n_8192),
.Y(n_8327)
);

INVx2_ASAP7_75t_L g8328 ( 
.A(n_8229),
.Y(n_8328)
);

NOR2xp33_ASAP7_75t_L g8329 ( 
.A(n_8278),
.B(n_8142),
.Y(n_8329)
);

INVx1_ASAP7_75t_L g8330 ( 
.A(n_8283),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_8174),
.Y(n_8331)
);

AND2x2_ASAP7_75t_L g8332 ( 
.A(n_8298),
.B(n_8079),
.Y(n_8332)
);

AOI22xp33_ASAP7_75t_L g8333 ( 
.A1(n_8173),
.A2(n_6472),
.B1(n_6445),
.B2(n_6760),
.Y(n_8333)
);

AND2x2_ASAP7_75t_L g8334 ( 
.A(n_8281),
.B(n_8085),
.Y(n_8334)
);

OR2x2_ASAP7_75t_L g8335 ( 
.A(n_8190),
.B(n_8105),
.Y(n_8335)
);

OR2x2_ASAP7_75t_L g8336 ( 
.A(n_8290),
.B(n_8124),
.Y(n_8336)
);

OAI21xp5_ASAP7_75t_SL g8337 ( 
.A1(n_8188),
.A2(n_8158),
.B(n_8151),
.Y(n_8337)
);

INVx2_ASAP7_75t_L g8338 ( 
.A(n_8305),
.Y(n_8338)
);

NAND2xp5_ASAP7_75t_L g8339 ( 
.A(n_8305),
.B(n_8138),
.Y(n_8339)
);

INVx1_ASAP7_75t_L g8340 ( 
.A(n_8196),
.Y(n_8340)
);

INVx2_ASAP7_75t_L g8341 ( 
.A(n_8285),
.Y(n_8341)
);

OAI221xp5_ASAP7_75t_L g8342 ( 
.A1(n_8179),
.A2(n_8160),
.B1(n_8156),
.B2(n_8113),
.C(n_8112),
.Y(n_8342)
);

OAI22xp5_ASAP7_75t_L g8343 ( 
.A1(n_8248),
.A2(n_7066),
.B1(n_6920),
.B2(n_7087),
.Y(n_8343)
);

INVx1_ASAP7_75t_L g8344 ( 
.A(n_8200),
.Y(n_8344)
);

AND2x2_ASAP7_75t_L g8345 ( 
.A(n_8301),
.B(n_8161),
.Y(n_8345)
);

INVx1_ASAP7_75t_L g8346 ( 
.A(n_8285),
.Y(n_8346)
);

INVx1_ASAP7_75t_L g8347 ( 
.A(n_8306),
.Y(n_8347)
);

NAND2xp5_ASAP7_75t_L g8348 ( 
.A(n_8306),
.B(n_8197),
.Y(n_8348)
);

INVx2_ASAP7_75t_L g8349 ( 
.A(n_8181),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_8199),
.Y(n_8350)
);

INVx1_ASAP7_75t_L g8351 ( 
.A(n_8180),
.Y(n_8351)
);

NAND2xp5_ASAP7_75t_L g8352 ( 
.A(n_8181),
.B(n_6980),
.Y(n_8352)
);

AOI22xp5_ASAP7_75t_L g8353 ( 
.A1(n_8243),
.A2(n_6988),
.B1(n_6996),
.B2(n_6987),
.Y(n_8353)
);

INVx2_ASAP7_75t_L g8354 ( 
.A(n_8194),
.Y(n_8354)
);

NOR2xp33_ASAP7_75t_L g8355 ( 
.A(n_8223),
.B(n_6997),
.Y(n_8355)
);

INVx1_ASAP7_75t_L g8356 ( 
.A(n_8191),
.Y(n_8356)
);

OAI21xp5_ASAP7_75t_SL g8357 ( 
.A1(n_8262),
.A2(n_7013),
.B(n_7002),
.Y(n_8357)
);

OAI21xp5_ASAP7_75t_L g8358 ( 
.A1(n_8175),
.A2(n_7009),
.B(n_7006),
.Y(n_8358)
);

AOI21xp33_ASAP7_75t_L g8359 ( 
.A1(n_8220),
.A2(n_7015),
.B(n_7047),
.Y(n_8359)
);

OAI322xp33_ASAP7_75t_L g8360 ( 
.A1(n_8234),
.A2(n_7024),
.A3(n_7027),
.B1(n_7041),
.B2(n_7038),
.C1(n_7061),
.C2(n_7043),
.Y(n_8360)
);

OR2x2_ASAP7_75t_L g8361 ( 
.A(n_8243),
.B(n_7073),
.Y(n_8361)
);

OR2x2_ASAP7_75t_L g8362 ( 
.A(n_8184),
.B(n_7076),
.Y(n_8362)
);

AND2x2_ASAP7_75t_L g8363 ( 
.A(n_8195),
.B(n_6664),
.Y(n_8363)
);

HB1xp67_ASAP7_75t_L g8364 ( 
.A(n_8288),
.Y(n_8364)
);

INVx2_ASAP7_75t_SL g8365 ( 
.A(n_8201),
.Y(n_8365)
);

INVx1_ASAP7_75t_L g8366 ( 
.A(n_8207),
.Y(n_8366)
);

NAND2xp5_ASAP7_75t_L g8367 ( 
.A(n_8224),
.B(n_8234),
.Y(n_8367)
);

INVx2_ASAP7_75t_L g8368 ( 
.A(n_8288),
.Y(n_8368)
);

INVx1_ASAP7_75t_L g8369 ( 
.A(n_8209),
.Y(n_8369)
);

OAI22xp5_ASAP7_75t_L g8370 ( 
.A1(n_8284),
.A2(n_6869),
.B1(n_6767),
.B2(n_6766),
.Y(n_8370)
);

INVx1_ASAP7_75t_L g8371 ( 
.A(n_8186),
.Y(n_8371)
);

AND2x2_ASAP7_75t_L g8372 ( 
.A(n_8218),
.B(n_6665),
.Y(n_8372)
);

INVx1_ASAP7_75t_L g8373 ( 
.A(n_8214),
.Y(n_8373)
);

INVx1_ASAP7_75t_L g8374 ( 
.A(n_8187),
.Y(n_8374)
);

OAI221xp5_ASAP7_75t_L g8375 ( 
.A1(n_8182),
.A2(n_7086),
.B1(n_7081),
.B2(n_7016),
.C(n_6449),
.Y(n_8375)
);

OR2x2_ASAP7_75t_L g8376 ( 
.A(n_8230),
.B(n_6431),
.Y(n_8376)
);

AND2x2_ASAP7_75t_L g8377 ( 
.A(n_8225),
.B(n_6665),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_8177),
.Y(n_8378)
);

AND2x2_ASAP7_75t_L g8379 ( 
.A(n_8238),
.B(n_6666),
.Y(n_8379)
);

AOI21xp5_ASAP7_75t_L g8380 ( 
.A1(n_8222),
.A2(n_6472),
.B(n_6445),
.Y(n_8380)
);

INVx1_ASAP7_75t_L g8381 ( 
.A(n_8254),
.Y(n_8381)
);

INVx1_ASAP7_75t_L g8382 ( 
.A(n_8244),
.Y(n_8382)
);

INVx1_ASAP7_75t_L g8383 ( 
.A(n_8193),
.Y(n_8383)
);

NAND2xp5_ASAP7_75t_L g8384 ( 
.A(n_8241),
.B(n_6586),
.Y(n_8384)
);

AND2x2_ASAP7_75t_L g8385 ( 
.A(n_8204),
.B(n_6666),
.Y(n_8385)
);

NAND2xp5_ASAP7_75t_SL g8386 ( 
.A(n_8241),
.B(n_6449),
.Y(n_8386)
);

NAND2xp5_ASAP7_75t_L g8387 ( 
.A(n_8291),
.B(n_6586),
.Y(n_8387)
);

AOI32xp33_ASAP7_75t_L g8388 ( 
.A1(n_8282),
.A2(n_6861),
.A3(n_6852),
.B1(n_6471),
.B2(n_6473),
.Y(n_8388)
);

INVx1_ASAP7_75t_L g8389 ( 
.A(n_8236),
.Y(n_8389)
);

NAND2xp5_ASAP7_75t_L g8390 ( 
.A(n_8215),
.B(n_6603),
.Y(n_8390)
);

AOI221xp5_ASAP7_75t_L g8391 ( 
.A1(n_8267),
.A2(n_6469),
.B1(n_6473),
.B2(n_6471),
.C(n_6465),
.Y(n_8391)
);

OAI31xp33_ASAP7_75t_L g8392 ( 
.A1(n_8265),
.A2(n_6852),
.A3(n_6603),
.B(n_6469),
.Y(n_8392)
);

INVx1_ASAP7_75t_L g8393 ( 
.A(n_8189),
.Y(n_8393)
);

AOI22xp5_ASAP7_75t_L g8394 ( 
.A1(n_8263),
.A2(n_8307),
.B1(n_8213),
.B2(n_8228),
.Y(n_8394)
);

INVx1_ASAP7_75t_L g8395 ( 
.A(n_8250),
.Y(n_8395)
);

OAI21xp5_ASAP7_75t_L g8396 ( 
.A1(n_8172),
.A2(n_6477),
.B(n_6465),
.Y(n_8396)
);

NAND2xp5_ASAP7_75t_L g8397 ( 
.A(n_8206),
.B(n_8264),
.Y(n_8397)
);

NAND2xp5_ASAP7_75t_L g8398 ( 
.A(n_8287),
.B(n_6603),
.Y(n_8398)
);

OAI21xp5_ASAP7_75t_L g8399 ( 
.A1(n_8203),
.A2(n_6481),
.B(n_6477),
.Y(n_8399)
);

NAND3xp33_ASAP7_75t_L g8400 ( 
.A(n_8228),
.B(n_6516),
.C(n_6514),
.Y(n_8400)
);

O2A1O1Ixp33_ASAP7_75t_SL g8401 ( 
.A1(n_8277),
.A2(n_6481),
.B(n_6484),
.C(n_6591),
.Y(n_8401)
);

AOI21xp5_ASAP7_75t_L g8402 ( 
.A1(n_8219),
.A2(n_6472),
.B(n_6445),
.Y(n_8402)
);

OR2x2_ASAP7_75t_L g8403 ( 
.A(n_8271),
.B(n_6438),
.Y(n_8403)
);

AOI222xp33_ASAP7_75t_L g8404 ( 
.A1(n_8299),
.A2(n_6484),
.B1(n_6543),
.B2(n_6546),
.C1(n_6542),
.C2(n_6520),
.Y(n_8404)
);

NAND2xp5_ASAP7_75t_SL g8405 ( 
.A(n_8309),
.B(n_6591),
.Y(n_8405)
);

AND2x2_ASAP7_75t_L g8406 ( 
.A(n_8310),
.B(n_6669),
.Y(n_8406)
);

AOI211xp5_ASAP7_75t_L g8407 ( 
.A1(n_8267),
.A2(n_6576),
.B(n_6583),
.C(n_6578),
.Y(n_8407)
);

NAND2x1_ASAP7_75t_SL g8408 ( 
.A(n_8256),
.B(n_6596),
.Y(n_8408)
);

INVx1_ASAP7_75t_L g8409 ( 
.A(n_8235),
.Y(n_8409)
);

INVx1_ASAP7_75t_L g8410 ( 
.A(n_8240),
.Y(n_8410)
);

INVx1_ASAP7_75t_L g8411 ( 
.A(n_8247),
.Y(n_8411)
);

AOI322xp5_ASAP7_75t_L g8412 ( 
.A1(n_8299),
.A2(n_6582),
.A3(n_6595),
.B1(n_6601),
.B2(n_6607),
.C1(n_6599),
.C2(n_6588),
.Y(n_8412)
);

NAND2xp5_ASAP7_75t_L g8413 ( 
.A(n_8266),
.B(n_6757),
.Y(n_8413)
);

NAND2xp5_ASAP7_75t_L g8414 ( 
.A(n_8249),
.B(n_6553),
.Y(n_8414)
);

INVx2_ASAP7_75t_L g8415 ( 
.A(n_8253),
.Y(n_8415)
);

OAI32xp33_ASAP7_75t_L g8416 ( 
.A1(n_8297),
.A2(n_6606),
.A3(n_6600),
.B1(n_6596),
.B2(n_6766),
.Y(n_8416)
);

INVx1_ASAP7_75t_L g8417 ( 
.A(n_8242),
.Y(n_8417)
);

INVx2_ASAP7_75t_SL g8418 ( 
.A(n_8233),
.Y(n_8418)
);

OAI222xp33_ASAP7_75t_L g8419 ( 
.A1(n_8183),
.A2(n_6606),
.B1(n_6600),
.B2(n_6767),
.C1(n_6242),
.C2(n_6224),
.Y(n_8419)
);

INVx2_ASAP7_75t_SL g8420 ( 
.A(n_8276),
.Y(n_8420)
);

OAI221xp5_ASAP7_75t_L g8421 ( 
.A1(n_8178),
.A2(n_6698),
.B1(n_6770),
.B2(n_6649),
.C(n_6615),
.Y(n_8421)
);

INVx1_ASAP7_75t_L g8422 ( 
.A(n_8272),
.Y(n_8422)
);

OAI21xp5_ASAP7_75t_L g8423 ( 
.A1(n_8232),
.A2(n_6721),
.B(n_6736),
.Y(n_8423)
);

OR2x2_ASAP7_75t_L g8424 ( 
.A(n_8260),
.B(n_6438),
.Y(n_8424)
);

NAND2xp5_ASAP7_75t_L g8425 ( 
.A(n_8289),
.B(n_6553),
.Y(n_8425)
);

INVx1_ASAP7_75t_L g8426 ( 
.A(n_8296),
.Y(n_8426)
);

AND2x2_ASAP7_75t_L g8427 ( 
.A(n_8273),
.B(n_6669),
.Y(n_8427)
);

AOI222xp33_ASAP7_75t_L g8428 ( 
.A1(n_8265),
.A2(n_8300),
.B1(n_8268),
.B2(n_8295),
.C1(n_8261),
.C2(n_8255),
.Y(n_8428)
);

INVx1_ASAP7_75t_SL g8429 ( 
.A(n_8274),
.Y(n_8429)
);

INVx1_ASAP7_75t_L g8430 ( 
.A(n_8210),
.Y(n_8430)
);

INVx1_ASAP7_75t_L g8431 ( 
.A(n_8231),
.Y(n_8431)
);

INVx1_ASAP7_75t_SL g8432 ( 
.A(n_8286),
.Y(n_8432)
);

INVx1_ASAP7_75t_L g8433 ( 
.A(n_8293),
.Y(n_8433)
);

AOI22xp33_ASAP7_75t_L g8434 ( 
.A1(n_8257),
.A2(n_6531),
.B1(n_6721),
.B2(n_6736),
.Y(n_8434)
);

HB1xp67_ASAP7_75t_L g8435 ( 
.A(n_8364),
.Y(n_8435)
);

OR2x2_ASAP7_75t_L g8436 ( 
.A(n_8376),
.B(n_8275),
.Y(n_8436)
);

INVxp67_ASAP7_75t_L g8437 ( 
.A(n_8348),
.Y(n_8437)
);

NAND2xp5_ASAP7_75t_L g8438 ( 
.A(n_8316),
.B(n_8176),
.Y(n_8438)
);

OAI221xp5_ASAP7_75t_L g8439 ( 
.A1(n_8314),
.A2(n_8237),
.B1(n_8269),
.B2(n_8245),
.C(n_8217),
.Y(n_8439)
);

OAI21xp5_ASAP7_75t_SL g8440 ( 
.A1(n_8394),
.A2(n_8313),
.B(n_8337),
.Y(n_8440)
);

NAND2xp5_ASAP7_75t_L g8441 ( 
.A(n_8346),
.B(n_8171),
.Y(n_8441)
);

INVx1_ASAP7_75t_L g8442 ( 
.A(n_8384),
.Y(n_8442)
);

INVx1_ASAP7_75t_SL g8443 ( 
.A(n_8322),
.Y(n_8443)
);

AND2x2_ASAP7_75t_L g8444 ( 
.A(n_8363),
.B(n_8208),
.Y(n_8444)
);

NOR2xp33_ASAP7_75t_L g8445 ( 
.A(n_8349),
.B(n_8294),
.Y(n_8445)
);

AND2x2_ASAP7_75t_L g8446 ( 
.A(n_8372),
.B(n_8212),
.Y(n_8446)
);

NAND2xp5_ASAP7_75t_L g8447 ( 
.A(n_8341),
.B(n_8279),
.Y(n_8447)
);

NAND4xp25_ASAP7_75t_L g8448 ( 
.A(n_8329),
.B(n_8246),
.C(n_8226),
.D(n_8259),
.Y(n_8448)
);

NAND2xp5_ASAP7_75t_L g8449 ( 
.A(n_8388),
.B(n_8205),
.Y(n_8449)
);

NAND2xp5_ASAP7_75t_SL g8450 ( 
.A(n_8338),
.B(n_8258),
.Y(n_8450)
);

AOI21xp5_ASAP7_75t_L g8451 ( 
.A1(n_8380),
.A2(n_8270),
.B(n_8292),
.Y(n_8451)
);

INVx1_ASAP7_75t_L g8452 ( 
.A(n_8414),
.Y(n_8452)
);

INVx1_ASAP7_75t_L g8453 ( 
.A(n_8387),
.Y(n_8453)
);

INVx2_ASAP7_75t_L g8454 ( 
.A(n_8424),
.Y(n_8454)
);

AOI21xp33_ASAP7_75t_SL g8455 ( 
.A1(n_8318),
.A2(n_8227),
.B(n_8304),
.Y(n_8455)
);

NAND2xp5_ASAP7_75t_L g8456 ( 
.A(n_8347),
.B(n_8280),
.Y(n_8456)
);

INVx1_ASAP7_75t_SL g8457 ( 
.A(n_8403),
.Y(n_8457)
);

INVx2_ASAP7_75t_L g8458 ( 
.A(n_8365),
.Y(n_8458)
);

AOI22xp5_ASAP7_75t_L g8459 ( 
.A1(n_8324),
.A2(n_6535),
.B1(n_6580),
.B2(n_6745),
.Y(n_8459)
);

NOR2x1_ASAP7_75t_SL g8460 ( 
.A(n_8405),
.B(n_8386),
.Y(n_8460)
);

NOR2xp33_ASAP7_75t_L g8461 ( 
.A(n_8321),
.B(n_6634),
.Y(n_8461)
);

AND2x2_ASAP7_75t_L g8462 ( 
.A(n_8377),
.B(n_6567),
.Y(n_8462)
);

AOI21xp5_ASAP7_75t_L g8463 ( 
.A1(n_8402),
.A2(n_6531),
.B(n_6610),
.Y(n_8463)
);

NAND2xp5_ASAP7_75t_L g8464 ( 
.A(n_8345),
.B(n_6535),
.Y(n_8464)
);

INVx3_ASAP7_75t_L g8465 ( 
.A(n_8368),
.Y(n_8465)
);

OAI22xp33_ASAP7_75t_L g8466 ( 
.A1(n_8394),
.A2(n_6224),
.B1(n_6243),
.B2(n_6236),
.Y(n_8466)
);

NOR2xp33_ASAP7_75t_L g8467 ( 
.A(n_8330),
.B(n_6763),
.Y(n_8467)
);

INVx2_ASAP7_75t_SL g8468 ( 
.A(n_8379),
.Y(n_8468)
);

INVx1_ASAP7_75t_L g8469 ( 
.A(n_8398),
.Y(n_8469)
);

NOR2xp67_ASAP7_75t_L g8470 ( 
.A(n_8400),
.B(n_8418),
.Y(n_8470)
);

INVxp33_ASAP7_75t_L g8471 ( 
.A(n_8425),
.Y(n_8471)
);

INVx1_ASAP7_75t_L g8472 ( 
.A(n_8390),
.Y(n_8472)
);

NAND2xp5_ASAP7_75t_SL g8473 ( 
.A(n_8323),
.B(n_6535),
.Y(n_8473)
);

A2O1A1Ixp33_ASAP7_75t_SL g8474 ( 
.A1(n_8342),
.A2(n_6251),
.B(n_6248),
.C(n_6611),
.Y(n_8474)
);

OAI21xp33_ASAP7_75t_L g8475 ( 
.A1(n_8351),
.A2(n_6705),
.B(n_6723),
.Y(n_8475)
);

AOI32xp33_ASAP7_75t_L g8476 ( 
.A1(n_8344),
.A2(n_6705),
.A3(n_6745),
.B1(n_6752),
.B2(n_6723),
.Y(n_8476)
);

INVx1_ASAP7_75t_L g8477 ( 
.A(n_8385),
.Y(n_8477)
);

AOI21xp33_ASAP7_75t_L g8478 ( 
.A1(n_8428),
.A2(n_6531),
.B(n_6614),
.Y(n_8478)
);

INVxp67_ASAP7_75t_L g8479 ( 
.A(n_8427),
.Y(n_8479)
);

NAND2xp33_ASAP7_75t_SL g8480 ( 
.A(n_8408),
.B(n_8335),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_8406),
.Y(n_8481)
);

OAI22xp33_ASAP7_75t_L g8482 ( 
.A1(n_8323),
.A2(n_6248),
.B1(n_6251),
.B2(n_6624),
.Y(n_8482)
);

OAI332xp33_ASAP7_75t_L g8483 ( 
.A1(n_8420),
.A2(n_6754),
.A3(n_6742),
.B1(n_6761),
.B2(n_6749),
.B3(n_6741),
.C1(n_6673),
.C2(n_6689),
.Y(n_8483)
);

AOI21xp5_ASAP7_75t_L g8484 ( 
.A1(n_8367),
.A2(n_6637),
.B(n_6635),
.Y(n_8484)
);

NAND2xp5_ASAP7_75t_L g8485 ( 
.A(n_8434),
.B(n_8325),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_8332),
.Y(n_8486)
);

NAND2xp5_ASAP7_75t_L g8487 ( 
.A(n_8334),
.B(n_6580),
.Y(n_8487)
);

AOI22xp5_ASAP7_75t_L g8488 ( 
.A1(n_8331),
.A2(n_6580),
.B1(n_6752),
.B2(n_6723),
.Y(n_8488)
);

NAND3xp33_ASAP7_75t_L g8489 ( 
.A(n_8333),
.B(n_8400),
.C(n_8315),
.Y(n_8489)
);

INVx1_ASAP7_75t_L g8490 ( 
.A(n_8339),
.Y(n_8490)
);

AND2x2_ASAP7_75t_L g8491 ( 
.A(n_8423),
.B(n_6567),
.Y(n_8491)
);

OAI33xp33_ASAP7_75t_L g8492 ( 
.A1(n_8370),
.A2(n_6700),
.A3(n_6651),
.B1(n_6706),
.B2(n_6692),
.B3(n_6646),
.Y(n_8492)
);

OR2x2_ASAP7_75t_L g8493 ( 
.A(n_8319),
.B(n_6648),
.Y(n_8493)
);

NOR2xp33_ASAP7_75t_L g8494 ( 
.A(n_8373),
.B(n_6718),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_8352),
.Y(n_8495)
);

OAI221xp5_ASAP7_75t_L g8496 ( 
.A1(n_8392),
.A2(n_6727),
.B1(n_6716),
.B2(n_6714),
.C(n_6732),
.Y(n_8496)
);

INVx2_ASAP7_75t_L g8497 ( 
.A(n_8328),
.Y(n_8497)
);

INVx3_ASAP7_75t_L g8498 ( 
.A(n_8336),
.Y(n_8498)
);

INVx1_ASAP7_75t_L g8499 ( 
.A(n_8413),
.Y(n_8499)
);

NAND2xp5_ASAP7_75t_L g8500 ( 
.A(n_8350),
.B(n_6738),
.Y(n_8500)
);

INVx2_ASAP7_75t_L g8501 ( 
.A(n_8361),
.Y(n_8501)
);

AO22x1_ASAP7_75t_L g8502 ( 
.A1(n_8366),
.A2(n_6769),
.B1(n_6740),
.B2(n_6752),
.Y(n_8502)
);

INVx1_ASAP7_75t_L g8503 ( 
.A(n_8326),
.Y(n_8503)
);

INVx1_ASAP7_75t_L g8504 ( 
.A(n_8369),
.Y(n_8504)
);

AND2x2_ASAP7_75t_L g8505 ( 
.A(n_8381),
.B(n_7053),
.Y(n_8505)
);

OAI21xp33_ASAP7_75t_L g8506 ( 
.A1(n_8356),
.A2(n_7053),
.B(n_7045),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_8311),
.Y(n_8507)
);

AOI22xp5_ASAP7_75t_L g8508 ( 
.A1(n_8327),
.A2(n_7045),
.B1(n_6356),
.B2(n_6375),
.Y(n_8508)
);

NOR2xp33_ASAP7_75t_L g8509 ( 
.A(n_8359),
.B(n_6648),
.Y(n_8509)
);

NAND4xp25_ASAP7_75t_L g8510 ( 
.A(n_8358),
.B(n_6658),
.C(n_6768),
.D(n_6054),
.Y(n_8510)
);

INVx1_ASAP7_75t_L g8511 ( 
.A(n_8397),
.Y(n_8511)
);

INVx1_ASAP7_75t_L g8512 ( 
.A(n_8312),
.Y(n_8512)
);

INVx2_ASAP7_75t_L g8513 ( 
.A(n_8411),
.Y(n_8513)
);

HB1xp67_ASAP7_75t_L g8514 ( 
.A(n_8343),
.Y(n_8514)
);

INVx1_ASAP7_75t_SL g8515 ( 
.A(n_8429),
.Y(n_8515)
);

NAND2xp5_ASAP7_75t_L g8516 ( 
.A(n_8417),
.B(n_6658),
.Y(n_8516)
);

AOI21xp5_ASAP7_75t_SL g8517 ( 
.A1(n_8317),
.A2(n_6285),
.B(n_6394),
.Y(n_8517)
);

INVx2_ASAP7_75t_L g8518 ( 
.A(n_8362),
.Y(n_8518)
);

INVxp67_ASAP7_75t_L g8519 ( 
.A(n_8355),
.Y(n_8519)
);

NOR4xp25_ASAP7_75t_SL g8520 ( 
.A(n_8357),
.B(n_6184),
.C(n_6196),
.D(n_6172),
.Y(n_8520)
);

NAND3xp33_ASAP7_75t_L g8521 ( 
.A(n_8320),
.B(n_6394),
.C(n_6285),
.Y(n_8521)
);

OAI22xp33_ASAP7_75t_L g8522 ( 
.A1(n_8409),
.A2(n_8410),
.B1(n_8353),
.B2(n_8354),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_8396),
.Y(n_8523)
);

HB1xp67_ASAP7_75t_L g8524 ( 
.A(n_8399),
.Y(n_8524)
);

OAI222xp33_ASAP7_75t_L g8525 ( 
.A1(n_8375),
.A2(n_6285),
.B1(n_6394),
.B2(n_6054),
.C1(n_6061),
.C2(n_6069),
.Y(n_8525)
);

AOI21xp5_ASAP7_75t_L g8526 ( 
.A1(n_8317),
.A2(n_6061),
.B(n_6051),
.Y(n_8526)
);

INVx1_ASAP7_75t_L g8527 ( 
.A(n_8401),
.Y(n_8527)
);

AOI22xp33_ASAP7_75t_L g8528 ( 
.A1(n_8383),
.A2(n_6067),
.B1(n_6069),
.B2(n_6051),
.Y(n_8528)
);

O2A1O1Ixp33_ASAP7_75t_SL g8529 ( 
.A1(n_8389),
.A2(n_8416),
.B(n_8419),
.C(n_8407),
.Y(n_8529)
);

OAI221xp5_ASAP7_75t_L g8530 ( 
.A1(n_8353),
.A2(n_6768),
.B1(n_6394),
.B2(n_6285),
.C(n_6577),
.Y(n_8530)
);

INVx1_ASAP7_75t_L g8531 ( 
.A(n_8360),
.Y(n_8531)
);

INVx2_ASAP7_75t_L g8532 ( 
.A(n_8382),
.Y(n_8532)
);

OAI22xp33_ASAP7_75t_L g8533 ( 
.A1(n_8393),
.A2(n_6577),
.B1(n_6574),
.B2(n_6285),
.Y(n_8533)
);

NOR3xp33_ASAP7_75t_L g8534 ( 
.A(n_8371),
.B(n_6070),
.C(n_6067),
.Y(n_8534)
);

NAND2xp5_ASAP7_75t_L g8535 ( 
.A(n_8378),
.B(n_6574),
.Y(n_8535)
);

INVx1_ASAP7_75t_L g8536 ( 
.A(n_8360),
.Y(n_8536)
);

INVx1_ASAP7_75t_L g8537 ( 
.A(n_8462),
.Y(n_8537)
);

INVx1_ASAP7_75t_L g8538 ( 
.A(n_8505),
.Y(n_8538)
);

NAND2xp5_ASAP7_75t_SL g8539 ( 
.A(n_8443),
.B(n_8391),
.Y(n_8539)
);

INVx1_ASAP7_75t_L g8540 ( 
.A(n_8487),
.Y(n_8540)
);

NAND2xp5_ASAP7_75t_L g8541 ( 
.A(n_8459),
.B(n_8476),
.Y(n_8541)
);

AND2x2_ASAP7_75t_L g8542 ( 
.A(n_8491),
.B(n_8415),
.Y(n_8542)
);

AND2x2_ASAP7_75t_L g8543 ( 
.A(n_8458),
.B(n_8486),
.Y(n_8543)
);

NAND2xp5_ASAP7_75t_L g8544 ( 
.A(n_8488),
.B(n_8432),
.Y(n_8544)
);

INVxp67_ASAP7_75t_L g8545 ( 
.A(n_8435),
.Y(n_8545)
);

NAND2xp5_ASAP7_75t_L g8546 ( 
.A(n_8475),
.B(n_8340),
.Y(n_8546)
);

INVxp67_ASAP7_75t_SL g8547 ( 
.A(n_8473),
.Y(n_8547)
);

NAND2xp5_ASAP7_75t_SL g8548 ( 
.A(n_8493),
.B(n_8404),
.Y(n_8548)
);

AOI22xp33_ASAP7_75t_L g8549 ( 
.A1(n_8506),
.A2(n_8374),
.B1(n_8422),
.B2(n_8395),
.Y(n_8549)
);

OAI221xp5_ASAP7_75t_L g8550 ( 
.A1(n_8440),
.A2(n_8421),
.B1(n_8426),
.B2(n_8433),
.C(n_8430),
.Y(n_8550)
);

AND2x4_ASAP7_75t_SL g8551 ( 
.A(n_8498),
.B(n_8431),
.Y(n_8551)
);

OAI21xp33_ASAP7_75t_L g8552 ( 
.A1(n_8471),
.A2(n_8412),
.B(n_8407),
.Y(n_8552)
);

NAND2xp5_ASAP7_75t_L g8553 ( 
.A(n_8502),
.B(n_8412),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_8464),
.Y(n_8554)
);

AOI21xp33_ASAP7_75t_L g8555 ( 
.A1(n_8457),
.A2(n_6070),
.B(n_6680),
.Y(n_8555)
);

INVxp67_ASAP7_75t_L g8556 ( 
.A(n_8445),
.Y(n_8556)
);

OAI31xp33_ASAP7_75t_L g8557 ( 
.A1(n_8478),
.A2(n_8480),
.A3(n_8439),
.B(n_8489),
.Y(n_8557)
);

OAI32xp33_ASAP7_75t_L g8558 ( 
.A1(n_8485),
.A2(n_6086),
.A3(n_6088),
.B1(n_6087),
.B2(n_6082),
.Y(n_8558)
);

OAI222xp33_ASAP7_75t_L g8559 ( 
.A1(n_8515),
.A2(n_6394),
.B1(n_6165),
.B2(n_6680),
.C1(n_6108),
.C2(n_6225),
.Y(n_8559)
);

INVxp67_ASAP7_75t_SL g8560 ( 
.A(n_8460),
.Y(n_8560)
);

AOI221xp5_ASAP7_75t_L g8561 ( 
.A1(n_8455),
.A2(n_6260),
.B1(n_6225),
.B2(n_6210),
.C(n_6087),
.Y(n_8561)
);

INVxp67_ASAP7_75t_SL g8562 ( 
.A(n_8470),
.Y(n_8562)
);

OR2x2_ASAP7_75t_L g8563 ( 
.A(n_8510),
.B(n_6554),
.Y(n_8563)
);

OAI22xp5_ASAP7_75t_L g8564 ( 
.A1(n_8437),
.A2(n_6086),
.B1(n_6090),
.B2(n_6088),
.Y(n_8564)
);

NAND2xp5_ASAP7_75t_L g8565 ( 
.A(n_8526),
.B(n_6090),
.Y(n_8565)
);

AOI221xp5_ASAP7_75t_L g8566 ( 
.A1(n_8529),
.A2(n_6260),
.B1(n_6225),
.B2(n_6093),
.C(n_6207),
.Y(n_8566)
);

NAND2xp5_ASAP7_75t_SL g8567 ( 
.A(n_8498),
.B(n_6225),
.Y(n_8567)
);

INVx1_ASAP7_75t_SL g8568 ( 
.A(n_8436),
.Y(n_8568)
);

AOI222xp33_ASAP7_75t_L g8569 ( 
.A1(n_8531),
.A2(n_6260),
.B1(n_6375),
.B2(n_6362),
.C1(n_6373),
.C2(n_6093),
.Y(n_8569)
);

INVx1_ASAP7_75t_L g8570 ( 
.A(n_8516),
.Y(n_8570)
);

OAI21xp33_ASAP7_75t_L g8571 ( 
.A1(n_8448),
.A2(n_6260),
.B(n_6207),
.Y(n_8571)
);

AOI32xp33_ASAP7_75t_L g8572 ( 
.A1(n_8503),
.A2(n_6207),
.A3(n_6319),
.B1(n_6375),
.B2(n_6373),
.Y(n_8572)
);

INVx1_ASAP7_75t_L g8573 ( 
.A(n_8535),
.Y(n_8573)
);

INVx2_ASAP7_75t_L g8574 ( 
.A(n_8465),
.Y(n_8574)
);

AOI21xp33_ASAP7_75t_L g8575 ( 
.A1(n_8461),
.A2(n_6022),
.B(n_6044),
.Y(n_8575)
);

BUFx2_ASAP7_75t_L g8576 ( 
.A(n_8465),
.Y(n_8576)
);

OAI22xp5_ASAP7_75t_L g8577 ( 
.A1(n_8528),
.A2(n_6022),
.B1(n_6375),
.B2(n_6196),
.Y(n_8577)
);

NAND2xp5_ASAP7_75t_L g8578 ( 
.A(n_8466),
.B(n_6554),
.Y(n_8578)
);

INVx2_ASAP7_75t_SL g8579 ( 
.A(n_8454),
.Y(n_8579)
);

INVx1_ASAP7_75t_SL g8580 ( 
.A(n_8444),
.Y(n_8580)
);

NOR2xp33_ASAP7_75t_L g8581 ( 
.A(n_8450),
.B(n_6184),
.Y(n_8581)
);

OAI211xp5_ASAP7_75t_L g8582 ( 
.A1(n_8517),
.A2(n_5878),
.B(n_5882),
.C(n_5881),
.Y(n_8582)
);

AND2x2_ASAP7_75t_L g8583 ( 
.A(n_8446),
.B(n_6554),
.Y(n_8583)
);

NAND2xp5_ASAP7_75t_L g8584 ( 
.A(n_8468),
.B(n_6554),
.Y(n_8584)
);

NAND2xp5_ASAP7_75t_L g8585 ( 
.A(n_8482),
.B(n_6554),
.Y(n_8585)
);

NAND3xp33_ASAP7_75t_SL g8586 ( 
.A(n_8463),
.B(n_6319),
.C(n_6083),
.Y(n_8586)
);

INVx1_ASAP7_75t_L g8587 ( 
.A(n_8514),
.Y(n_8587)
);

NAND2xp33_ASAP7_75t_L g8588 ( 
.A(n_8534),
.B(n_6362),
.Y(n_8588)
);

INVx1_ASAP7_75t_L g8589 ( 
.A(n_8527),
.Y(n_8589)
);

AOI22xp5_ASAP7_75t_L g8590 ( 
.A1(n_8481),
.A2(n_6356),
.B1(n_6146),
.B2(n_6168),
.Y(n_8590)
);

OAI21xp5_ASAP7_75t_L g8591 ( 
.A1(n_8479),
.A2(n_8509),
.B(n_8438),
.Y(n_8591)
);

NAND2xp5_ASAP7_75t_L g8592 ( 
.A(n_8536),
.B(n_6617),
.Y(n_8592)
);

OAI211xp5_ASAP7_75t_SL g8593 ( 
.A1(n_8441),
.A2(n_5834),
.B(n_5842),
.C(n_5839),
.Y(n_8593)
);

INVxp67_ASAP7_75t_L g8594 ( 
.A(n_8467),
.Y(n_8594)
);

OAI31xp33_ASAP7_75t_L g8595 ( 
.A1(n_8489),
.A2(n_6322),
.A3(n_6328),
.B(n_6324),
.Y(n_8595)
);

INVx1_ASAP7_75t_L g8596 ( 
.A(n_8524),
.Y(n_8596)
);

NAND2xp5_ASAP7_75t_L g8597 ( 
.A(n_8497),
.B(n_6617),
.Y(n_8597)
);

OAI221xp5_ASAP7_75t_L g8598 ( 
.A1(n_8530),
.A2(n_6165),
.B1(n_5875),
.B2(n_6083),
.C(n_6197),
.Y(n_8598)
);

AOI221x1_ASAP7_75t_L g8599 ( 
.A1(n_8448),
.A2(n_6340),
.B1(n_6343),
.B2(n_6333),
.C(n_6332),
.Y(n_8599)
);

AOI221x1_ASAP7_75t_L g8600 ( 
.A1(n_8451),
.A2(n_6340),
.B1(n_6343),
.B2(n_6333),
.C(n_6332),
.Y(n_8600)
);

AND2x2_ASAP7_75t_L g8601 ( 
.A(n_8513),
.B(n_6617),
.Y(n_8601)
);

INVx1_ASAP7_75t_L g8602 ( 
.A(n_8456),
.Y(n_8602)
);

OAI21xp33_ASAP7_75t_L g8603 ( 
.A1(n_8447),
.A2(n_6207),
.B(n_6146),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_8477),
.Y(n_8604)
);

OAI21xp33_ASAP7_75t_L g8605 ( 
.A1(n_8490),
.A2(n_6168),
.B(n_6282),
.Y(n_8605)
);

AND2x2_ASAP7_75t_L g8606 ( 
.A(n_8532),
.B(n_6617),
.Y(n_8606)
);

NOR3xp33_ASAP7_75t_L g8607 ( 
.A(n_8442),
.B(n_6102),
.C(n_6193),
.Y(n_8607)
);

AND2x2_ASAP7_75t_L g8608 ( 
.A(n_8504),
.B(n_6617),
.Y(n_8608)
);

AOI21xp33_ASAP7_75t_L g8609 ( 
.A1(n_8522),
.A2(n_6044),
.B(n_6076),
.Y(n_8609)
);

OAI322xp33_ASAP7_75t_L g8610 ( 
.A1(n_8533),
.A2(n_6354),
.A3(n_6351),
.B1(n_6357),
.B2(n_6360),
.C1(n_6352),
.C2(n_6345),
.Y(n_8610)
);

NAND2xp5_ASAP7_75t_L g8611 ( 
.A(n_8523),
.B(n_6211),
.Y(n_8611)
);

HB1xp67_ASAP7_75t_L g8612 ( 
.A(n_8521),
.Y(n_8612)
);

AOI21xp5_ASAP7_75t_L g8613 ( 
.A1(n_8449),
.A2(n_6199),
.B(n_6197),
.Y(n_8613)
);

INVx1_ASAP7_75t_L g8614 ( 
.A(n_8500),
.Y(n_8614)
);

INVxp67_ASAP7_75t_SL g8615 ( 
.A(n_8494),
.Y(n_8615)
);

NAND2xp5_ASAP7_75t_L g8616 ( 
.A(n_8474),
.B(n_8484),
.Y(n_8616)
);

OAI22xp5_ASAP7_75t_L g8617 ( 
.A1(n_8508),
.A2(n_6199),
.B1(n_6211),
.B2(n_6206),
.Y(n_8617)
);

INVx1_ASAP7_75t_L g8618 ( 
.A(n_8453),
.Y(n_8618)
);

INVx1_ASAP7_75t_L g8619 ( 
.A(n_8501),
.Y(n_8619)
);

AOI22xp5_ASAP7_75t_L g8620 ( 
.A1(n_8469),
.A2(n_6168),
.B1(n_6282),
.B2(n_6322),
.Y(n_8620)
);

NAND2xp5_ASAP7_75t_L g8621 ( 
.A(n_8483),
.B(n_6253),
.Y(n_8621)
);

AOI21xp33_ASAP7_75t_SL g8622 ( 
.A1(n_8507),
.A2(n_6102),
.B(n_6148),
.Y(n_8622)
);

INVx1_ASAP7_75t_L g8623 ( 
.A(n_8472),
.Y(n_8623)
);

INVx1_ASAP7_75t_L g8624 ( 
.A(n_8511),
.Y(n_8624)
);

INVx1_ASAP7_75t_L g8625 ( 
.A(n_8452),
.Y(n_8625)
);

INVx1_ASAP7_75t_SL g8626 ( 
.A(n_8518),
.Y(n_8626)
);

OAI211xp5_ASAP7_75t_L g8627 ( 
.A1(n_8519),
.A2(n_5980),
.B(n_6328),
.C(n_6324),
.Y(n_8627)
);

AOI322xp5_ASAP7_75t_L g8628 ( 
.A1(n_8547),
.A2(n_8512),
.A3(n_8495),
.B1(n_8499),
.B2(n_8520),
.C1(n_8492),
.C2(n_8525),
.Y(n_8628)
);

CKINVDCx14_ASAP7_75t_R g8629 ( 
.A(n_8576),
.Y(n_8629)
);

NOR2xp33_ASAP7_75t_L g8630 ( 
.A(n_8568),
.B(n_8580),
.Y(n_8630)
);

OAI322xp33_ASAP7_75t_L g8631 ( 
.A1(n_8545),
.A2(n_8496),
.A3(n_8521),
.B1(n_8520),
.B2(n_6357),
.C1(n_6388),
.C2(n_6354),
.Y(n_8631)
);

HB1xp67_ASAP7_75t_L g8632 ( 
.A(n_8583),
.Y(n_8632)
);

AND2x2_ASAP7_75t_L g8633 ( 
.A(n_8543),
.B(n_6168),
.Y(n_8633)
);

OAI22xp33_ASAP7_75t_SL g8634 ( 
.A1(n_8567),
.A2(n_6212),
.B1(n_6213),
.B2(n_6206),
.Y(n_8634)
);

OAI221xp5_ASAP7_75t_L g8635 ( 
.A1(n_8557),
.A2(n_8595),
.B1(n_8603),
.B2(n_8552),
.C(n_8560),
.Y(n_8635)
);

AOI21xp5_ASAP7_75t_L g8636 ( 
.A1(n_8548),
.A2(n_6213),
.B(n_6212),
.Y(n_8636)
);

NOR2xp33_ASAP7_75t_SL g8637 ( 
.A(n_8568),
.B(n_5955),
.Y(n_8637)
);

OAI21xp33_ASAP7_75t_L g8638 ( 
.A1(n_8587),
.A2(n_6351),
.B(n_6345),
.Y(n_8638)
);

NAND2xp5_ASAP7_75t_L g8639 ( 
.A(n_8608),
.B(n_8601),
.Y(n_8639)
);

NAND2xp5_ASAP7_75t_L g8640 ( 
.A(n_8606),
.B(n_6230),
.Y(n_8640)
);

OAI211xp5_ASAP7_75t_L g8641 ( 
.A1(n_8557),
.A2(n_6233),
.B(n_6235),
.C(n_6230),
.Y(n_8641)
);

OAI21xp5_ASAP7_75t_SL g8642 ( 
.A1(n_8626),
.A2(n_5768),
.B(n_6337),
.Y(n_8642)
);

NAND3xp33_ASAP7_75t_L g8643 ( 
.A(n_8549),
.B(n_6235),
.C(n_6233),
.Y(n_8643)
);

NOR2x1_ASAP7_75t_L g8644 ( 
.A(n_8574),
.B(n_6244),
.Y(n_8644)
);

INVx1_ASAP7_75t_L g8645 ( 
.A(n_8584),
.Y(n_8645)
);

NAND3xp33_ASAP7_75t_SL g8646 ( 
.A(n_8626),
.B(n_8553),
.C(n_8616),
.Y(n_8646)
);

OAI22xp5_ASAP7_75t_L g8647 ( 
.A1(n_8620),
.A2(n_6244),
.B1(n_6253),
.B2(n_6247),
.Y(n_8647)
);

NAND2xp5_ASAP7_75t_SL g8648 ( 
.A(n_8566),
.B(n_6247),
.Y(n_8648)
);

OAI22xp5_ASAP7_75t_L g8649 ( 
.A1(n_8590),
.A2(n_6258),
.B1(n_6283),
.B2(n_6259),
.Y(n_8649)
);

AOI21xp5_ASAP7_75t_L g8650 ( 
.A1(n_8562),
.A2(n_8541),
.B(n_8539),
.Y(n_8650)
);

INVx1_ASAP7_75t_L g8651 ( 
.A(n_8565),
.Y(n_8651)
);

NAND2xp5_ASAP7_75t_L g8652 ( 
.A(n_8537),
.B(n_6258),
.Y(n_8652)
);

AOI221xp5_ASAP7_75t_L g8653 ( 
.A1(n_8555),
.A2(n_6026),
.B1(n_6044),
.B2(n_6360),
.C(n_6352),
.Y(n_8653)
);

NAND2xp5_ASAP7_75t_SL g8654 ( 
.A(n_8595),
.B(n_6259),
.Y(n_8654)
);

OAI22xp33_ASAP7_75t_L g8655 ( 
.A1(n_8592),
.A2(n_6383),
.B1(n_6387),
.B2(n_6372),
.Y(n_8655)
);

OAI21xp33_ASAP7_75t_L g8656 ( 
.A1(n_8579),
.A2(n_6383),
.B(n_6372),
.Y(n_8656)
);

OAI211xp5_ASAP7_75t_L g8657 ( 
.A1(n_8591),
.A2(n_6283),
.B(n_6293),
.C(n_6286),
.Y(n_8657)
);

AOI221xp5_ASAP7_75t_L g8658 ( 
.A1(n_8609),
.A2(n_6026),
.B1(n_6388),
.B2(n_6395),
.C(n_6387),
.Y(n_8658)
);

OAI221xp5_ASAP7_75t_L g8659 ( 
.A1(n_8605),
.A2(n_6293),
.B1(n_6297),
.B2(n_6294),
.C(n_6286),
.Y(n_8659)
);

OAI22xp33_ASAP7_75t_L g8660 ( 
.A1(n_8563),
.A2(n_6395),
.B1(n_6297),
.B2(n_6302),
.Y(n_8660)
);

NAND2xp5_ASAP7_75t_SL g8661 ( 
.A(n_8561),
.B(n_6294),
.Y(n_8661)
);

NAND2xp33_ASAP7_75t_L g8662 ( 
.A(n_8597),
.B(n_6302),
.Y(n_8662)
);

OAI221xp5_ASAP7_75t_L g8663 ( 
.A1(n_8571),
.A2(n_6313),
.B1(n_6327),
.B2(n_6321),
.C(n_6308),
.Y(n_8663)
);

OAI311xp33_ASAP7_75t_L g8664 ( 
.A1(n_8585),
.A2(n_5726),
.A3(n_5805),
.B1(n_5802),
.C1(n_5722),
.Y(n_8664)
);

INVx2_ASAP7_75t_L g8665 ( 
.A(n_8538),
.Y(n_8665)
);

OAI221xp5_ASAP7_75t_SL g8666 ( 
.A1(n_8572),
.A2(n_5771),
.B1(n_6337),
.B2(n_6321),
.C(n_6313),
.Y(n_8666)
);

OAI221xp5_ASAP7_75t_SL g8667 ( 
.A1(n_8627),
.A2(n_6308),
.B1(n_6339),
.B2(n_6330),
.C(n_6327),
.Y(n_8667)
);

OAI21xp33_ASAP7_75t_L g8668 ( 
.A1(n_8544),
.A2(n_6339),
.B(n_6330),
.Y(n_8668)
);

AOI222xp33_ASAP7_75t_L g8669 ( 
.A1(n_8588),
.A2(n_6366),
.B1(n_6355),
.B2(n_6376),
.C1(n_6371),
.C2(n_6350),
.Y(n_8669)
);

NAND2xp5_ASAP7_75t_L g8670 ( 
.A(n_8551),
.B(n_6350),
.Y(n_8670)
);

AOI211xp5_ASAP7_75t_L g8671 ( 
.A1(n_8550),
.A2(n_6148),
.B(n_6366),
.C(n_6355),
.Y(n_8671)
);

INVx1_ASAP7_75t_SL g8672 ( 
.A(n_8542),
.Y(n_8672)
);

INVx1_ASAP7_75t_L g8673 ( 
.A(n_8578),
.Y(n_8673)
);

OAI222xp33_ASAP7_75t_L g8674 ( 
.A1(n_8598),
.A2(n_6325),
.B1(n_6377),
.B2(n_6378),
.C1(n_6376),
.C2(n_6371),
.Y(n_8674)
);

OAI222xp33_ASAP7_75t_L g8675 ( 
.A1(n_8589),
.A2(n_6325),
.B1(n_6380),
.B2(n_6389),
.C1(n_6378),
.C2(n_6377),
.Y(n_8675)
);

INVx1_ASAP7_75t_L g8676 ( 
.A(n_8621),
.Y(n_8676)
);

AOI221xp5_ASAP7_75t_L g8677 ( 
.A1(n_8558),
.A2(n_8564),
.B1(n_8581),
.B2(n_8596),
.C(n_8612),
.Y(n_8677)
);

AOI221xp5_ASAP7_75t_SL g8678 ( 
.A1(n_8613),
.A2(n_6389),
.B1(n_6380),
.B2(n_6342),
.C(n_5800),
.Y(n_8678)
);

INVxp67_ASAP7_75t_L g8679 ( 
.A(n_8604),
.Y(n_8679)
);

INVx2_ASAP7_75t_L g8680 ( 
.A(n_8619),
.Y(n_8680)
);

NAND2xp5_ASAP7_75t_L g8681 ( 
.A(n_8556),
.B(n_6363),
.Y(n_8681)
);

OAI221xp5_ASAP7_75t_L g8682 ( 
.A1(n_8546),
.A2(n_5710),
.B1(n_6186),
.B2(n_5992),
.C(n_5862),
.Y(n_8682)
);

A2O1A1Ixp33_ASAP7_75t_L g8683 ( 
.A1(n_8618),
.A2(n_6193),
.B(n_6214),
.C(n_6095),
.Y(n_8683)
);

OAI22xp5_ASAP7_75t_L g8684 ( 
.A1(n_8554),
.A2(n_8623),
.B1(n_8540),
.B2(n_8602),
.Y(n_8684)
);

AOI22xp33_ASAP7_75t_L g8685 ( 
.A1(n_8593),
.A2(n_6026),
.B1(n_6363),
.B2(n_6317),
.Y(n_8685)
);

AOI221xp5_ASAP7_75t_L g8686 ( 
.A1(n_8586),
.A2(n_6317),
.B1(n_6267),
.B2(n_6390),
.C(n_6263),
.Y(n_8686)
);

AOI211xp5_ASAP7_75t_L g8687 ( 
.A1(n_8625),
.A2(n_6214),
.B(n_5702),
.C(n_5819),
.Y(n_8687)
);

OAI211xp5_ASAP7_75t_L g8688 ( 
.A1(n_8615),
.A2(n_6186),
.B(n_6076),
.C(n_6005),
.Y(n_8688)
);

A2O1A1Ixp33_ASAP7_75t_SL g8689 ( 
.A1(n_8594),
.A2(n_5620),
.B(n_5627),
.C(n_5600),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8611),
.Y(n_8690)
);

OAI22xp5_ASAP7_75t_L g8691 ( 
.A1(n_8582),
.A2(n_6370),
.B1(n_6367),
.B2(n_6307),
.Y(n_8691)
);

INVx1_ASAP7_75t_L g8692 ( 
.A(n_8570),
.Y(n_8692)
);

INVx1_ASAP7_75t_L g8693 ( 
.A(n_8624),
.Y(n_8693)
);

INVx1_ASAP7_75t_L g8694 ( 
.A(n_8617),
.Y(n_8694)
);

XOR2x2_ASAP7_75t_SL g8695 ( 
.A(n_8573),
.B(n_5783),
.Y(n_8695)
);

AOI21xp5_ASAP7_75t_L g8696 ( 
.A1(n_8614),
.A2(n_6076),
.B(n_6101),
.Y(n_8696)
);

AOI21xp5_ASAP7_75t_L g8697 ( 
.A1(n_8575),
.A2(n_6076),
.B(n_6101),
.Y(n_8697)
);

AOI221xp5_ASAP7_75t_L g8698 ( 
.A1(n_8577),
.A2(n_6317),
.B1(n_6267),
.B2(n_6390),
.C(n_6263),
.Y(n_8698)
);

OAI22xp5_ASAP7_75t_L g8699 ( 
.A1(n_8622),
.A2(n_6370),
.B1(n_6367),
.B2(n_6307),
.Y(n_8699)
);

AND2x2_ASAP7_75t_L g8700 ( 
.A(n_8569),
.B(n_6342),
.Y(n_8700)
);

AOI221xp5_ASAP7_75t_L g8701 ( 
.A1(n_8559),
.A2(n_6267),
.B1(n_6390),
.B2(n_6263),
.C(n_5998),
.Y(n_8701)
);

O2A1O1Ixp33_ASAP7_75t_L g8702 ( 
.A1(n_8610),
.A2(n_6186),
.B(n_6114),
.C(n_6170),
.Y(n_8702)
);

INVx1_ASAP7_75t_L g8703 ( 
.A(n_8599),
.Y(n_8703)
);

AOI21xp33_ASAP7_75t_SL g8704 ( 
.A1(n_8607),
.A2(n_6095),
.B(n_6114),
.Y(n_8704)
);

CKINVDCx20_ASAP7_75t_R g8705 ( 
.A(n_8600),
.Y(n_8705)
);

OR2x2_ASAP7_75t_L g8706 ( 
.A(n_8568),
.B(n_6114),
.Y(n_8706)
);

NOR2xp33_ASAP7_75t_L g8707 ( 
.A(n_8568),
.B(n_6170),
.Y(n_8707)
);

OAI21xp33_ASAP7_75t_L g8708 ( 
.A1(n_8587),
.A2(n_6326),
.B(n_6232),
.Y(n_8708)
);

AOI222xp33_ASAP7_75t_L g8709 ( 
.A1(n_8588),
.A2(n_5627),
.B1(n_5637),
.B2(n_5650),
.C1(n_5645),
.C2(n_5634),
.Y(n_8709)
);

AOI221xp5_ASAP7_75t_L g8710 ( 
.A1(n_8555),
.A2(n_6170),
.B1(n_6109),
.B2(n_6107),
.C(n_6101),
.Y(n_8710)
);

OAI22xp5_ASAP7_75t_L g8711 ( 
.A1(n_8568),
.A2(n_6326),
.B1(n_6334),
.B2(n_6232),
.Y(n_8711)
);

NOR2xp33_ASAP7_75t_L g8712 ( 
.A(n_8568),
.B(n_6127),
.Y(n_8712)
);

OAI221xp5_ASAP7_75t_L g8713 ( 
.A1(n_8557),
.A2(n_6186),
.B1(n_5751),
.B2(n_5786),
.C(n_5795),
.Y(n_8713)
);

INVx1_ASAP7_75t_L g8714 ( 
.A(n_8583),
.Y(n_8714)
);

A2O1A1Ixp33_ASAP7_75t_L g8715 ( 
.A1(n_8595),
.A2(n_6334),
.B(n_5966),
.C(n_5969),
.Y(n_8715)
);

NOR4xp25_ASAP7_75t_L g8716 ( 
.A(n_8635),
.B(n_5637),
.C(n_5645),
.D(n_5634),
.Y(n_8716)
);

AOI221xp5_ASAP7_75t_L g8717 ( 
.A1(n_8631),
.A2(n_6109),
.B1(n_6107),
.B2(n_6202),
.C(n_6127),
.Y(n_8717)
);

NOR3xp33_ASAP7_75t_SL g8718 ( 
.A(n_8646),
.B(n_5967),
.C(n_5736),
.Y(n_8718)
);

AND3x2_ASAP7_75t_L g8719 ( 
.A(n_8632),
.B(n_5292),
.C(n_5287),
.Y(n_8719)
);

OAI321xp33_ASAP7_75t_L g8720 ( 
.A1(n_8712),
.A2(n_5976),
.A3(n_5979),
.B1(n_6013),
.B2(n_5861),
.C(n_5846),
.Y(n_8720)
);

OAI21xp33_ASAP7_75t_L g8721 ( 
.A1(n_8637),
.A2(n_5799),
.B(n_5787),
.Y(n_8721)
);

OAI211xp5_ASAP7_75t_SL g8722 ( 
.A1(n_8628),
.A2(n_8677),
.B(n_8629),
.C(n_8650),
.Y(n_8722)
);

AOI21xp33_ASAP7_75t_SL g8723 ( 
.A1(n_8706),
.A2(n_6127),
.B(n_6198),
.Y(n_8723)
);

AOI21xp5_ASAP7_75t_L g8724 ( 
.A1(n_8630),
.A2(n_6109),
.B(n_6107),
.Y(n_8724)
);

NAND4xp75_ASAP7_75t_L g8725 ( 
.A(n_8693),
.B(n_6198),
.C(n_6348),
.D(n_6329),
.Y(n_8725)
);

OAI21x1_ASAP7_75t_SL g8726 ( 
.A1(n_8636),
.A2(n_5966),
.B(n_5895),
.Y(n_8726)
);

NOR2x1_ASAP7_75t_L g8727 ( 
.A(n_8705),
.B(n_6202),
.Y(n_8727)
);

OAI21xp33_ASAP7_75t_SL g8728 ( 
.A1(n_8710),
.A2(n_8685),
.B(n_8707),
.Y(n_8728)
);

NAND2xp5_ASAP7_75t_L g8729 ( 
.A(n_8633),
.B(n_6202),
.Y(n_8729)
);

OAI322xp33_ASAP7_75t_L g8730 ( 
.A1(n_8679),
.A2(n_5969),
.A3(n_5650),
.B1(n_5729),
.B2(n_5673),
.C1(n_5749),
.C2(n_5687),
.Y(n_8730)
);

OAI21xp5_ASAP7_75t_L g8731 ( 
.A1(n_8672),
.A2(n_5644),
.B(n_6198),
.Y(n_8731)
);

AND2x2_ASAP7_75t_L g8732 ( 
.A(n_8665),
.B(n_6198),
.Y(n_8732)
);

OAI22xp5_ASAP7_75t_L g8733 ( 
.A1(n_8666),
.A2(n_5978),
.B1(n_5886),
.B2(n_5808),
.Y(n_8733)
);

AOI21xp5_ASAP7_75t_L g8734 ( 
.A1(n_8684),
.A2(n_8670),
.B(n_8681),
.Y(n_8734)
);

AOI22xp5_ASAP7_75t_L g8735 ( 
.A1(n_8708),
.A2(n_6329),
.B1(n_6348),
.B2(n_6358),
.Y(n_8735)
);

NOR4xp25_ASAP7_75t_L g8736 ( 
.A(n_8703),
.B(n_5673),
.C(n_5687),
.D(n_5671),
.Y(n_8736)
);

AOI222xp33_ASAP7_75t_L g8737 ( 
.A1(n_8658),
.A2(n_5770),
.B1(n_5671),
.B2(n_5772),
.C1(n_5749),
.C2(n_5729),
.Y(n_8737)
);

NAND2xp5_ASAP7_75t_L g8738 ( 
.A(n_8700),
.B(n_5961),
.Y(n_8738)
);

AND2x2_ASAP7_75t_L g8739 ( 
.A(n_8680),
.B(n_5313),
.Y(n_8739)
);

AOI222xp33_ASAP7_75t_L g8740 ( 
.A1(n_8654),
.A2(n_5797),
.B1(n_5772),
.B2(n_5813),
.C1(n_5809),
.C2(n_5770),
.Y(n_8740)
);

AOI22xp5_ASAP7_75t_L g8741 ( 
.A1(n_8692),
.A2(n_6329),
.B1(n_6348),
.B2(n_6358),
.Y(n_8741)
);

AOI21xp33_ASAP7_75t_L g8742 ( 
.A1(n_8684),
.A2(n_6348),
.B(n_6329),
.Y(n_8742)
);

OAI211xp5_ASAP7_75t_L g8743 ( 
.A1(n_8694),
.A2(n_6010),
.B(n_5999),
.C(n_5958),
.Y(n_8743)
);

AND2x2_ASAP7_75t_L g8744 ( 
.A(n_8651),
.B(n_5313),
.Y(n_8744)
);

O2A1O1Ixp33_ASAP7_75t_L g8745 ( 
.A1(n_8714),
.A2(n_5809),
.B(n_5813),
.C(n_5797),
.Y(n_8745)
);

AOI211xp5_ASAP7_75t_L g8746 ( 
.A1(n_8660),
.A2(n_5829),
.B(n_5863),
.C(n_5850),
.Y(n_8746)
);

AOI221xp5_ASAP7_75t_L g8747 ( 
.A1(n_8655),
.A2(n_5863),
.B1(n_5850),
.B2(n_5829),
.C(n_5959),
.Y(n_8747)
);

AOI221xp5_ASAP7_75t_L g8748 ( 
.A1(n_8674),
.A2(n_8638),
.B1(n_8656),
.B2(n_8668),
.C(n_8667),
.Y(n_8748)
);

OR2x2_ASAP7_75t_L g8749 ( 
.A(n_8711),
.B(n_6358),
.Y(n_8749)
);

OA211x2_ASAP7_75t_L g8750 ( 
.A1(n_8639),
.A2(n_5750),
.B(n_5950),
.C(n_5388),
.Y(n_8750)
);

A2O1A1Ixp33_ASAP7_75t_L g8751 ( 
.A1(n_8671),
.A2(n_5930),
.B(n_5927),
.C(n_5737),
.Y(n_8751)
);

NAND2xp5_ASAP7_75t_L g8752 ( 
.A(n_8678),
.B(n_6358),
.Y(n_8752)
);

AOI22xp5_ASAP7_75t_L g8753 ( 
.A1(n_8711),
.A2(n_6369),
.B1(n_6252),
.B2(n_6290),
.Y(n_8753)
);

NAND2xp5_ASAP7_75t_SL g8754 ( 
.A(n_8695),
.B(n_5898),
.Y(n_8754)
);

OAI211xp5_ASAP7_75t_L g8755 ( 
.A1(n_8676),
.A2(n_6369),
.B(n_5743),
.C(n_6252),
.Y(n_8755)
);

AOI22xp5_ASAP7_75t_L g8756 ( 
.A1(n_8642),
.A2(n_6369),
.B1(n_6252),
.B2(n_6290),
.Y(n_8756)
);

OR2x6_ASAP7_75t_L g8757 ( 
.A(n_8690),
.B(n_6369),
.Y(n_8757)
);

NAND2xp5_ASAP7_75t_L g8758 ( 
.A(n_8644),
.B(n_6252),
.Y(n_8758)
);

INVxp67_ASAP7_75t_L g8759 ( 
.A(n_8652),
.Y(n_8759)
);

AOI322xp5_ASAP7_75t_L g8760 ( 
.A1(n_8648),
.A2(n_8661),
.A3(n_8673),
.B1(n_8645),
.B2(n_8662),
.C1(n_8640),
.C2(n_8701),
.Y(n_8760)
);

O2A1O1Ixp33_ASAP7_75t_L g8761 ( 
.A1(n_8649),
.A2(n_6290),
.B(n_6270),
.C(n_5162),
.Y(n_8761)
);

NAND2xp5_ASAP7_75t_L g8762 ( 
.A(n_8657),
.B(n_6270),
.Y(n_8762)
);

AOI22xp5_ASAP7_75t_SL g8763 ( 
.A1(n_8634),
.A2(n_5380),
.B1(n_6290),
.B2(n_6270),
.Y(n_8763)
);

O2A1O1Ixp5_ASAP7_75t_SL g8764 ( 
.A1(n_8641),
.A2(n_6270),
.B(n_5225),
.C(n_5235),
.Y(n_8764)
);

OAI221xp5_ASAP7_75t_L g8765 ( 
.A1(n_8643),
.A2(n_5030),
.B1(n_5162),
.B2(n_5542),
.C(n_5539),
.Y(n_8765)
);

NOR3x1_ASAP7_75t_L g8766 ( 
.A(n_8689),
.B(n_5261),
.C(n_5546),
.Y(n_8766)
);

AOI221xp5_ASAP7_75t_L g8767 ( 
.A1(n_8647),
.A2(n_5544),
.B1(n_5411),
.B2(n_5225),
.C(n_5247),
.Y(n_8767)
);

NOR3x1_ASAP7_75t_L g8768 ( 
.A(n_8663),
.B(n_5261),
.C(n_5552),
.Y(n_8768)
);

NAND3xp33_ASAP7_75t_L g8769 ( 
.A(n_8697),
.B(n_5162),
.C(n_5030),
.Y(n_8769)
);

A2O1A1Ixp33_ASAP7_75t_L g8770 ( 
.A1(n_8702),
.A2(n_5084),
.B(n_5069),
.C(n_5226),
.Y(n_8770)
);

OAI21xp33_ASAP7_75t_L g8771 ( 
.A1(n_8704),
.A2(n_5410),
.B(n_5544),
.Y(n_8771)
);

AOI221xp5_ASAP7_75t_L g8772 ( 
.A1(n_8675),
.A2(n_5411),
.B1(n_5226),
.B2(n_5256),
.C(n_5247),
.Y(n_8772)
);

NAND2xp5_ASAP7_75t_L g8773 ( 
.A(n_8699),
.B(n_5254),
.Y(n_8773)
);

OAI221xp5_ASAP7_75t_L g8774 ( 
.A1(n_8659),
.A2(n_8715),
.B1(n_8682),
.B2(n_8691),
.C(n_8696),
.Y(n_8774)
);

OAI31xp33_ASAP7_75t_L g8775 ( 
.A1(n_8664),
.A2(n_5410),
.A3(n_5515),
.B(n_5533),
.Y(n_8775)
);

AOI21xp5_ASAP7_75t_L g8776 ( 
.A1(n_8686),
.A2(n_5272),
.B(n_5490),
.Y(n_8776)
);

NAND2xp5_ASAP7_75t_SL g8777 ( 
.A(n_8687),
.B(n_5533),
.Y(n_8777)
);

NOR3xp33_ASAP7_75t_L g8778 ( 
.A(n_8713),
.B(n_5412),
.C(n_5403),
.Y(n_8778)
);

NOR2xp33_ASAP7_75t_L g8779 ( 
.A(n_8688),
.B(n_5158),
.Y(n_8779)
);

AOI21xp5_ASAP7_75t_L g8780 ( 
.A1(n_8669),
.A2(n_5330),
.B(n_5363),
.Y(n_8780)
);

NAND3xp33_ASAP7_75t_L g8781 ( 
.A(n_8653),
.B(n_5363),
.C(n_5559),
.Y(n_8781)
);

NOR2xp67_ASAP7_75t_SL g8782 ( 
.A(n_8698),
.B(n_5537),
.Y(n_8782)
);

AOI211x1_ASAP7_75t_L g8783 ( 
.A1(n_8709),
.A2(n_5235),
.B(n_5266),
.C(n_5256),
.Y(n_8783)
);

NAND2xp5_ASAP7_75t_L g8784 ( 
.A(n_8716),
.B(n_8718),
.Y(n_8784)
);

OAI222xp33_ASAP7_75t_L g8785 ( 
.A1(n_8774),
.A2(n_8683),
.B1(n_5537),
.B2(n_5557),
.C1(n_5394),
.C2(n_5459),
.Y(n_8785)
);

OAI211xp5_ASAP7_75t_L g8786 ( 
.A1(n_8748),
.A2(n_8722),
.B(n_8760),
.C(n_8728),
.Y(n_8786)
);

OAI221xp5_ASAP7_75t_L g8787 ( 
.A1(n_8775),
.A2(n_5557),
.B1(n_5394),
.B2(n_5363),
.C(n_5270),
.Y(n_8787)
);

A2O1A1Ixp33_ASAP7_75t_L g8788 ( 
.A1(n_8724),
.A2(n_5084),
.B(n_5069),
.C(n_5266),
.Y(n_8788)
);

OAI32xp33_ASAP7_75t_L g8789 ( 
.A1(n_8729),
.A2(n_5459),
.A3(n_5453),
.B1(n_5425),
.B2(n_5418),
.Y(n_8789)
);

A2O1A1Ixp33_ASAP7_75t_L g8790 ( 
.A1(n_8779),
.A2(n_5270),
.B(n_5280),
.C(n_5268),
.Y(n_8790)
);

OAI211xp5_ASAP7_75t_SL g8791 ( 
.A1(n_8759),
.A2(n_5393),
.B(n_5375),
.C(n_5357),
.Y(n_8791)
);

AOI211xp5_ASAP7_75t_L g8792 ( 
.A1(n_8734),
.A2(n_5119),
.B(n_4899),
.C(n_5506),
.Y(n_8792)
);

OAI22xp5_ASAP7_75t_L g8793 ( 
.A1(n_8738),
.A2(n_5453),
.B1(n_5216),
.B2(n_5418),
.Y(n_8793)
);

AOI21xp33_ASAP7_75t_L g8794 ( 
.A1(n_8727),
.A2(n_5363),
.B(n_5553),
.Y(n_8794)
);

NOR3x1_ASAP7_75t_L g8795 ( 
.A(n_8777),
.B(n_5308),
.C(n_5119),
.Y(n_8795)
);

AOI22xp33_ASAP7_75t_L g8796 ( 
.A1(n_8778),
.A2(n_5330),
.B1(n_5553),
.B2(n_5316),
.Y(n_8796)
);

NAND2xp5_ASAP7_75t_L g8797 ( 
.A(n_8719),
.B(n_5254),
.Y(n_8797)
);

AND2x2_ASAP7_75t_L g8798 ( 
.A(n_8739),
.B(n_5081),
.Y(n_8798)
);

NAND2xp5_ASAP7_75t_L g8799 ( 
.A(n_8732),
.B(n_5262),
.Y(n_8799)
);

A2O1A1Ixp33_ASAP7_75t_L g8800 ( 
.A1(n_8771),
.A2(n_5280),
.B(n_5284),
.C(n_5268),
.Y(n_8800)
);

OAI221xp5_ASAP7_75t_L g8801 ( 
.A1(n_8770),
.A2(n_5296),
.B1(n_5299),
.B2(n_5295),
.C(n_5284),
.Y(n_8801)
);

NOR2xp33_ASAP7_75t_L g8802 ( 
.A(n_8773),
.B(n_5262),
.Y(n_8802)
);

INVx1_ASAP7_75t_L g8803 ( 
.A(n_8752),
.Y(n_8803)
);

OAI211xp5_ASAP7_75t_L g8804 ( 
.A1(n_8736),
.A2(n_5330),
.B(n_5316),
.C(n_5315),
.Y(n_8804)
);

NOR3xp33_ASAP7_75t_L g8805 ( 
.A(n_8754),
.B(n_5308),
.C(n_5127),
.Y(n_8805)
);

NAND2xp5_ASAP7_75t_L g8806 ( 
.A(n_8744),
.B(n_5264),
.Y(n_8806)
);

AOI21xp5_ASAP7_75t_L g8807 ( 
.A1(n_8758),
.A2(n_5330),
.B(n_5553),
.Y(n_8807)
);

OAI211xp5_ASAP7_75t_L g8808 ( 
.A1(n_8742),
.A2(n_5316),
.B(n_5315),
.C(n_5296),
.Y(n_8808)
);

INVxp67_ASAP7_75t_L g8809 ( 
.A(n_8782),
.Y(n_8809)
);

O2A1O1Ixp33_ASAP7_75t_SL g8810 ( 
.A1(n_8749),
.A2(n_5425),
.B(n_5407),
.C(n_5264),
.Y(n_8810)
);

OAI21xp33_ASAP7_75t_L g8811 ( 
.A1(n_8721),
.A2(n_5362),
.B(n_5342),
.Y(n_8811)
);

NAND4xp25_ASAP7_75t_SL g8812 ( 
.A(n_8762),
.B(n_5407),
.C(n_5515),
.D(n_5295),
.Y(n_8812)
);

OAI211xp5_ASAP7_75t_SL g8813 ( 
.A1(n_8731),
.A2(n_5548),
.B(n_5541),
.C(n_5477),
.Y(n_8813)
);

NAND2xp5_ASAP7_75t_L g8814 ( 
.A(n_8783),
.B(n_5275),
.Y(n_8814)
);

INVx1_ASAP7_75t_L g8815 ( 
.A(n_8726),
.Y(n_8815)
);

OAI211xp5_ASAP7_75t_L g8816 ( 
.A1(n_8781),
.A2(n_5316),
.B(n_5315),
.C(n_5299),
.Y(n_8816)
);

OAI211xp5_ASAP7_75t_SL g8817 ( 
.A1(n_8776),
.A2(n_5405),
.B(n_5317),
.C(n_5323),
.Y(n_8817)
);

NOR3x1_ASAP7_75t_L g8818 ( 
.A(n_8743),
.B(n_5326),
.C(n_5325),
.Y(n_8818)
);

AOI211xp5_ASAP7_75t_SL g8819 ( 
.A1(n_8720),
.A2(n_5317),
.B(n_5323),
.C(n_5314),
.Y(n_8819)
);

HB1xp67_ASAP7_75t_L g8820 ( 
.A(n_8766),
.Y(n_8820)
);

AOI21xp33_ASAP7_75t_L g8821 ( 
.A1(n_8763),
.A2(n_5553),
.B(n_5315),
.Y(n_8821)
);

NAND2xp5_ASAP7_75t_SL g8822 ( 
.A(n_8717),
.B(n_5275),
.Y(n_8822)
);

OR2x2_ASAP7_75t_L g8823 ( 
.A(n_8751),
.B(n_5302),
.Y(n_8823)
);

OAI211xp5_ASAP7_75t_L g8824 ( 
.A1(n_8772),
.A2(n_5314),
.B(n_5336),
.C(n_5333),
.Y(n_8824)
);

INVx1_ASAP7_75t_L g8825 ( 
.A(n_8745),
.Y(n_8825)
);

INVx1_ASAP7_75t_L g8826 ( 
.A(n_8750),
.Y(n_8826)
);

NOR4xp25_ASAP7_75t_L g8827 ( 
.A(n_8755),
.B(n_5336),
.C(n_5338),
.D(n_5333),
.Y(n_8827)
);

OAI21xp33_ASAP7_75t_SL g8828 ( 
.A1(n_8764),
.A2(n_5046),
.B(n_5043),
.Y(n_8828)
);

OAI221xp5_ASAP7_75t_L g8829 ( 
.A1(n_8746),
.A2(n_5341),
.B1(n_5346),
.B2(n_5339),
.C(n_5338),
.Y(n_8829)
);

OAI22xp5_ASAP7_75t_L g8830 ( 
.A1(n_8741),
.A2(n_8733),
.B1(n_8735),
.B2(n_8725),
.Y(n_8830)
);

AOI221xp5_ASAP7_75t_L g8831 ( 
.A1(n_8723),
.A2(n_5551),
.B1(n_5346),
.B2(n_5358),
.C(n_5341),
.Y(n_8831)
);

AOI21xp5_ASAP7_75t_L g8832 ( 
.A1(n_8769),
.A2(n_8780),
.B(n_8761),
.Y(n_8832)
);

AOI22xp5_ASAP7_75t_L g8833 ( 
.A1(n_8767),
.A2(n_5215),
.B1(n_5358),
.B2(n_5339),
.Y(n_8833)
);

OAI21xp5_ASAP7_75t_L g8834 ( 
.A1(n_8747),
.A2(n_5127),
.B(n_5253),
.Y(n_8834)
);

OAI21xp33_ASAP7_75t_L g8835 ( 
.A1(n_8756),
.A2(n_5081),
.B(n_5147),
.Y(n_8835)
);

INVx1_ASAP7_75t_L g8836 ( 
.A(n_8768),
.Y(n_8836)
);

AOI222xp33_ASAP7_75t_L g8837 ( 
.A1(n_8765),
.A2(n_5551),
.B1(n_5382),
.B2(n_5545),
.C1(n_5389),
.C2(n_5390),
.Y(n_8837)
);

OAI21xp33_ASAP7_75t_L g8838 ( 
.A1(n_8740),
.A2(n_5147),
.B(n_5146),
.Y(n_8838)
);

NAND2xp5_ASAP7_75t_SL g8839 ( 
.A(n_8826),
.B(n_8737),
.Y(n_8839)
);

NAND2xp5_ASAP7_75t_L g8840 ( 
.A(n_8820),
.B(n_8753),
.Y(n_8840)
);

NAND2xp5_ASAP7_75t_L g8841 ( 
.A(n_8809),
.B(n_8757),
.Y(n_8841)
);

NAND4xp25_ASAP7_75t_L g8842 ( 
.A(n_8786),
.B(n_8730),
.C(n_8757),
.D(n_4891),
.Y(n_8842)
);

AOI211xp5_ASAP7_75t_L g8843 ( 
.A1(n_8830),
.A2(n_8757),
.B(n_5377),
.C(n_5382),
.Y(n_8843)
);

NAND2xp5_ASAP7_75t_L g8844 ( 
.A(n_8803),
.B(n_5302),
.Y(n_8844)
);

NAND4xp25_ASAP7_75t_L g8845 ( 
.A(n_8784),
.B(n_4891),
.C(n_5377),
.D(n_5373),
.Y(n_8845)
);

INVx2_ASAP7_75t_L g8846 ( 
.A(n_8823),
.Y(n_8846)
);

NAND4xp25_ASAP7_75t_L g8847 ( 
.A(n_8819),
.B(n_5385),
.C(n_5389),
.D(n_5373),
.Y(n_8847)
);

NOR3xp33_ASAP7_75t_SL g8848 ( 
.A(n_8836),
.B(n_5390),
.C(n_5385),
.Y(n_8848)
);

OAI22xp33_ASAP7_75t_L g8849 ( 
.A1(n_8797),
.A2(n_8787),
.B1(n_8825),
.B2(n_8815),
.Y(n_8849)
);

NOR2xp33_ASAP7_75t_SL g8850 ( 
.A(n_8785),
.B(n_5391),
.Y(n_8850)
);

A2O1A1Ixp33_ASAP7_75t_L g8851 ( 
.A1(n_8832),
.A2(n_5396),
.B(n_5397),
.C(n_5395),
.Y(n_8851)
);

NOR3x1_ASAP7_75t_L g8852 ( 
.A(n_8822),
.B(n_5326),
.C(n_5325),
.Y(n_8852)
);

AOI221xp5_ASAP7_75t_L g8853 ( 
.A1(n_8827),
.A2(n_5397),
.B1(n_5404),
.B2(n_5396),
.C(n_5395),
.Y(n_8853)
);

AND2x2_ASAP7_75t_L g8854 ( 
.A(n_8798),
.B(n_8790),
.Y(n_8854)
);

NAND3xp33_ASAP7_75t_SL g8855 ( 
.A(n_8805),
.B(n_5406),
.C(n_5404),
.Y(n_8855)
);

OAI221xp5_ASAP7_75t_L g8856 ( 
.A1(n_8799),
.A2(n_5409),
.B1(n_5413),
.B2(n_5408),
.C(n_5406),
.Y(n_8856)
);

NOR3xp33_ASAP7_75t_L g8857 ( 
.A(n_8802),
.B(n_5046),
.C(n_5043),
.Y(n_8857)
);

NAND2xp5_ASAP7_75t_L g8858 ( 
.A(n_8814),
.B(n_5320),
.Y(n_8858)
);

OAI211xp5_ASAP7_75t_SL g8859 ( 
.A1(n_8837),
.A2(n_5409),
.B(n_5413),
.C(n_5408),
.Y(n_8859)
);

NAND5xp2_ASAP7_75t_L g8860 ( 
.A(n_8831),
.B(n_5500),
.C(n_5549),
.D(n_5430),
.E(n_5432),
.Y(n_8860)
);

AOI211xp5_ASAP7_75t_L g8861 ( 
.A1(n_8812),
.A2(n_5419),
.B(n_5430),
.C(n_5428),
.Y(n_8861)
);

NAND3xp33_ASAP7_75t_L g8862 ( 
.A(n_8816),
.B(n_5428),
.C(n_5419),
.Y(n_8862)
);

NOR2xp33_ASAP7_75t_L g8863 ( 
.A(n_8806),
.B(n_5320),
.Y(n_8863)
);

AOI211xp5_ASAP7_75t_L g8864 ( 
.A1(n_8810),
.A2(n_8801),
.B(n_8817),
.C(n_8808),
.Y(n_8864)
);

INVx2_ASAP7_75t_L g8865 ( 
.A(n_8818),
.Y(n_8865)
);

NOR2xp33_ASAP7_75t_L g8866 ( 
.A(n_8838),
.B(n_5345),
.Y(n_8866)
);

NAND3xp33_ASAP7_75t_SL g8867 ( 
.A(n_8833),
.B(n_5433),
.C(n_5432),
.Y(n_8867)
);

NOR2xp67_ASAP7_75t_L g8868 ( 
.A(n_8828),
.B(n_5345),
.Y(n_8868)
);

NOR2x1_ASAP7_75t_L g8869 ( 
.A(n_8800),
.B(n_5215),
.Y(n_8869)
);

NAND2xp5_ASAP7_75t_L g8870 ( 
.A(n_8835),
.B(n_5347),
.Y(n_8870)
);

NAND2xp5_ASAP7_75t_SL g8871 ( 
.A(n_8792),
.B(n_5347),
.Y(n_8871)
);

INVx2_ASAP7_75t_SL g8872 ( 
.A(n_8793),
.Y(n_8872)
);

NAND4xp25_ASAP7_75t_L g8873 ( 
.A(n_8795),
.B(n_5434),
.C(n_5435),
.D(n_5433),
.Y(n_8873)
);

NAND2xp5_ASAP7_75t_L g8874 ( 
.A(n_8824),
.B(n_5374),
.Y(n_8874)
);

NAND2x1_ASAP7_75t_SL g8875 ( 
.A(n_8788),
.B(n_5374),
.Y(n_8875)
);

NAND4xp25_ASAP7_75t_SL g8876 ( 
.A(n_8807),
.B(n_5435),
.C(n_5436),
.D(n_5434),
.Y(n_8876)
);

NOR2x1_ASAP7_75t_L g8877 ( 
.A(n_8829),
.B(n_5215),
.Y(n_8877)
);

NOR2x1_ASAP7_75t_L g8878 ( 
.A(n_8813),
.B(n_5436),
.Y(n_8878)
);

NAND4xp25_ASAP7_75t_L g8879 ( 
.A(n_8811),
.B(n_5454),
.C(n_5462),
.D(n_5442),
.Y(n_8879)
);

NAND4xp75_ASAP7_75t_L g8880 ( 
.A(n_8834),
.B(n_5274),
.C(n_5293),
.D(n_5228),
.Y(n_8880)
);

INVx1_ASAP7_75t_L g8881 ( 
.A(n_8789),
.Y(n_8881)
);

NAND4xp25_ASAP7_75t_L g8882 ( 
.A(n_8843),
.B(n_8791),
.C(n_8794),
.D(n_8821),
.Y(n_8882)
);

OAI211xp5_ASAP7_75t_L g8883 ( 
.A1(n_8839),
.A2(n_8840),
.B(n_8841),
.C(n_8881),
.Y(n_8883)
);

NAND2xp5_ASAP7_75t_L g8884 ( 
.A(n_8865),
.B(n_8821),
.Y(n_8884)
);

NAND3xp33_ASAP7_75t_SL g8885 ( 
.A(n_8846),
.B(n_8796),
.C(n_8804),
.Y(n_8885)
);

NAND4xp25_ASAP7_75t_L g8886 ( 
.A(n_8842),
.B(n_5454),
.C(n_5462),
.D(n_5442),
.Y(n_8886)
);

OAI211xp5_ASAP7_75t_L g8887 ( 
.A1(n_8842),
.A2(n_5465),
.B(n_5474),
.C(n_5464),
.Y(n_8887)
);

NOR2xp67_ASAP7_75t_L g8888 ( 
.A(n_8872),
.B(n_5400),
.Y(n_8888)
);

NAND2xp5_ASAP7_75t_L g8889 ( 
.A(n_8868),
.B(n_5400),
.Y(n_8889)
);

INVx1_ASAP7_75t_SL g8890 ( 
.A(n_8854),
.Y(n_8890)
);

OAI211xp5_ASAP7_75t_SL g8891 ( 
.A1(n_8849),
.A2(n_5465),
.B(n_5474),
.C(n_5464),
.Y(n_8891)
);

OAI211xp5_ASAP7_75t_SL g8892 ( 
.A1(n_8864),
.A2(n_5496),
.B(n_5498),
.C(n_5483),
.Y(n_8892)
);

NOR3xp33_ASAP7_75t_L g8893 ( 
.A(n_8844),
.B(n_5257),
.C(n_4569),
.Y(n_8893)
);

AOI221xp5_ASAP7_75t_L g8894 ( 
.A1(n_8866),
.A2(n_5498),
.B1(n_5496),
.B2(n_5483),
.C(n_5528),
.Y(n_8894)
);

INVxp67_ASAP7_75t_SL g8895 ( 
.A(n_8858),
.Y(n_8895)
);

NAND3xp33_ASAP7_75t_L g8896 ( 
.A(n_8848),
.B(n_8850),
.C(n_8873),
.Y(n_8896)
);

AOI211xp5_ASAP7_75t_SL g8897 ( 
.A1(n_8870),
.A2(n_5545),
.B(n_5528),
.C(n_5427),
.Y(n_8897)
);

NOR4xp25_ASAP7_75t_L g8898 ( 
.A(n_8867),
.B(n_5427),
.C(n_5469),
.D(n_5424),
.Y(n_8898)
);

OAI221xp5_ASAP7_75t_L g8899 ( 
.A1(n_8874),
.A2(n_8875),
.B1(n_8851),
.B2(n_8869),
.C(n_8847),
.Y(n_8899)
);

XNOR2x1_ASAP7_75t_L g8900 ( 
.A(n_8878),
.B(n_5391),
.Y(n_8900)
);

NAND4xp25_ASAP7_75t_L g8901 ( 
.A(n_8863),
.B(n_5469),
.C(n_5471),
.D(n_5424),
.Y(n_8901)
);

INVxp33_ASAP7_75t_L g8902 ( 
.A(n_8877),
.Y(n_8902)
);

INVx1_ASAP7_75t_L g8903 ( 
.A(n_8855),
.Y(n_8903)
);

AOI221xp5_ASAP7_75t_L g8904 ( 
.A1(n_8871),
.A2(n_5471),
.B1(n_5473),
.B2(n_5529),
.C(n_5493),
.Y(n_8904)
);

NOR2x1p5_ASAP7_75t_L g8905 ( 
.A(n_8879),
.B(n_5473),
.Y(n_8905)
);

NOR3xp33_ASAP7_75t_L g8906 ( 
.A(n_8876),
.B(n_8859),
.C(n_8860),
.Y(n_8906)
);

NAND3xp33_ASAP7_75t_SL g8907 ( 
.A(n_8861),
.B(n_8862),
.C(n_8853),
.Y(n_8907)
);

NOR2x1p5_ASAP7_75t_L g8908 ( 
.A(n_8845),
.B(n_5493),
.Y(n_8908)
);

NAND3xp33_ASAP7_75t_L g8909 ( 
.A(n_8856),
.B(n_5511),
.C(n_5495),
.Y(n_8909)
);

AOI22xp5_ASAP7_75t_L g8910 ( 
.A1(n_8880),
.A2(n_5511),
.B1(n_5527),
.B2(n_5495),
.Y(n_8910)
);

AOI211x1_ASAP7_75t_L g8911 ( 
.A1(n_8852),
.A2(n_5500),
.B(n_5549),
.C(n_5146),
.Y(n_8911)
);

NAND4xp75_ASAP7_75t_L g8912 ( 
.A(n_8857),
.B(n_5274),
.C(n_5293),
.D(n_5228),
.Y(n_8912)
);

OAI221xp5_ASAP7_75t_L g8913 ( 
.A1(n_8842),
.A2(n_5529),
.B1(n_5527),
.B2(n_5391),
.C(n_5274),
.Y(n_8913)
);

AOI21xp5_ASAP7_75t_L g8914 ( 
.A1(n_8841),
.A2(n_5206),
.B(n_5179),
.Y(n_8914)
);

NAND4xp75_ASAP7_75t_L g8915 ( 
.A(n_8839),
.B(n_5274),
.C(n_5293),
.D(n_5228),
.Y(n_8915)
);

OAI21xp5_ASAP7_75t_L g8916 ( 
.A1(n_8839),
.A2(n_5257),
.B(n_4564),
.Y(n_8916)
);

AOI21xp5_ASAP7_75t_L g8917 ( 
.A1(n_8841),
.A2(n_5206),
.B(n_5179),
.Y(n_8917)
);

NOR3xp33_ASAP7_75t_L g8918 ( 
.A(n_8849),
.B(n_4569),
.C(n_5136),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_8841),
.Y(n_8919)
);

AOI211xp5_ASAP7_75t_L g8920 ( 
.A1(n_8849),
.A2(n_5516),
.B(n_5523),
.C(n_5518),
.Y(n_8920)
);

AND2x2_ASAP7_75t_SL g8921 ( 
.A(n_8919),
.B(n_5234),
.Y(n_8921)
);

NOR2x1_ASAP7_75t_SL g8922 ( 
.A(n_8883),
.B(n_5391),
.Y(n_8922)
);

INVx1_ASAP7_75t_L g8923 ( 
.A(n_8888),
.Y(n_8923)
);

AOI22xp5_ASAP7_75t_L g8924 ( 
.A1(n_8890),
.A2(n_5111),
.B1(n_5206),
.B2(n_5293),
.Y(n_8924)
);

NOR2x1_ASAP7_75t_L g8925 ( 
.A(n_8903),
.B(n_5111),
.Y(n_8925)
);

AND3x4_ASAP7_75t_L g8926 ( 
.A(n_8906),
.B(n_4649),
.C(n_4634),
.Y(n_8926)
);

NOR2x1_ASAP7_75t_L g8927 ( 
.A(n_8884),
.B(n_8896),
.Y(n_8927)
);

AOI22xp5_ASAP7_75t_L g8928 ( 
.A1(n_8895),
.A2(n_5228),
.B1(n_4529),
.B2(n_5234),
.Y(n_8928)
);

AOI22xp5_ASAP7_75t_L g8929 ( 
.A1(n_8886),
.A2(n_4529),
.B1(n_5234),
.B2(n_5236),
.Y(n_8929)
);

AO22x2_ASAP7_75t_L g8930 ( 
.A1(n_8885),
.A2(n_4933),
.B1(n_4934),
.B2(n_4907),
.Y(n_8930)
);

AND2x2_ASAP7_75t_L g8931 ( 
.A(n_8900),
.B(n_5234),
.Y(n_8931)
);

OR2x2_ASAP7_75t_L g8932 ( 
.A(n_8889),
.B(n_5307),
.Y(n_8932)
);

INVx2_ASAP7_75t_L g8933 ( 
.A(n_8908),
.Y(n_8933)
);

NOR2x1_ASAP7_75t_L g8934 ( 
.A(n_8899),
.B(n_5502),
.Y(n_8934)
);

AND2x4_ASAP7_75t_L g8935 ( 
.A(n_8905),
.B(n_4758),
.Y(n_8935)
);

INVxp33_ASAP7_75t_SL g8936 ( 
.A(n_8902),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_8891),
.Y(n_8937)
);

AOI22xp5_ASAP7_75t_L g8938 ( 
.A1(n_8918),
.A2(n_4529),
.B1(n_5236),
.B2(n_5502),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_8887),
.Y(n_8939)
);

NOR2x1_ASAP7_75t_L g8940 ( 
.A(n_8907),
.B(n_5517),
.Y(n_8940)
);

INVx3_ASAP7_75t_L g8941 ( 
.A(n_8892),
.Y(n_8941)
);

AOI221xp5_ASAP7_75t_L g8942 ( 
.A1(n_8882),
.A2(n_8913),
.B1(n_8898),
.B2(n_8911),
.C(n_8920),
.Y(n_8942)
);

AOI22xp5_ASAP7_75t_L g8943 ( 
.A1(n_8909),
.A2(n_5236),
.B1(n_5517),
.B2(n_5519),
.Y(n_8943)
);

NOR2x1_ASAP7_75t_L g8944 ( 
.A(n_8915),
.B(n_5532),
.Y(n_8944)
);

AOI22xp33_ASAP7_75t_SL g8945 ( 
.A1(n_8916),
.A2(n_5236),
.B1(n_5514),
.B2(n_5504),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8910),
.Y(n_8946)
);

OR2x2_ASAP7_75t_L g8947 ( 
.A(n_8901),
.B(n_5307),
.Y(n_8947)
);

NOR2x1_ASAP7_75t_L g8948 ( 
.A(n_8912),
.B(n_5532),
.Y(n_8948)
);

NOR2x1_ASAP7_75t_L g8949 ( 
.A(n_8923),
.B(n_8914),
.Y(n_8949)
);

NOR4xp25_ASAP7_75t_SL g8950 ( 
.A(n_8939),
.B(n_8904),
.C(n_8894),
.D(n_8897),
.Y(n_8950)
);

NOR2x1_ASAP7_75t_L g8951 ( 
.A(n_8927),
.B(n_8946),
.Y(n_8951)
);

AND2x4_ASAP7_75t_L g8952 ( 
.A(n_8925),
.B(n_8893),
.Y(n_8952)
);

NAND4xp75_ASAP7_75t_L g8953 ( 
.A(n_8933),
.B(n_8917),
.C(n_5514),
.D(n_5504),
.Y(n_8953)
);

AOI211xp5_ASAP7_75t_L g8954 ( 
.A1(n_8942),
.A2(n_5518),
.B(n_5523),
.C(n_5516),
.Y(n_8954)
);

NOR3xp33_ASAP7_75t_L g8955 ( 
.A(n_8941),
.B(n_4569),
.C(n_5136),
.Y(n_8955)
);

INVxp67_ASAP7_75t_L g8956 ( 
.A(n_8937),
.Y(n_8956)
);

NAND3xp33_ASAP7_75t_L g8957 ( 
.A(n_8940),
.B(n_8934),
.C(n_8948),
.Y(n_8957)
);

NAND4xp75_ASAP7_75t_L g8958 ( 
.A(n_8936),
.B(n_5514),
.C(n_5504),
.D(n_5361),
.Y(n_8958)
);

AND2x4_ASAP7_75t_L g8959 ( 
.A(n_8922),
.B(n_4758),
.Y(n_8959)
);

INVx1_ASAP7_75t_L g8960 ( 
.A(n_8930),
.Y(n_8960)
);

AND2x4_ASAP7_75t_L g8961 ( 
.A(n_8931),
.B(n_4758),
.Y(n_8961)
);

NOR3xp33_ASAP7_75t_L g8962 ( 
.A(n_8944),
.B(n_5137),
.C(n_4564),
.Y(n_8962)
);

NOR4xp25_ASAP7_75t_L g8963 ( 
.A(n_8932),
.B(n_4934),
.C(n_4951),
.D(n_4933),
.Y(n_8963)
);

NAND2xp5_ASAP7_75t_L g8964 ( 
.A(n_8930),
.B(n_5307),
.Y(n_8964)
);

NOR3xp33_ASAP7_75t_L g8965 ( 
.A(n_8947),
.B(n_5137),
.C(n_4564),
.Y(n_8965)
);

NAND2xp5_ASAP7_75t_L g8966 ( 
.A(n_8935),
.B(n_5307),
.Y(n_8966)
);

NOR3xp33_ASAP7_75t_L g8967 ( 
.A(n_8926),
.B(n_8938),
.C(n_8929),
.Y(n_8967)
);

NOR2xp67_ASAP7_75t_L g8968 ( 
.A(n_8943),
.B(n_4966),
.Y(n_8968)
);

NOR3xp33_ASAP7_75t_L g8969 ( 
.A(n_8945),
.B(n_4602),
.C(n_4559),
.Y(n_8969)
);

NAND2xp5_ASAP7_75t_L g8970 ( 
.A(n_8951),
.B(n_8921),
.Y(n_8970)
);

CKINVDCx5p33_ASAP7_75t_R g8971 ( 
.A(n_8956),
.Y(n_8971)
);

NOR3xp33_ASAP7_75t_L g8972 ( 
.A(n_8949),
.B(n_8924),
.C(n_8928),
.Y(n_8972)
);

NOR2x1_ASAP7_75t_L g8973 ( 
.A(n_8957),
.B(n_5532),
.Y(n_8973)
);

OAI211xp5_ASAP7_75t_SL g8974 ( 
.A1(n_8960),
.A2(n_4976),
.B(n_4978),
.C(n_4974),
.Y(n_8974)
);

OR2x2_ASAP7_75t_L g8975 ( 
.A(n_8959),
.B(n_5307),
.Y(n_8975)
);

INVx1_ASAP7_75t_L g8976 ( 
.A(n_8952),
.Y(n_8976)
);

INVxp67_ASAP7_75t_L g8977 ( 
.A(n_8952),
.Y(n_8977)
);

INVxp33_ASAP7_75t_L g8978 ( 
.A(n_8967),
.Y(n_8978)
);

NOR3xp33_ASAP7_75t_L g8979 ( 
.A(n_8965),
.B(n_4559),
.C(n_4602),
.Y(n_8979)
);

OAI221xp5_ASAP7_75t_L g8980 ( 
.A1(n_8962),
.A2(n_5190),
.B1(n_5514),
.B2(n_5504),
.C(n_5484),
.Y(n_8980)
);

AOI221xp5_ASAP7_75t_L g8981 ( 
.A1(n_8963),
.A2(n_4978),
.B1(n_4976),
.B2(n_5519),
.C(n_5536),
.Y(n_8981)
);

INVx1_ASAP7_75t_L g8982 ( 
.A(n_8968),
.Y(n_8982)
);

NAND4xp75_ASAP7_75t_L g8983 ( 
.A(n_8950),
.B(n_5361),
.C(n_5484),
.D(n_5456),
.Y(n_8983)
);

AO22x1_ASAP7_75t_L g8984 ( 
.A1(n_8969),
.A2(n_4667),
.B1(n_4703),
.B2(n_4649),
.Y(n_8984)
);

NOR3xp33_ASAP7_75t_L g8985 ( 
.A(n_8953),
.B(n_4559),
.C(n_5171),
.Y(n_8985)
);

INVxp33_ASAP7_75t_L g8986 ( 
.A(n_8966),
.Y(n_8986)
);

NAND4xp75_ASAP7_75t_L g8987 ( 
.A(n_8964),
.B(n_5484),
.C(n_5456),
.D(n_5361),
.Y(n_8987)
);

AND2x2_ASAP7_75t_SL g8988 ( 
.A(n_8976),
.B(n_8955),
.Y(n_8988)
);

XOR2x1_ASAP7_75t_L g8989 ( 
.A(n_8982),
.B(n_8961),
.Y(n_8989)
);

OR2x6_ASAP7_75t_L g8990 ( 
.A(n_8970),
.B(n_8961),
.Y(n_8990)
);

INVx2_ASAP7_75t_L g8991 ( 
.A(n_8971),
.Y(n_8991)
);

NAND3x1_ASAP7_75t_L g8992 ( 
.A(n_8972),
.B(n_8954),
.C(n_8958),
.Y(n_8992)
);

INVx1_ASAP7_75t_L g8993 ( 
.A(n_8977),
.Y(n_8993)
);

AND2x4_ASAP7_75t_L g8994 ( 
.A(n_8975),
.B(n_4758),
.Y(n_8994)
);

CKINVDCx14_ASAP7_75t_R g8995 ( 
.A(n_8978),
.Y(n_8995)
);

INVx1_ASAP7_75t_L g8996 ( 
.A(n_8973),
.Y(n_8996)
);

NOR3xp33_ASAP7_75t_L g8997 ( 
.A(n_8986),
.B(n_5204),
.C(n_5171),
.Y(n_8997)
);

INVx3_ASAP7_75t_L g8998 ( 
.A(n_8983),
.Y(n_8998)
);

HB1xp67_ASAP7_75t_L g8999 ( 
.A(n_8985),
.Y(n_8999)
);

OR2x2_ASAP7_75t_L g9000 ( 
.A(n_8984),
.B(n_5352),
.Y(n_9000)
);

AND2x4_ASAP7_75t_L g9001 ( 
.A(n_8979),
.B(n_4758),
.Y(n_9001)
);

NOR3xp33_ASAP7_75t_SL g9002 ( 
.A(n_8974),
.B(n_4607),
.C(n_4658),
.Y(n_9002)
);

AND4x1_ASAP7_75t_L g9003 ( 
.A(n_8981),
.B(n_4607),
.C(n_5352),
.D(n_4658),
.Y(n_9003)
);

NOR2x1_ASAP7_75t_L g9004 ( 
.A(n_8987),
.B(n_8980),
.Y(n_9004)
);

NOR3xp33_ASAP7_75t_L g9005 ( 
.A(n_8977),
.B(n_5204),
.C(n_4594),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8993),
.Y(n_9006)
);

INVx3_ASAP7_75t_SL g9007 ( 
.A(n_8990),
.Y(n_9007)
);

INVx2_ASAP7_75t_L g9008 ( 
.A(n_8989),
.Y(n_9008)
);

CKINVDCx20_ASAP7_75t_R g9009 ( 
.A(n_8995),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8999),
.Y(n_9010)
);

HB1xp67_ASAP7_75t_L g9011 ( 
.A(n_8990),
.Y(n_9011)
);

INVx2_ASAP7_75t_L g9012 ( 
.A(n_8998),
.Y(n_9012)
);

AND2x2_ASAP7_75t_L g9013 ( 
.A(n_8991),
.B(n_5190),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_8988),
.Y(n_9014)
);

INVx1_ASAP7_75t_L g9015 ( 
.A(n_8992),
.Y(n_9015)
);

INVx1_ASAP7_75t_L g9016 ( 
.A(n_9004),
.Y(n_9016)
);

INVx2_ASAP7_75t_L g9017 ( 
.A(n_8996),
.Y(n_9017)
);

AND3x4_ASAP7_75t_L g9018 ( 
.A(n_9001),
.B(n_4667),
.C(n_4649),
.Y(n_9018)
);

OAI22xp5_ASAP7_75t_L g9019 ( 
.A1(n_9000),
.A2(n_5484),
.B1(n_5456),
.B2(n_5361),
.Y(n_9019)
);

XOR2x1_ASAP7_75t_L g9020 ( 
.A(n_9011),
.B(n_8994),
.Y(n_9020)
);

INVxp67_ASAP7_75t_SL g9021 ( 
.A(n_9008),
.Y(n_9021)
);

INVx1_ASAP7_75t_L g9022 ( 
.A(n_9006),
.Y(n_9022)
);

INVx4_ASAP7_75t_L g9023 ( 
.A(n_9007),
.Y(n_9023)
);

AND2x2_ASAP7_75t_SL g9024 ( 
.A(n_9012),
.B(n_8997),
.Y(n_9024)
);

INVx2_ASAP7_75t_L g9025 ( 
.A(n_9009),
.Y(n_9025)
);

HB1xp67_ASAP7_75t_L g9026 ( 
.A(n_9016),
.Y(n_9026)
);

AND2x2_ASAP7_75t_L g9027 ( 
.A(n_9017),
.B(n_9002),
.Y(n_9027)
);

NOR2x1p5_ASAP7_75t_L g9028 ( 
.A(n_9014),
.B(n_9015),
.Y(n_9028)
);

HB1xp67_ASAP7_75t_L g9029 ( 
.A(n_9010),
.Y(n_9029)
);

INVx2_ASAP7_75t_SL g9030 ( 
.A(n_9028),
.Y(n_9030)
);

NAND2xp5_ASAP7_75t_L g9031 ( 
.A(n_9026),
.B(n_9013),
.Y(n_9031)
);

AOI221xp5_ASAP7_75t_L g9032 ( 
.A1(n_9021),
.A2(n_9019),
.B1(n_9018),
.B2(n_9005),
.C(n_9003),
.Y(n_9032)
);

CKINVDCx5p33_ASAP7_75t_R g9033 ( 
.A(n_9029),
.Y(n_9033)
);

HB1xp67_ASAP7_75t_L g9034 ( 
.A(n_9033),
.Y(n_9034)
);

NAND3xp33_ASAP7_75t_L g9035 ( 
.A(n_9030),
.B(n_9023),
.C(n_9025),
.Y(n_9035)
);

HB1xp67_ASAP7_75t_L g9036 ( 
.A(n_9031),
.Y(n_9036)
);

NAND2xp5_ASAP7_75t_L g9037 ( 
.A(n_9032),
.B(n_9022),
.Y(n_9037)
);

INVx1_ASAP7_75t_L g9038 ( 
.A(n_9035),
.Y(n_9038)
);

INVx1_ASAP7_75t_L g9039 ( 
.A(n_9034),
.Y(n_9039)
);

AOI21xp5_ASAP7_75t_L g9040 ( 
.A1(n_9037),
.A2(n_9024),
.B(n_9027),
.Y(n_9040)
);

HB1xp67_ASAP7_75t_L g9041 ( 
.A(n_9038),
.Y(n_9041)
);

OAI22x1_ASAP7_75t_L g9042 ( 
.A1(n_9041),
.A2(n_9039),
.B1(n_9036),
.B2(n_9020),
.Y(n_9042)
);

AOI221xp5_ASAP7_75t_L g9043 ( 
.A1(n_9042),
.A2(n_9040),
.B1(n_5536),
.B2(n_5519),
.C(n_4999),
.Y(n_9043)
);

OAI222xp33_ASAP7_75t_L g9044 ( 
.A1(n_9043),
.A2(n_4732),
.B1(n_4667),
.B2(n_4703),
.C1(n_4714),
.C2(n_4724),
.Y(n_9044)
);

OAI21xp5_ASAP7_75t_L g9045 ( 
.A1(n_9044),
.A2(n_5335),
.B(n_4691),
.Y(n_9045)
);

INVx1_ASAP7_75t_L g9046 ( 
.A(n_9045),
.Y(n_9046)
);

AO21x2_ASAP7_75t_L g9047 ( 
.A1(n_9046),
.A2(n_4594),
.B(n_5535),
.Y(n_9047)
);

OAI21xp5_ASAP7_75t_L g9048 ( 
.A1(n_9046),
.A2(n_4691),
.B(n_4668),
.Y(n_9048)
);

OAI221xp5_ASAP7_75t_R g9049 ( 
.A1(n_9048),
.A2(n_9047),
.B1(n_5352),
.B2(n_4607),
.C(n_5536),
.Y(n_9049)
);

AOI22xp5_ASAP7_75t_L g9050 ( 
.A1(n_9049),
.A2(n_2540),
.B1(n_2549),
.B2(n_2551),
.Y(n_9050)
);

AOI211xp5_ASAP7_75t_L g9051 ( 
.A1(n_9050),
.A2(n_2540),
.B(n_2549),
.C(n_2551),
.Y(n_9051)
);


endmodule