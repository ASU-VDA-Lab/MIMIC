module real_jpeg_15237_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_27;
wire n_32;
wire n_20;
wire n_19;
wire n_26;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AO22x1_ASAP7_75t_SL g11 ( 
.A1(n_0),
.A2(n_1),
.B1(n_12),
.B2(n_13),
.Y(n_11)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

OA22x2_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_4),
.B1(n_13),
.B2(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx2_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

OR2x4_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_16),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_16),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_3),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

AOI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_14),
.B(n_23),
.C(n_32),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_10),
.Y(n_8)
);

OR2x4_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_10),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_19),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_21),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);


endmodule