module real_jpeg_18056_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_616;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_1),
.B(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_2),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_2),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_2),
.Y(n_476)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_3),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_3),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_3),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_4),
.A2(n_89),
.B1(n_279),
.B2(n_281),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_4),
.A2(n_281),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_4),
.A2(n_281),
.B1(n_490),
.B2(n_492),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g548 ( 
.A1(n_4),
.A2(n_281),
.B1(n_549),
.B2(n_552),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_5),
.A2(n_376),
.B1(n_378),
.B2(n_379),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_5),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g428 ( 
.A1(n_5),
.A2(n_378),
.B1(n_429),
.B2(n_434),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_5),
.A2(n_378),
.B1(n_541),
.B2(n_544),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_5),
.A2(n_378),
.B1(n_582),
.B2(n_585),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_56),
.B1(n_77),
.B2(n_80),
.Y(n_76)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_6),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_6),
.A2(n_80),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_6),
.A2(n_80),
.B1(n_242),
.B2(n_274),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_6),
.A2(n_80),
.B1(n_361),
.B2(n_364),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_44),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_7),
.A2(n_39),
.B1(n_118),
.B2(n_122),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_7),
.A2(n_39),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_7),
.A2(n_39),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_50),
.B1(n_54),
.B2(n_55),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_54),
.B1(n_130),
.B2(n_133),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_8),
.A2(n_54),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_8),
.A2(n_54),
.B1(n_267),
.B2(n_269),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_9),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_9),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_88),
.B1(n_178),
.B2(n_181),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_9),
.A2(n_88),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_9),
.A2(n_88),
.B1(n_309),
.B2(n_312),
.Y(n_308)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_10),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_10),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_10),
.Y(n_208)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_10),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_10),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_10),
.Y(n_519)
);

BUFx5_ASAP7_75t_L g221 ( 
.A(n_11),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g319 ( 
.A(n_11),
.Y(n_319)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_11),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_12),
.A2(n_325),
.B1(n_326),
.B2(n_328),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_12),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_12),
.A2(n_328),
.B1(n_408),
.B2(n_413),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_12),
.A2(n_328),
.B1(n_482),
.B2(n_488),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_12),
.A2(n_328),
.B1(n_564),
.B2(n_567),
.Y(n_563)
);

OAI32xp33_ASAP7_75t_L g342 ( 
.A1(n_13),
.A2(n_343),
.A3(n_347),
.B1(n_349),
.B2(n_355),
.Y(n_342)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_13),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_13),
.A2(n_40),
.B1(n_354),
.B2(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_13),
.B(n_26),
.Y(n_439)
);

OAI32xp33_ASAP7_75t_L g461 ( 
.A1(n_13),
.A2(n_198),
.A3(n_462),
.B1(n_467),
.B2(n_470),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_13),
.A2(n_354),
.B1(n_497),
.B2(n_499),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_13),
.B(n_140),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_13),
.B(n_318),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_13),
.B(n_93),
.Y(n_597)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_15),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_16),
.Y(n_101)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_16),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_619),
.Y(n_21)
);

OAI221xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_67),
.B1(n_70),
.B2(n_298),
.C(n_613),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_23),
.B(n_67),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_24),
.B(n_291),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_24),
.B(n_291),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_48),
.Y(n_24)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_25),
.A2(n_58),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_38),
.Y(n_25)
);

OR2x6_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_26),
.B(n_49),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_26),
.A2(n_57),
.B1(n_374),
.B2(n_381),
.Y(n_373)
);

AO22x2_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_28),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_32),
.Y(n_180)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_33),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_33),
.Y(n_200)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_35),
.Y(n_163)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_41),
.Y(n_380)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_47),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_48),
.A2(n_68),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_57),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_52),
.Y(n_377)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_68),
.B(n_69),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_68),
.B1(n_76),
.B2(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_58),
.A2(n_69),
.B(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_58),
.A2(n_84),
.B(n_251),
.Y(n_292)
);

OAI22x1_ASAP7_75t_SL g323 ( 
.A1(n_58),
.A2(n_68),
.B1(n_278),
.B2(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_58),
.A2(n_68),
.B1(n_375),
.B2(n_401),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_63),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_63),
.Y(n_405)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_64),
.Y(n_348)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_289),
.C(n_297),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_252),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_72),
.A2(n_615),
.B(n_616),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_188),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_73),
.B(n_188),
.Y(n_616)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_175),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_82),
.B2(n_174),
.Y(n_74)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_75),
.B(n_92),
.C(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_75),
.A2(n_174),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_75),
.B(n_82),
.C(n_175),
.Y(n_290)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2x1_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_91),
.Y(n_82)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_83),
.Y(n_296)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_89),
.B(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_127),
.B1(n_128),
.B2(n_173),
.Y(n_91)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_92),
.B(n_176),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_104),
.B(n_116),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_93),
.B(n_206),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_93),
.B(n_273),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_93),
.A2(n_104),
.B1(n_537),
.B2(n_540),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_93),
.A2(n_104),
.B1(n_481),
.B2(n_540),
.Y(n_557)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_94),
.B(n_117),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_94),
.A2(n_241),
.B1(n_247),
.B2(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_94),
.A2(n_247),
.B1(n_480),
.B2(n_489),
.Y(n_479)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_97),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_97),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_97),
.Y(n_311)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_97),
.Y(n_554)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_101),
.Y(n_234)
);

INVx5_ASAP7_75t_L g314 ( 
.A(n_101),
.Y(n_314)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_101),
.Y(n_523)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_101),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_104),
.B(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_104),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_104),
.A2(n_213),
.B(n_504),
.Y(n_503)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_110),
.B2(n_113),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_106),
.Y(n_531)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_108),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_108),
.Y(n_539)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AO22x2_ASAP7_75t_L g140 ( 
.A1(n_115),
.A2(n_141),
.B1(n_144),
.B2(n_147),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_115),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_115),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_115),
.Y(n_545)
);

INVxp33_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g399 ( 
.A1(n_117),
.A2(n_247),
.B(n_248),
.Y(n_399)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_120),
.Y(n_212)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_127),
.B(n_173),
.C(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

AO21x1_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_138),
.B(n_164),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_129),
.B(n_140),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_129),
.Y(n_284)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_177),
.B(n_186),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_138),
.A2(n_140),
.B1(n_177),
.B2(n_196),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_SL g293 ( 
.A1(n_138),
.A2(n_140),
.B(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_138),
.A2(n_164),
.B(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_139),
.A2(n_165),
.B1(n_197),
.B2(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_139),
.A2(n_166),
.B(n_187),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_139),
.A2(n_165),
.B1(n_335),
.B2(n_407),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_139),
.A2(n_165),
.B1(n_407),
.B2(n_428),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_139),
.A2(n_165),
.B1(n_428),
.B2(n_496),
.Y(n_495)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_152),
.Y(n_139)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_145),
.Y(n_276)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_146),
.Y(n_246)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_156),
.B1(n_160),
.B2(n_162),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_158),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_159),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_159),
.Y(n_353)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_162),
.Y(n_340)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_166),
.Y(n_294)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_170),
.Y(n_412)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_179),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_185),
.Y(n_416)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.C(n_214),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_190),
.Y(n_288)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_203),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_203),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_213),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_205),
.B(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_208),
.Y(n_469)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_214),
.A2(n_215),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_238),
.B(n_249),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_216),
.A2(n_217),
.B1(n_249),
.B2(n_250),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_L g384 ( 
.A1(n_216),
.A2(n_217),
.B1(n_240),
.B2(n_385),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_222),
.B(n_232),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_221),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_222),
.B(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_222),
.A2(n_548),
.B(n_555),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_222),
.A2(n_318),
.B1(n_354),
.B2(n_581),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_222),
.A2(n_563),
.B1(n_581),
.B2(n_595),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_225),
.Y(n_566)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_226),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_227),
.Y(n_571)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_228),
.Y(n_596)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_232),
.Y(n_478)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_237),
.Y(n_367)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_237),
.Y(n_587)
);

INVxp33_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_240),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B(n_248),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_243),
.Y(n_488)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_285),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_253),
.B(n_285),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_255),
.A2(n_257),
.B1(n_258),
.B2(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_255),
.Y(n_448)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_259),
.B(n_447),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_277),
.C(n_282),
.Y(n_259)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_260),
.B(n_387),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_271),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g331 ( 
.A(n_261),
.B(n_271),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_262),
.Y(n_555)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_263),
.Y(n_441)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_265),
.A2(n_360),
.B(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_266),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_270),
.Y(n_534)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_277),
.B(n_283),
.Y(n_387)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g613 ( 
.A1(n_289),
.A2(n_297),
.B(n_614),
.C(n_617),
.D(n_618),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_290),
.B(n_291),
.Y(n_617)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.CI(n_295),
.CON(n_291),
.SN(n_291)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_450),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_391),
.B(n_442),
.C(n_443),
.D(n_449),
.Y(n_300)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_301),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_382),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_302),
.B(n_382),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_330),
.C(n_332),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_304),
.A2(n_330),
.B1(n_331),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_322),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_305),
.B(n_323),
.C(n_329),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_320),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_306),
.B(n_320),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B(n_315),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_307),
.A2(n_308),
.B1(n_360),
.B2(n_368),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_307),
.A2(n_315),
.B(n_478),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_307),
.A2(n_562),
.B1(n_572),
.B2(n_573),
.Y(n_561)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_314),
.Y(n_592)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx6_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_329),
.Y(n_322)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_324),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_341),
.C(n_373),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_333),
.B(n_373),
.Y(n_397)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_359),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_342),
.B(n_359),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_346),
.Y(n_433)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_354),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_354),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_354),
.B(n_530),
.Y(n_529)
);

OAI21xp33_ASAP7_75t_SL g537 ( 
.A1(n_354),
.A2(n_529),
.B(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_367),
.Y(n_551)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_372),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_383),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g390 ( 
.A(n_383),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_386),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_386),
.C(n_388),
.Y(n_445)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.C(n_418),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_392),
.B(n_395),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.C(n_417),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_396),
.B(n_420),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_398),
.B(n_417),
.Y(n_420)
);

MAJx2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.C(n_406),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_399),
.B(n_406),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_400),
.B(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_421),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_419),
.B(n_421),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_424),
.C(n_426),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g609 ( 
.A(n_422),
.B(n_610),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_424),
.A2(n_425),
.B1(n_426),
.B2(n_611),
.Y(n_610)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_426),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_438),
.C(n_440),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_429),
.Y(n_499)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_438),
.A2(n_439),
.B1(n_440),
.B2(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_440),
.Y(n_508)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

NOR3xp33_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_452),
.C(n_455),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_445),
.B(n_446),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_456),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_607),
.B(n_612),
.Y(n_456)
);

AOI21x1_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_510),
.B(n_606),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_500),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_459),
.B(n_500),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_479),
.C(n_495),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_460),
.B(n_603),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_477),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_461),
.B(n_477),
.Y(n_502)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_466),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_479),
.B(n_495),
.Y(n_603)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_489),
.Y(n_504)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_505),
.B1(n_506),
.B2(n_509),
.Y(n_500)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_501),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_502),
.B(n_503),
.C(n_505),
.Y(n_608)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_511),
.A2(n_601),
.B(n_605),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_512),
.A2(n_559),
.B(n_600),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_546),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_513),
.B(n_546),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_535),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_514),
.A2(n_535),
.B1(n_536),
.B2(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_514),
.Y(n_577)
);

OAI32xp33_ASAP7_75t_L g514 ( 
.A1(n_515),
.A2(n_520),
.A3(n_524),
.B1(n_529),
.B2(n_532),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx8_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_547),
.B(n_556),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_547),
.B(n_557),
.C(n_558),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_548),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_558),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_560),
.A2(n_578),
.B(n_599),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_576),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_561),
.B(n_576),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_579),
.A2(n_593),
.B(n_598),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_580),
.B(n_588),
.Y(n_579)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_589),
.B(n_590),
.Y(n_588)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_594),
.B(n_597),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_594),
.B(n_597),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_SL g601 ( 
.A(n_602),
.B(n_604),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_602),
.B(n_604),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_608),
.B(n_609),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_609),
.Y(n_612)
);


endmodule