module fake_jpeg_17889_n_20 (n_3, n_2, n_1, n_0, n_4, n_5, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_20;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_9;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx16f_ASAP7_75t_L g6 ( 
.A(n_2),
.Y(n_6)
);

AOI22xp33_ASAP7_75t_SL g7 ( 
.A1(n_1),
.A2(n_2),
.B1(n_0),
.B2(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_0),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_SL g10 ( 
.A1(n_4),
.A2(n_0),
.B1(n_2),
.B2(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_6),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_13),
.B1(n_14),
.B2(n_3),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_4),
.Y(n_13)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_3),
.C(n_8),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_7),
.B(n_10),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_16),
.B(n_12),
.C(n_6),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_18),
.B(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_19),
.B(n_3),
.Y(n_20)
);


endmodule