module fake_jpeg_29412_n_536 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_536);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_536;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_331;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_15),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_81),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_55),
.Y(n_164)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_62),
.Y(n_108)
);

INVx11_ASAP7_75t_SL g61 ( 
.A(n_28),
.Y(n_61)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_18),
.B(n_14),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_63),
.B(n_26),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_67),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_66),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_18),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_77),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_75),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_79),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_85),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_14),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_82),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_21),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_13),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_101),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_30),
.B(n_13),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_29),
.Y(n_107)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_30),
.B1(n_43),
.B2(n_26),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_117),
.A2(n_143),
.B1(n_69),
.B2(n_83),
.Y(n_208)
);

INVx6_ASAP7_75t_SL g118 ( 
.A(n_61),
.Y(n_118)
);

INVx6_ASAP7_75t_SL g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_55),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_119),
.B(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_56),
.B(n_35),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_130),
.B(n_140),
.Y(n_218)
);

AO22x2_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_50),
.B1(n_43),
.B2(n_53),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_137),
.A2(n_148),
.B1(n_90),
.B2(n_92),
.Y(n_191)
);

CKINVDCx12_ASAP7_75t_R g142 ( 
.A(n_78),
.Y(n_142)
);

CKINVDCx12_ASAP7_75t_R g195 ( 
.A(n_142),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_68),
.A2(n_26),
.B1(n_43),
.B2(n_53),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_71),
.A2(n_52),
.B1(n_49),
.B2(n_19),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_55),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_98),
.B(n_36),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_154),
.B(n_166),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_78),
.Y(n_156)
);

CKINVDCx9p33_ASAP7_75t_R g223 ( 
.A(n_156),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_57),
.B(n_46),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_162),
.B(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_65),
.B(n_46),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_74),
.B(n_36),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_112),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_183),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_108),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_172),
.B(n_187),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_137),
.A2(n_99),
.B1(n_94),
.B2(n_102),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_173),
.A2(n_198),
.B1(n_207),
.B2(n_210),
.Y(n_257)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_175),
.Y(n_253)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

INVx4_ASAP7_75t_SL g233 ( 
.A(n_176),
.Y(n_233)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_126),
.Y(n_177)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

CKINVDCx6p67_ASAP7_75t_R g178 ( 
.A(n_159),
.Y(n_178)
);

INVx4_ASAP7_75t_SL g246 ( 
.A(n_178),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_113),
.B(n_107),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_182),
.B(n_186),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_114),
.A2(n_19),
.B1(n_42),
.B2(n_104),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_122),
.B(n_37),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_37),
.Y(n_187)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_188),
.Y(n_260)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_42),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_193),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_191),
.A2(n_208),
.B1(n_222),
.B2(n_82),
.Y(n_239)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_137),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

CKINVDCx12_ASAP7_75t_R g197 ( 
.A(n_115),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_197),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_79),
.B1(n_76),
.B2(n_88),
.Y(n_198)
);

AND2x2_ASAP7_75t_SL g200 ( 
.A(n_158),
.B(n_75),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_200),
.B(n_210),
.C(n_181),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_114),
.A2(n_136),
.B(n_143),
.C(n_123),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_211),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_116),
.B(n_27),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_216),
.Y(n_245)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

BUFx16f_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_133),
.Y(n_206)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_97),
.B1(n_91),
.B2(n_103),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_139),
.A2(n_100),
.B1(n_93),
.B2(n_73),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_209),
.A2(n_213),
.B1(n_144),
.B2(n_127),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_145),
.A2(n_89),
.B1(n_105),
.B2(n_106),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_146),
.A2(n_48),
.B1(n_41),
.B2(n_27),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_212),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_160),
.A2(n_93),
.B1(n_59),
.B2(n_73),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_214),
.Y(n_252)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_155),
.B(n_41),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_169),
.Y(n_221)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_221),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_145),
.A2(n_52),
.B1(n_66),
.B2(n_59),
.Y(n_222)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_156),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_225),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_164),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_147),
.B1(n_168),
.B2(n_151),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_229),
.A2(n_168),
.B1(n_153),
.B2(n_192),
.Y(n_282)
);

A2O1A1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_201),
.A2(n_223),
.B(n_173),
.C(n_191),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_230),
.A2(n_254),
.B(n_178),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_239),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_148),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_235),
.B(n_183),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_147),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_190),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_223),
.A2(n_161),
.B1(n_146),
.B2(n_164),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g256 ( 
.A1(n_202),
.A2(n_151),
.B1(n_109),
.B2(n_170),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_215),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_200),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_184),
.B(n_22),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_265),
.B(n_268),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_171),
.B(n_22),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_270),
.A2(n_289),
.B(n_262),
.Y(n_319)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_271),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_272),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_273),
.A2(n_256),
.B1(n_240),
.B2(n_230),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_226),
.B(n_171),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_274),
.B(n_276),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_178),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_275),
.B(n_284),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_217),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_277),
.Y(n_323)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx11_ASAP7_75t_SL g279 ( 
.A(n_246),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_279),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_241),
.B(n_200),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_287),
.Y(n_311)
);

INVx11_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_282),
.A2(n_266),
.B1(n_240),
.B2(n_257),
.Y(n_322)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_245),
.B(n_206),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_241),
.A2(n_211),
.B1(n_157),
.B2(n_163),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_285),
.A2(n_292),
.B1(n_257),
.B2(n_266),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_288),
.C(n_302),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_242),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_195),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_247),
.A2(n_220),
.B(n_178),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_204),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_291),
.Y(n_329)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_239),
.A2(n_157),
.B1(n_163),
.B2(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_234),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_293),
.B(n_300),
.Y(n_318)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_294),
.B(n_295),
.Y(n_321)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_248),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_250),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_296),
.Y(n_306)
);

BUFx12f_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_298),
.Y(n_337)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_267),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_299),
.B(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_264),
.B(n_219),
.Y(n_300)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_233),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_301),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_247),
.B(n_174),
.C(n_189),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_247),
.B(n_219),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_305),
.A2(n_331),
.B1(n_333),
.B2(n_334),
.Y(n_345)
);

MAJx2_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_230),
.C(n_252),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_299),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_272),
.A2(n_235),
.B(n_230),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_315),
.A2(n_327),
.B(n_297),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_335),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_319),
.A2(n_293),
.B(n_291),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_286),
.B(n_234),
.C(n_259),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_328),
.C(n_336),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g360 ( 
.A(n_322),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_275),
.A2(n_259),
.B(n_249),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_324),
.A2(n_270),
.B(n_289),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_304),
.A2(n_236),
.B(n_262),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_237),
.C(n_228),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_297),
.A2(n_256),
.B1(n_180),
.B2(n_175),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_297),
.A2(n_273),
.B1(n_280),
.B2(n_269),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_269),
.A2(n_188),
.B1(n_185),
.B2(n_194),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_287),
.B(n_48),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_302),
.B(n_260),
.C(n_232),
.Y(n_336)
);

AOI21xp33_ASAP7_75t_L g338 ( 
.A1(n_309),
.A2(n_303),
.B(n_296),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_330),
.B(n_325),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_321),
.Y(n_341)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_341),
.Y(n_372)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_323),
.Y(n_342)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_301),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_343),
.B(n_349),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_355),
.Y(n_394)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_321),
.Y(n_347)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_347),
.Y(n_379)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_307),
.Y(n_348)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_348),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_319),
.A2(n_285),
.B(n_292),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_323),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_350),
.Y(n_371)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_351),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_352),
.B(n_356),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_353),
.Y(n_377)
);

AND2x6_ASAP7_75t_L g354 ( 
.A(n_306),
.B(n_205),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_362),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_271),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_310),
.B(n_295),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_306),
.Y(n_357)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_369),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_283),
.B1(n_281),
.B2(n_294),
.Y(n_359)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_359),
.Y(n_393)
);

OAI32xp33_ASAP7_75t_L g361 ( 
.A1(n_333),
.A2(n_298),
.A3(n_66),
.B1(n_277),
.B2(n_278),
.Y(n_361)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_310),
.B(n_260),
.C(n_232),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_336),
.C(n_320),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_308),
.B(n_298),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_366),
.Y(n_391)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_365),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_233),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_325),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_368),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_311),
.B(n_298),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_316),
.B(n_141),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g416 ( 
.A(n_370),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_312),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_385),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_388),
.C(n_392),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_339),
.B(n_312),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_339),
.B(n_318),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_386),
.B(n_387),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_352),
.B(n_318),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_363),
.B(n_311),
.C(n_328),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_345),
.A2(n_322),
.B1(n_334),
.B2(n_315),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_389),
.A2(n_348),
.B1(n_258),
.B2(n_238),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_340),
.B(n_317),
.C(n_332),
.Y(n_392)
);

NAND2x1p5_ASAP7_75t_L g395 ( 
.A(n_346),
.B(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_314),
.Y(n_396)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_396),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_344),
.B(n_337),
.Y(n_400)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_355),
.B(n_307),
.Y(n_401)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_399),
.A2(n_369),
.B1(n_349),
.B2(n_355),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_402),
.A2(n_407),
.B1(n_410),
.B2(n_414),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_396),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_403),
.B(n_408),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_326),
.Y(n_405)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_406),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_376),
.A2(n_369),
.B1(n_361),
.B2(n_360),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g408 ( 
.A(n_394),
.B(n_343),
.CI(n_331),
.CON(n_408),
.SN(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_377),
.A2(n_360),
.B1(n_353),
.B2(n_354),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_381),
.B(n_307),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_420),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_375),
.A2(n_365),
.B(n_332),
.Y(n_413)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_413),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_342),
.B1(n_350),
.B2(n_317),
.Y(n_414)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_205),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_426),
.Y(n_448)
);

FAx1_ASAP7_75t_SL g417 ( 
.A(n_394),
.B(n_348),
.CI(n_110),
.CON(n_417),
.SN(n_417)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_417),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_372),
.B1(n_379),
.B2(n_371),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_253),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_419),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_375),
.A2(n_176),
.B(n_12),
.Y(n_420)
);

A2O1A1O1Ixp25_ASAP7_75t_L g422 ( 
.A1(n_395),
.A2(n_179),
.B(n_177),
.C(n_12),
.D(n_13),
.Y(n_422)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_422),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_11),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_428),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_212),
.Y(n_425)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_425),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g426 ( 
.A(n_385),
.B(n_110),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_401),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_429),
.Y(n_440)
);

INVx3_ASAP7_75t_SL g433 ( 
.A(n_425),
.Y(n_433)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_433),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_416),
.B(n_383),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_446),
.Y(n_462)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_442),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_384),
.C(n_386),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_447),
.C(n_451),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_445),
.A2(n_402),
.B1(n_389),
.B2(n_407),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_409),
.B(n_387),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_388),
.C(n_421),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_392),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_424),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_398),
.C(n_394),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_410),
.B(n_382),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_453),
.B(n_418),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_458),
.Y(n_478)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_450),
.B(n_415),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_461),
.Y(n_485)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_439),
.Y(n_460)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_426),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_408),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_466),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_437),
.A2(n_414),
.B1(n_411),
.B2(n_430),
.Y(n_464)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_464),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_408),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_468),
.Y(n_479)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_398),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_438),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_469),
.B(n_470),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_436),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_471),
.B(n_472),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_432),
.B(n_417),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_474),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_467),
.B(n_435),
.C(n_434),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_454),
.A2(n_438),
.B(n_469),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_456),
.A2(n_437),
.B1(n_452),
.B2(n_445),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_480),
.A2(n_429),
.B1(n_440),
.B2(n_461),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_435),
.C(n_434),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_489),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_455),
.A2(n_442),
.B(n_395),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_484),
.A2(n_440),
.B(n_422),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_448),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_486),
.B(n_458),
.C(n_462),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_468),
.B(n_417),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_493),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_485),
.Y(n_510)
);

BUFx24_ASAP7_75t_SL g493 ( 
.A(n_481),
.Y(n_493)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_494),
.Y(n_512)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_496),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_449),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_478),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_499),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_373),
.C(n_378),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_378),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_500),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_167),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_501),
.B(n_0),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_487),
.A2(n_153),
.B1(n_1),
.B2(n_5),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_503),
.A2(n_504),
.B1(n_52),
.B2(n_1),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_475),
.A2(n_484),
.B1(n_488),
.B2(n_478),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_494),
.A2(n_479),
.B(n_486),
.Y(n_507)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_507),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_510),
.B(n_511),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_490),
.A2(n_485),
.B(n_110),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_513),
.B(n_515),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g514 ( 
.A1(n_504),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_514)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_6),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_497),
.A2(n_0),
.B(n_6),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_512),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_519),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_502),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_501),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_523),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_521),
.B(n_509),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_522),
.C(n_523),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_518),
.A2(n_509),
.B(n_505),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_526),
.A2(n_514),
.B(n_8),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_528),
.B(n_530),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_529),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_7),
.C(n_8),
.Y(n_530)
);

NOR3xp33_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_527),
.C(n_8),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_533),
.A2(n_531),
.B(n_9),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g535 ( 
.A(n_534),
.B(n_7),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_535),
.A2(n_9),
.B(n_10),
.Y(n_536)
);


endmodule