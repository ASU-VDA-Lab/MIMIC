module fake_jpeg_30627_n_143 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx24_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_38),
.Y(n_50)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_12),
.B(n_5),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_40),
.Y(n_45)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_20),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_14),
.B1(n_23),
.B2(n_19),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_48),
.A2(n_49),
.B1(n_37),
.B2(n_39),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_14),
.B1(n_23),
.B2(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_28),
.B(n_13),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_26),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_25),
.B(n_33),
.C(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_56),
.B(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_25),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_60),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_5),
.Y(n_58)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_19),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_36),
.C(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_63),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_48),
.B(n_36),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_67),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_32),
.C(n_31),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_24),
.B(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_72),
.Y(n_87)
);

XNOR2x1_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_22),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_78),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_42),
.B1(n_24),
.B2(n_53),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_34),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_42),
.B1(n_29),
.B2(n_30),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_56),
.B1(n_59),
.B2(n_73),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_104),
.B1(n_106),
.B2(n_107),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.C(n_87),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_100),
.C(n_105),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_67),
.C(n_72),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_102),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_65),
.B1(n_69),
.B2(n_68),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_85),
.B(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_82),
.A2(n_78),
.B(n_70),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_105),
.A2(n_81),
.B(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_84),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_116),
.C(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_81),
.B1(n_95),
.B2(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_96),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_102),
.B(n_100),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_124),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_120),
.B(n_122),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_123),
.C(n_108),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g122 ( 
.A1(n_109),
.A2(n_80),
.B(n_92),
.C(n_79),
.D(n_9),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_113),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_129),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_123),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_112),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_128),
.B(n_117),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_128),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_111),
.B1(n_110),
.B2(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_126),
.Y(n_135)
);

OAI221xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_114),
.C(n_92),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_137),
.A2(n_133),
.B(n_131),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_139),
.B(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_11),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_74),
.Y(n_142)
);

BUFx24_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);


endmodule