module fake_netlist_1_1029_n_32 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_4), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_9), .B(n_3), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_9), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_10), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
INVx5_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
CKINVDCx8_ASAP7_75t_R g17 ( .A(n_14), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_13), .B(n_0), .Y(n_18) );
AND2x2_ASAP7_75t_L g19 ( .A(n_15), .B(n_1), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_15), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_11), .B1(n_12), .B2(n_5), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_16), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_23), .Y(n_25) );
XNOR2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_21), .Y(n_26) );
NOR2x1p5_ASAP7_75t_L g27 ( .A(n_26), .B(n_24), .Y(n_27) );
OAI322xp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_18), .A3(n_20), .B1(n_19), .B2(n_24), .C1(n_8), .C2(n_1), .Y(n_28) );
NAND3xp33_ASAP7_75t_SL g29 ( .A(n_28), .B(n_20), .C(n_6), .Y(n_29) );
OAI221xp5_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_2), .B1(n_6), .B2(n_7), .C(n_8), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_29), .Y(n_31) );
AOI22xp5_ASAP7_75t_SL g32 ( .A1(n_31), .A2(n_30), .B1(n_2), .B2(n_10), .Y(n_32) );
endmodule