module fake_jpeg_3119_n_101 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_32),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_30),
.B1(n_35),
.B2(n_38),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_44),
.B1(n_37),
.B2(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_29),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_31),
.B1(n_35),
.B2(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_52),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_40),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_42),
.B(n_45),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_1),
.B(n_2),
.Y(n_66)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_53),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_48),
.B1(n_45),
.B2(n_37),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_4),
.Y(n_74)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_40),
.C(n_11),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_52),
.B(n_5),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_70),
.B1(n_71),
.B2(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_4),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_5),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_6),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

OAI32xp33_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_84),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_20),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_91),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_21),
.B(n_25),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_86),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_92),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_89),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_93),
.C(n_84),
.Y(n_99)
);

O2A1O1Ixp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_88),
.B(n_83),
.C(n_79),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_87),
.Y(n_101)
);


endmodule