module real_jpeg_25592_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_1),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_137),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_51),
.B1(n_52),
.B2(n_137),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_137),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_2),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_2),
.A2(n_28),
.B1(n_57),
.B2(n_58),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_2),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_43),
.B(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_3),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_3),
.B(n_31),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_134),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_3),
.B(n_53),
.C(n_58),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_3),
.B(n_66),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_108),
.B1(n_227),
.B2(n_234),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_6),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_127),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_127),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_127),
.Y(n_271)
);

INVx8_ASAP7_75t_SL g37 ( 
.A(n_7),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_8),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_26),
.B1(n_125),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_8),
.A2(n_51),
.B1(n_52),
.B2(n_125),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g224 ( 
.A1(n_8),
.A2(n_57),
.B1(n_58),
.B2(n_125),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_9),
.A2(n_41),
.B1(n_57),
.B2(n_58),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_9),
.A2(n_41),
.B1(n_51),
.B2(n_52),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_73),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_10),
.A2(n_51),
.B1(n_52),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_73),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_12),
.A2(n_51),
.B1(n_52),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_12),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_61),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_294)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_15),
.Y(n_117)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_15),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_84),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_78),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_20),
.A2(n_21),
.B1(n_74),
.B2(n_326),
.Y(n_332)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_45),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_47),
.C(n_62),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_31),
.B2(n_40),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_24),
.A2(n_30),
.B(n_75),
.Y(n_74)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_27),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_29),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_29),
.A2(n_40),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_29),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_29),
.A2(n_31),
.B1(n_136),
.B2(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_29),
.A2(n_31),
.B1(n_144),
.B2(n_271),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_29),
.A2(n_271),
.B(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_29),
.A2(n_88),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_38),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_30),
.A2(n_130),
.B1(n_131),
.B2(n_135),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_30),
.B(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_32),
.A2(n_33),
.B1(n_67),
.B2(n_68),
.Y(n_71)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_32),
.A2(n_36),
.B(n_133),
.C(n_151),
.Y(n_150)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_32),
.B(n_134),
.CON(n_179),
.SN(n_179)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_33),
.B(n_35),
.C(n_146),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g178 ( 
.A1(n_33),
.A2(n_52),
.A3(n_67),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_44),
.B(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_62),
.B2(n_63),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_74),
.C(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_46),
.A2(n_47),
.B1(n_79),
.B2(n_329),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_56),
.B(n_59),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_49),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_49),
.A2(n_60),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_49),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_49),
.A2(n_188),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_49),
.A2(n_187),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_49),
.A2(n_186),
.B1(n_187),
.B2(n_207),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_49),
.A2(n_187),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_49),
.A2(n_121),
.B(n_265),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_52),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_51),
.B(n_68),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_52),
.B(n_209),
.Y(n_208)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_56)
);

BUFx24_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_56),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_56),
.B(n_59),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_56),
.B(n_134),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_57),
.B(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_64),
.A2(n_123),
.B(n_126),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_66),
.B(n_70),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_65),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_66),
.B(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_66),
.A2(n_70),
.B1(n_170),
.B2(n_179),
.Y(n_184)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_69),
.A2(n_128),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_72),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_74),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_74),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_78),
.B(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_79),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_81),
.A2(n_123),
.B1(n_128),
.B2(n_297),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_83),
.A2(n_123),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI321xp33_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_323),
.A3(n_333),
.B1(n_336),
.B2(n_337),
.C(n_340),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_302),
.B(n_322),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_279),
.B(n_301),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_171),
.B(n_255),
.C(n_278),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_156),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_156),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_140),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_118),
.B1(n_138),
.B2(n_139),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_101),
.B(n_139),
.C(n_140),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_102),
.B(n_107),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_103),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_104),
.B(n_309),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_112),
.B(n_114),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_108),
.A2(n_114),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_108),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_108),
.A2(n_224),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_108),
.A2(n_182),
.B(n_235),
.Y(n_287)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_109),
.B(n_115),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_109),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_111),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_117),
.Y(n_219)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.C(n_129),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_119),
.A2(n_120),
.B1(n_122),
.B2(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_128),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_134),
.B(n_235),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_149),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_147),
.B2(n_148),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_143),
.B(n_147),
.C(n_149),
.Y(n_276)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_152),
.B1(n_153),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_155),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_162),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_157),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_162),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_166),
.B1(n_167),
.B2(n_193),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_165),
.B(n_218),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_250),
.B(n_254),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_201),
.B(n_249),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_189),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_176),
.B(n_189),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_184),
.C(n_185),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_177),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_184),
.B(n_185),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_190),
.B(n_197),
.C(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_196),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_199),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_244),
.B(n_248),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_220),
.B(n_243),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_204),
.B(n_210),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_208),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_230),
.B(n_242),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_229),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_237),
.B(n_241),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_252),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_257),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_276),
.B2(n_277),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_267),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_267),
.C(n_277),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_266),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_261),
.B(n_266),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_263),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_275),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_280),
.B(n_281),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_300),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_288),
.B1(n_298),
.B2(n_299),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_299),
.C(n_300),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_286),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_287),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_286),
.A2(n_316),
.B(n_317),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_292),
.C(n_295),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_294),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_303),
.B(n_304),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_320),
.B2(n_321),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_312),
.B1(n_318),
.B2(n_319),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_307),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_319),
.C(n_321),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_310),
.B(n_311),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_325),
.C(n_330),
.Y(n_324)
);

FAx1_ASAP7_75t_L g335 ( 
.A(n_311),
.B(n_325),
.CI(n_330),
.CON(n_335),
.SN(n_335)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_331),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_324),
.B(n_331),
.Y(n_337)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_335),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_335),
.Y(n_338)
);


endmodule