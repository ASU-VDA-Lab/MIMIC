module fake_jpeg_19703_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_288;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_303;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_18),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_22),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_69),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_53),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_48),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_33),
.B1(n_19),
.B2(n_23),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_49),
.A2(n_67),
.B1(n_18),
.B2(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_19),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_60),
.B1(n_65),
.B2(n_31),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_61),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_56),
.Y(n_76)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_33),
.B1(n_23),
.B2(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_34),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_37),
.A2(n_26),
.B1(n_34),
.B2(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_28),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_20),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_81),
.B1(n_88),
.B2(n_77),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_80),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_53),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_45),
.C(n_71),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_29),
.B1(n_20),
.B2(n_18),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_41),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_119),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_98),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_102),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_62),
.C(n_43),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_62),
.C(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_101),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_47),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_21),
.B(n_50),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_72),
.A2(n_61),
.B(n_31),
.C(n_68),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_80),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_105),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_43),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_111),
.B1(n_86),
.B2(n_70),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_41),
.C(n_43),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_52),
.B1(n_64),
.B2(n_58),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_114),
.B1(n_94),
.B2(n_75),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_82),
.A2(n_52),
.B1(n_58),
.B2(n_66),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_31),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_41),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_90),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_140),
.Y(n_146)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_129),
.Y(n_162)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_96),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_132),
.A2(n_137),
.B1(n_111),
.B2(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_136),
.A2(n_138),
.B1(n_113),
.B2(n_114),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_85),
.B1(n_86),
.B2(n_93),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_107),
.A2(n_86),
.B1(n_85),
.B2(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_97),
.B(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_31),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_142),
.B(n_144),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_50),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_30),
.Y(n_144)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_105),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_106),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_137),
.B1(n_126),
.B2(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_120),
.B(n_100),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_164),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_151),
.A2(n_165),
.B1(n_138),
.B2(n_140),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_115),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_156),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_101),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_131),
.B(n_102),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_159),
.A2(n_167),
.B(n_127),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_124),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_170),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_118),
.B1(n_103),
.B2(n_91),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_166),
.Y(n_195)
);

AOI31xp33_ASAP7_75t_SL g167 ( 
.A1(n_126),
.A2(n_83),
.A3(n_93),
.B(n_21),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

NOR2x1_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_83),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_21),
.B(n_30),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_169),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_21),
.C(n_83),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_123),
.C(n_21),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g172 ( 
.A1(n_130),
.A2(n_30),
.A3(n_27),
.B1(n_93),
.B2(n_21),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_91),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_139),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_177),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_139),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_159),
.A2(n_127),
.B1(n_143),
.B2(n_136),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_179),
.A2(n_180),
.B(n_188),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_133),
.B1(n_132),
.B2(n_144),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_197),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_151),
.B1(n_160),
.B2(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_171),
.C(n_159),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_27),
.C(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_165),
.Y(n_194)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_129),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_156),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_174),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_208),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_158),
.Y(n_200)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_200),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_10),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_202),
.A2(n_211),
.B1(n_185),
.B2(n_179),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_178),
.B(n_168),
.C(n_154),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_160),
.Y(n_209)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_154),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_166),
.B1(n_147),
.B2(n_155),
.Y(n_211)
);

AOI322xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_166),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_7),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_128),
.C(n_30),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_213),
.B(n_218),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_180),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_219),
.A2(n_191),
.B(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_223),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_203),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_216),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_227),
.B(n_236),
.Y(n_249)
);

AND2x2_ASAP7_75t_SL g228 ( 
.A(n_209),
.B(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_229),
.A2(n_235),
.B1(n_207),
.B2(n_205),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_199),
.A2(n_196),
.B1(n_177),
.B2(n_197),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_211),
.B1(n_217),
.B2(n_4),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_232),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_202),
.A2(n_187),
.B1(n_27),
.B2(n_0),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_27),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_220),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_215),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_213),
.C(n_201),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_241),
.A2(n_230),
.B1(n_232),
.B2(n_238),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_243),
.B(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_216),
.C(n_206),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_248),
.C(n_252),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_206),
.Y(n_245)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_229),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_10),
.C(n_3),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_10),
.C(n_4),
.Y(n_252)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_223),
.B(n_11),
.Y(n_254)
);

XOR2x1_ASAP7_75t_SL g265 ( 
.A(n_254),
.B(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_11),
.C(n_7),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_256),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_261),
.B1(n_268),
.B2(n_249),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_238),
.B1(n_231),
.B2(n_222),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_255),
.A2(n_228),
.B(n_221),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_235),
.B(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_242),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_0),
.B1(n_9),
.B2(n_12),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_265),
.A2(n_252),
.B1(n_248),
.B2(n_256),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_249),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_253),
.A2(n_231),
.B1(n_228),
.B2(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_15),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_267),
.A2(n_245),
.B1(n_257),
.B2(n_262),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_280),
.B1(n_268),
.B2(n_261),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_234),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_273),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_279),
.C(n_12),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_278),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_276),
.A2(n_266),
.B1(n_265),
.B2(n_260),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_266),
.C(n_244),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_13),
.C(n_14),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_8),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_273),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_283),
.B(n_286),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_SL g285 ( 
.A(n_270),
.B(n_269),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_12),
.C(n_13),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_288),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_291),
.B(n_294),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_272),
.B(n_275),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_295),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_13),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_15),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_299),
.C(n_289),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_294),
.A2(n_14),
.B(n_15),
.Y(n_299)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_298),
.B(n_14),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_303),
.A2(n_0),
.B(n_301),
.Y(n_304)
);


endmodule