module fake_jpeg_7920_n_140 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_140);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_140;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx10_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx4f_ASAP7_75t_SL g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_32),
.Y(n_51)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_36),
.B(n_21),
.Y(n_39)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_3),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_50),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_16),
.B1(n_21),
.B2(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_16),
.B1(n_37),
.B2(n_31),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_2),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_18),
.B(n_26),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_32),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_27),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_66),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_55),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_3),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_33),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_44),
.B(n_14),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_69),
.B1(n_42),
.B2(n_40),
.Y(n_85)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_51),
.A2(n_30),
.B1(n_37),
.B2(n_32),
.Y(n_59)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_68),
.A3(n_41),
.B1(n_32),
.B2(n_35),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_5),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_6),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_52),
.A2(n_19),
.B1(n_25),
.B2(n_13),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_25),
.B1(n_13),
.B2(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_74),
.B1(n_83),
.B2(n_43),
.Y(n_96)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

OAI32xp33_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_13),
.A3(n_15),
.B1(n_28),
.B2(n_29),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_57),
.B(n_61),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_86),
.A2(n_88),
.B(n_90),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_55),
.C(n_67),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_91),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_92),
.B(n_96),
.Y(n_99)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_59),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_43),
.Y(n_104)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_91),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_103),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_108),
.B1(n_88),
.B2(n_96),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_106),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_79),
.C(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_78),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_97),
.A2(n_89),
.B1(n_93),
.B2(n_98),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_70),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_105),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_107),
.C(n_108),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_112),
.B(n_113),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_75),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.C(n_54),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_99),
.A2(n_86),
.B1(n_81),
.B2(n_90),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_64),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_120),
.C(n_122),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_62),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_19),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_56),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_123),
.A2(n_13),
.B(n_59),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_126),
.B1(n_121),
.B2(n_8),
.Y(n_129)
);

AOI21x1_ASAP7_75t_SL g126 ( 
.A1(n_119),
.A2(n_111),
.B(n_115),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_128),
.C(n_28),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_130),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_48),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_7),
.B(n_9),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_10),
.B(n_32),
.C(n_38),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_127),
.B1(n_12),
.B2(n_10),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_134),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_129),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_136),
.B(n_29),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_38),
.Y(n_140)
);


endmodule