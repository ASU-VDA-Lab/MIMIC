module fake_jpeg_3626_n_104 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_38),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_29),
.Y(n_48)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_31),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_33),
.B1(n_31),
.B2(n_35),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_55),
.B1(n_46),
.B2(n_36),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_40),
.B1(n_32),
.B2(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

NOR3xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_6),
.C(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_60),
.B(n_14),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_64),
.Y(n_66)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_49),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_75),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_5),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_49),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_59),
.B(n_66),
.Y(n_79)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_82),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_79),
.A2(n_86),
.B(n_12),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_63),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_20),
.C(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_76),
.B(n_8),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_8),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

AOI322xp5_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_13),
.A3(n_21),
.B1(n_22),
.B2(n_24),
.C1(n_26),
.C2(n_28),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_94),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_96),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_83),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_86),
.B1(n_92),
.B2(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_91),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g104 ( 
.A(n_103),
.Y(n_104)
);


endmodule