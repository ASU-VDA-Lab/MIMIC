module fake_jpeg_25768_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

AND2x4_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_1),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_43),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_47)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_20),
.B(n_1),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_46),
.A2(n_55),
.B1(n_63),
.B2(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.C(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_19),
.B1(n_18),
.B2(n_30),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_40),
.B1(n_21),
.B2(n_22),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_55)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_20),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_60),
.B(n_15),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_27),
.B1(n_24),
.B2(n_6),
.Y(n_89)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_41),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_31),
.B1(n_21),
.B2(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_80),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_59),
.B(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_82),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_49),
.A2(n_45),
.B1(n_17),
.B2(n_23),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_23),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_84),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_17),
.B1(n_26),
.B2(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_85),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_88),
.B(n_55),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_62),
.B1(n_57),
.B2(n_58),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_54),
.A3(n_63),
.B1(n_47),
.B2(n_67),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_54),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_97),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_76),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_99),
.B(n_104),
.Y(n_133)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_107),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_59),
.B(n_63),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_109),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_78),
.B(n_47),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_42),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_71),
.B(n_47),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_126),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_87),
.B1(n_73),
.B2(n_82),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_87),
.C(n_73),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_99),
.C(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_102),
.A2(n_57),
.B1(n_85),
.B2(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_79),
.B1(n_46),
.B2(n_83),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_83),
.B1(n_79),
.B2(n_56),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_127),
.B(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_15),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_92),
.A2(n_56),
.B1(n_37),
.B2(n_42),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_123),
.B1(n_115),
.B2(n_133),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_132),
.A2(n_96),
.B(n_103),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_137),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_101),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_136),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_110),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_105),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_145),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_131),
.C(n_115),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_141),
.B(n_151),
.C(n_153),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_123),
.B1(n_100),
.B2(n_112),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_94),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_94),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_149),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_41),
.CI(n_42),
.CON(n_149),
.SN(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_37),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_104),
.C(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_113),
.B(n_90),
.C(n_107),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_154),
.A2(n_64),
.B1(n_53),
.B2(n_86),
.Y(n_163)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_165),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_161),
.B(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_93),
.B1(n_90),
.B2(n_56),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_93),
.B(n_5),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_4),
.B(n_5),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_6),
.B(n_7),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_64),
.B1(n_27),
.B2(n_14),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_27),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_151),
.C(n_153),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_139),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_170),
.Y(n_177)
);

A2O1A1O1Ixp25_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_135),
.B(n_138),
.C(n_142),
.D(n_150),
.Y(n_179)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_171),
.C(n_166),
.Y(n_194)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_134),
.B(n_149),
.C(n_148),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_181),
.Y(n_191)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_168),
.B(n_160),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_155),
.B(n_154),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g197 ( 
.A(n_183),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_14),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_149),
.C(n_8),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_6),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_174),
.B(n_167),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_186),
.Y(n_204)
);

NAND4xp25_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_157),
.C(n_169),
.D(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_190),
.B(n_195),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_192),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_185),
.C(n_178),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_181),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_196)
);

AOI31xp67_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_9),
.A3(n_11),
.B(n_12),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_204),
.C(n_194),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_202),
.Y(n_212)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_197),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_11),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_173),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_205),
.B(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_207),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_196),
.B(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_209),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_189),
.C(n_187),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_196),
.B(n_176),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_211),
.A2(n_203),
.B1(n_176),
.B2(n_204),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

AOI21x1_ASAP7_75t_L g216 ( 
.A1(n_212),
.A2(n_12),
.B(n_13),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_12),
.B(n_13),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_220),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_13),
.Y(n_220)
);

BUFx24_ASAP7_75t_SL g222 ( 
.A(n_219),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_214),
.B(n_217),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_221),
.Y(n_225)
);


endmodule