module fake_ariane_577_n_1240 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1240);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1240;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_611;
wire n_365;
wire n_238;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1218;
wire n_221;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_1072;
wire n_695;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_1103;
wire n_825;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_617;
wire n_543;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_73),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_86),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_94),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_40),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_154),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_66),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_28),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_87),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_64),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_111),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_61),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_79),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_55),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_32),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_9),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_28),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_34),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_34),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_103),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_147),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_119),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_40),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_131),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_109),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_142),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_99),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_83),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_181),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_167),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_31),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_56),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_114),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_120),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_157),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_149),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_49),
.Y(n_237)
);

INVxp33_ASAP7_75t_SL g238 ( 
.A(n_122),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_183),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_88),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_13),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_164),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_165),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_160),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_33),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_139),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_161),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_130),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_54),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_16),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_74),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_68),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_43),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_170),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_190),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_110),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_135),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_180),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_129),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_117),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_107),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_32),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_124),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_92),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_116),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_47),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_71),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_50),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_115),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_24),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_145),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_118),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_174),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_58),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_1),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_39),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_80),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_3),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_41),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_72),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_153),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_95),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_9),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_144),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_98),
.Y(n_294)
);

BUFx10_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_52),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_125),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_127),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_159),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_84),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_23),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_162),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_89),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_4),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_59),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_27),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_158),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_188),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_48),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_136),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_219),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_268),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_225),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_228),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_227),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_232),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_240),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_221),
.B(n_0),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_193),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_195),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_256),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_271),
.Y(n_327)
);

NAND2xp33_ASAP7_75t_R g328 ( 
.A(n_191),
.B(n_197),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_198),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_211),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_195),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_213),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_198),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_208),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_253),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_208),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_278),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_235),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_214),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_285),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_285),
.B(n_0),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_246),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_255),
.B(n_1),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_277),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_261),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_215),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_215),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_215),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_235),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_272),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_277),
.B(n_2),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_196),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_295),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_288),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_279),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_L g362 ( 
.A(n_279),
.B(n_2),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_292),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_192),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_194),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_298),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_255),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_305),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_307),
.B(n_3),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_269),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_289),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_199),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_201),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_210),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_205),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_209),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_216),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_217),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_218),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_224),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_206),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_231),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_226),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_191),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_250),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_230),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_242),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_220),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_222),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_243),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_248),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_262),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_282),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_291),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_250),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_197),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_293),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_308),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_309),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_223),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_200),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_396),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_314),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_342),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_SL g408 ( 
.A(n_397),
.B(n_200),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_400),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_377),
.B(n_202),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_342),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_342),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_400),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_310),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_353),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_238),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_312),
.A2(n_238),
.B1(n_203),
.B2(n_204),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_373),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_375),
.B(n_311),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_328),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_347),
.B(n_266),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_266),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_378),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_380),
.A2(n_235),
.B(n_294),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g432 ( 
.A1(n_381),
.A2(n_235),
.B(n_203),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_384),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_331),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_393),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_399),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_401),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_332),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_335),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_338),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_340),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_341),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g453 ( 
.A(n_349),
.B(n_265),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_344),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_317),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_319),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_320),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_322),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_345),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_379),
.B(n_202),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_352),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_354),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_315),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_359),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_330),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_323),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_369),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_329),
.Y(n_471)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_385),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_457),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_425),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_389),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_424),
.A2(n_397),
.B1(n_357),
.B2(n_324),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_424),
.B(n_356),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_457),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_469),
.B(n_390),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_469),
.B(n_402),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_456),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_469),
.A2(n_357),
.B1(n_324),
.B2(n_348),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_316),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_435),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_469),
.B(n_464),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_453),
.B(n_318),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g491 ( 
.A(n_405),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_426),
.B(n_235),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_463),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_458),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_435),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_458),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_415),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_415),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_469),
.B(n_333),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_456),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_425),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_416),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_435),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_460),
.B(n_463),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_404),
.B(n_362),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g510 ( 
.A(n_404),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_422),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_460),
.B(n_343),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_463),
.B(n_346),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_456),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_463),
.B(n_467),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_467),
.B(n_355),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_435),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_467),
.B(n_360),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_469),
.B(n_366),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_406),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_430),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_459),
.B(n_361),
.Y(n_527)
);

AND2x6_ASAP7_75t_L g528 ( 
.A(n_426),
.B(n_300),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_433),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_428),
.Y(n_531)
);

INVx8_ASAP7_75t_L g532 ( 
.A(n_426),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_432),
.B(n_204),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_443),
.Y(n_534)
);

OAI22xp33_ASAP7_75t_L g535 ( 
.A1(n_472),
.A2(n_339),
.B1(n_334),
.B2(n_336),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_443),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_426),
.A2(n_334),
.B1(n_336),
.B2(n_339),
.Y(n_538)
);

AO22x2_ASAP7_75t_L g539 ( 
.A1(n_466),
.A2(n_383),
.B1(n_382),
.B2(n_321),
.Y(n_539)
);

INVx1_ASAP7_75t_SL g540 ( 
.A(n_471),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_443),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_433),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_477),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_497),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_498),
.Y(n_546)
);

AO22x2_ASAP7_75t_L g547 ( 
.A1(n_539),
.A2(n_421),
.B1(n_321),
.B2(n_326),
.Y(n_547)
);

AO22x2_ASAP7_75t_L g548 ( 
.A1(n_539),
.A2(n_421),
.B1(n_326),
.B2(n_327),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_499),
.A2(n_419),
.B1(n_467),
.B2(n_468),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_503),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_504),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_491),
.Y(n_552)
);

NAND2x1p5_ASAP7_75t_L g553 ( 
.A(n_515),
.B(n_459),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_508),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_515),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

OAI221xp5_ASAP7_75t_L g557 ( 
.A1(n_510),
.A2(n_466),
.B1(n_417),
.B2(n_423),
.C(n_465),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_528),
.A2(n_408),
.B1(n_363),
.B2(n_459),
.Y(n_558)
);

NAND2xp33_ASAP7_75t_L g559 ( 
.A(n_478),
.B(n_464),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_514),
.Y(n_560)
);

AO22x2_ASAP7_75t_L g561 ( 
.A1(n_539),
.A2(n_327),
.B1(n_461),
.B2(n_312),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_480),
.A2(n_464),
.B1(n_410),
.B2(n_462),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_486),
.B(n_465),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_518),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_524),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_526),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_510),
.B(n_464),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_531),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_530),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_543),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_480),
.B(n_464),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_480),
.A2(n_464),
.B1(n_403),
.B2(n_445),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_499),
.B(n_370),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_540),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_477),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_527),
.B(n_507),
.Y(n_576)
);

BUFx8_ASAP7_75t_L g577 ( 
.A(n_486),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_525),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_485),
.B(n_368),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_473),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_525),
.Y(n_581)
);

AO22x2_ASAP7_75t_L g582 ( 
.A1(n_539),
.A2(n_461),
.B1(n_470),
.B2(n_383),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_490),
.B(n_409),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_475),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_523),
.A2(n_363),
.B1(n_440),
.B2(n_438),
.Y(n_585)
);

OR2x2_ASAP7_75t_SL g586 ( 
.A(n_490),
.B(n_370),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_479),
.B(n_470),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_481),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_532),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_507),
.B(n_437),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_487),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_507),
.B(n_429),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_523),
.B(n_371),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_409),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_496),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_493),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_512),
.B(n_446),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_482),
.B(n_414),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_506),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_L g601 ( 
.A1(n_513),
.A2(n_438),
.B(n_437),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_519),
.B(n_429),
.Y(n_602)
);

AO22x2_ASAP7_75t_L g603 ( 
.A1(n_538),
.A2(n_382),
.B1(n_371),
.B2(n_429),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_517),
.Y(n_604)
);

AO22x2_ASAP7_75t_L g605 ( 
.A1(n_535),
.A2(n_429),
.B1(n_445),
.B2(n_442),
.Y(n_605)
);

AO22x2_ASAP7_75t_L g606 ( 
.A1(n_528),
.A2(n_442),
.B1(n_444),
.B2(n_441),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_522),
.B(n_439),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_532),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_482),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_474),
.Y(n_610)
);

NAND2x1_ASAP7_75t_L g611 ( 
.A(n_476),
.B(n_446),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_528),
.B(n_439),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_483),
.B(n_528),
.Y(n_614)
);

NAND2x1p5_ASAP7_75t_L g615 ( 
.A(n_483),
.B(n_414),
.Y(n_615)
);

AO22x2_ASAP7_75t_L g616 ( 
.A1(n_528),
.A2(n_444),
.B1(n_441),
.B2(n_440),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_532),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_474),
.Y(n_618)
);

OAI221xp5_ASAP7_75t_L g619 ( 
.A1(n_533),
.A2(n_417),
.B1(n_423),
.B2(n_455),
.C(n_448),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_489),
.B(n_313),
.Y(n_620)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_528),
.A2(n_455),
.B1(n_454),
.B2(n_451),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_474),
.Y(n_622)
);

NAND2x1p5_ASAP7_75t_L g623 ( 
.A(n_488),
.B(n_456),
.Y(n_623)
);

AO22x2_ASAP7_75t_L g624 ( 
.A1(n_489),
.A2(n_454),
.B1(n_451),
.B2(n_450),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_501),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_501),
.B(n_446),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_492),
.B(n_446),
.Y(n_627)
);

AO22x2_ASAP7_75t_L g628 ( 
.A1(n_492),
.A2(n_448),
.B1(n_450),
.B2(n_436),
.Y(n_628)
);

OAI221xp5_ASAP7_75t_L g629 ( 
.A1(n_533),
.A2(n_456),
.B1(n_452),
.B2(n_449),
.C(n_447),
.Y(n_629)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_501),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_492),
.B(n_446),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_488),
.Y(n_632)
);

BUFx6f_ASAP7_75t_SL g633 ( 
.A(n_492),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_502),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_492),
.B(n_446),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_509),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_492),
.B(n_456),
.Y(n_637)
);

OAI221xp5_ASAP7_75t_L g638 ( 
.A1(n_533),
.A2(n_452),
.B1(n_449),
.B2(n_447),
.C(n_436),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_509),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_502),
.Y(n_640)
);

AO22x2_ASAP7_75t_L g641 ( 
.A1(n_509),
.A2(n_452),
.B1(n_449),
.B2(n_447),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_SL g642 ( 
.A(n_589),
.B(n_520),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_576),
.B(n_520),
.Y(n_643)
);

AND2x2_ASAP7_75t_SL g644 ( 
.A(n_589),
.B(n_476),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_608),
.B(n_484),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_563),
.B(n_434),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_612),
.B(n_484),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_607),
.B(n_520),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_617),
.B(n_484),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_609),
.B(n_484),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_SL g651 ( 
.A(n_630),
.B(n_484),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_549),
.B(n_500),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_562),
.B(n_500),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_555),
.B(n_500),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_593),
.B(n_521),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_590),
.B(n_505),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_593),
.B(n_476),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_558),
.B(n_500),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_590),
.B(n_500),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_568),
.B(n_574),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_573),
.B(n_594),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_567),
.B(n_516),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_SL g663 ( 
.A(n_552),
.B(n_516),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_567),
.B(n_516),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_572),
.B(n_516),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_585),
.B(n_516),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_SL g667 ( 
.A(n_579),
.B(n_545),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_583),
.B(n_495),
.Y(n_668)
);

AND2x4_ASAP7_75t_L g669 ( 
.A(n_593),
.B(n_505),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_613),
.B(n_495),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_613),
.B(n_495),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_620),
.B(n_541),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_553),
.B(n_541),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_593),
.B(n_541),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_602),
.B(n_542),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g676 ( 
.A(n_546),
.B(n_542),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_595),
.B(n_542),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_618),
.B(n_529),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_625),
.B(n_614),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_550),
.B(n_434),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_551),
.B(n_434),
.Y(n_681)
);

NAND2xp33_ASAP7_75t_SL g682 ( 
.A(n_554),
.B(n_207),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_556),
.B(n_436),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_640),
.B(n_577),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_560),
.B(n_537),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_640),
.B(n_529),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_640),
.B(n_534),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_577),
.B(n_534),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_SL g689 ( 
.A(n_564),
.B(n_207),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_610),
.B(n_536),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_565),
.B(n_536),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_566),
.B(n_537),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_569),
.B(n_432),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_570),
.B(n_251),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_597),
.B(n_600),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_SL g696 ( 
.A(n_633),
.B(n_251),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_605),
.B(n_432),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_601),
.B(n_274),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_587),
.B(n_274),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_599),
.B(n_615),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_571),
.B(n_610),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_637),
.B(n_275),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_637),
.B(n_275),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_627),
.B(n_431),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_604),
.B(n_276),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_557),
.B(n_431),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_627),
.B(n_276),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_580),
.B(n_431),
.Y(n_708)
);

NAND2xp33_ASAP7_75t_SL g709 ( 
.A(n_633),
.B(n_280),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_622),
.B(n_280),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_636),
.B(n_406),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_580),
.B(n_584),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_639),
.B(n_281),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_632),
.B(n_281),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_634),
.B(n_283),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_588),
.B(n_283),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_SL g717 ( 
.A(n_611),
.B(n_229),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_591),
.B(n_233),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_592),
.B(n_407),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_596),
.B(n_234),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_626),
.B(n_236),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_623),
.B(n_237),
.Y(n_722)
);

NAND2xp33_ASAP7_75t_SL g723 ( 
.A(n_611),
.B(n_239),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_631),
.B(n_244),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_635),
.B(n_598),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_544),
.B(n_245),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_605),
.B(n_4),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_SL g728 ( 
.A(n_575),
.B(n_247),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_578),
.B(n_249),
.Y(n_729)
);

XNOR2xp5_ASAP7_75t_L g730 ( 
.A(n_547),
.B(n_254),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_581),
.B(n_257),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_SL g732 ( 
.A(n_619),
.B(n_258),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_641),
.B(n_259),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_SL g734 ( 
.A(n_606),
.B(n_616),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_606),
.B(n_260),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_641),
.B(n_263),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_616),
.B(n_264),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_708),
.A2(n_407),
.B(n_412),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_695),
.A2(n_559),
.B(n_629),
.Y(n_739)
);

OAI21x1_ASAP7_75t_L g740 ( 
.A1(n_693),
.A2(n_420),
.B(n_412),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_646),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_712),
.Y(n_742)
);

BUFx2_ASAP7_75t_SL g743 ( 
.A(n_660),
.Y(n_743)
);

A2O1A1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_661),
.A2(n_638),
.B(n_624),
.C(n_621),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_656),
.Y(n_745)
);

AO21x2_ASAP7_75t_L g746 ( 
.A1(n_733),
.A2(n_624),
.B(n_621),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_648),
.B(n_603),
.Y(n_747)
);

OAI22x1_ASAP7_75t_L g748 ( 
.A1(n_730),
.A2(n_727),
.B1(n_548),
.B2(n_547),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_656),
.B(n_586),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_R g750 ( 
.A(n_669),
.B(n_548),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_643),
.B(n_603),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_706),
.A2(n_628),
.B(n_301),
.Y(n_752)
);

AOI21xp5_ASAP7_75t_L g753 ( 
.A1(n_676),
.A2(n_628),
.B(n_303),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_675),
.A2(n_267),
.B(n_270),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_669),
.B(n_582),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_684),
.B(n_582),
.Y(n_756)
);

OAI21x1_ASAP7_75t_SL g757 ( 
.A1(n_685),
.A2(n_407),
.B(n_412),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_663),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_725),
.A2(n_413),
.B(n_420),
.Y(n_759)
);

AND3x4_ASAP7_75t_L g760 ( 
.A(n_711),
.B(n_561),
.C(n_6),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_680),
.B(n_561),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_642),
.A2(n_299),
.B(n_286),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_651),
.Y(n_763)
);

OAI21x1_ASAP7_75t_L g764 ( 
.A1(n_653),
.A2(n_420),
.B(n_418),
.Y(n_764)
);

AOI21x1_ASAP7_75t_SL g765 ( 
.A1(n_737),
.A2(n_5),
.B(n_6),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_665),
.A2(n_418),
.B(n_413),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_699),
.B(n_7),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_681),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_652),
.A2(n_297),
.B(n_290),
.Y(n_769)
);

OAI21x1_ASAP7_75t_L g770 ( 
.A1(n_690),
.A2(n_418),
.B(n_413),
.Y(n_770)
);

OAI22x1_ASAP7_75t_L g771 ( 
.A1(n_688),
.A2(n_273),
.B1(n_296),
.B2(n_306),
.Y(n_771)
);

NAND2x1_ASAP7_75t_L g772 ( 
.A(n_711),
.B(n_411),
.Y(n_772)
);

OAI21x1_ASAP7_75t_SL g773 ( 
.A1(n_683),
.A2(n_7),
.B(n_8),
.Y(n_773)
);

CKINVDCx6p67_ASAP7_75t_R g774 ( 
.A(n_694),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_719),
.Y(n_775)
);

AND3x2_ASAP7_75t_L g776 ( 
.A(n_697),
.B(n_8),
.C(n_10),
.Y(n_776)
);

AOI221xp5_ASAP7_75t_SL g777 ( 
.A1(n_698),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_777)
);

INVx3_ASAP7_75t_SL g778 ( 
.A(n_714),
.Y(n_778)
);

INVx5_ASAP7_75t_L g779 ( 
.A(n_704),
.Y(n_779)
);

OAI21x1_ASAP7_75t_L g780 ( 
.A1(n_690),
.A2(n_82),
.B(n_186),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_734),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_672),
.A2(n_411),
.B(n_81),
.Y(n_782)
);

AO32x2_ASAP7_75t_L g783 ( 
.A1(n_735),
.A2(n_12),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_783)
);

AOI221x1_ASAP7_75t_L g784 ( 
.A1(n_732),
.A2(n_411),
.B1(n_17),
.B2(n_18),
.C(n_19),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_659),
.B(n_15),
.Y(n_785)
);

AND3x4_ASAP7_75t_L g786 ( 
.A(n_719),
.B(n_17),
.C(n_18),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_644),
.B(n_19),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_644),
.B(n_20),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_704),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_655),
.A2(n_677),
.A3(n_657),
.B(n_674),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_682),
.B(n_411),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_679),
.A2(n_96),
.B(n_185),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_667),
.A2(n_411),
.B(n_93),
.Y(n_793)
);

NAND3xp33_ASAP7_75t_L g794 ( 
.A(n_689),
.B(n_411),
.C(n_21),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_705),
.A2(n_701),
.B1(n_666),
.B2(n_716),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_SL g796 ( 
.A1(n_721),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_700),
.A2(n_97),
.B(n_182),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_718),
.B(n_22),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_645),
.A2(n_100),
.B(n_178),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_662),
.B(n_23),
.Y(n_800)
);

AOI211x1_ASAP7_75t_L g801 ( 
.A1(n_720),
.A2(n_710),
.B(n_713),
.C(n_654),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_647),
.A2(n_91),
.B(n_177),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_789),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_739),
.A2(n_692),
.B(n_691),
.Y(n_804)
);

OAI21x1_ASAP7_75t_L g805 ( 
.A1(n_738),
.A2(n_736),
.B(n_733),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_779),
.B(n_736),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_779),
.B(n_670),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_789),
.Y(n_808)
);

OAI21x1_ASAP7_75t_L g809 ( 
.A1(n_740),
.A2(n_649),
.B(n_724),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_779),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_764),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_768),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_790),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_SL g814 ( 
.A1(n_787),
.A2(n_722),
.B(n_668),
.C(n_678),
.Y(n_814)
);

AOI222xp33_ASAP7_75t_L g815 ( 
.A1(n_748),
.A2(n_709),
.B1(n_696),
.B2(n_658),
.C1(n_703),
.C2(n_702),
.Y(n_815)
);

INVx4_ASAP7_75t_L g816 ( 
.A(n_763),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_766),
.Y(n_817)
);

AOI22xp5_ASAP7_75t_L g818 ( 
.A1(n_760),
.A2(n_707),
.B1(n_728),
.B2(n_664),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_752),
.A2(n_686),
.B(n_687),
.Y(n_819)
);

OAI21x1_ASAP7_75t_L g820 ( 
.A1(n_757),
.A2(n_650),
.B(n_673),
.Y(n_820)
);

AOI221xp5_ASAP7_75t_SL g821 ( 
.A1(n_798),
.A2(n_715),
.B1(n_729),
.B2(n_726),
.C(n_731),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_745),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_790),
.Y(n_823)
);

BUFx12f_ASAP7_75t_L g824 ( 
.A(n_749),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_759),
.A2(n_671),
.B(n_723),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_746),
.Y(n_826)
);

BUFx2_ASAP7_75t_SL g827 ( 
.A(n_758),
.Y(n_827)
);

AOI21x1_ASAP7_75t_L g828 ( 
.A1(n_791),
.A2(n_717),
.B(n_101),
.Y(n_828)
);

OAI21x1_ASAP7_75t_L g829 ( 
.A1(n_770),
.A2(n_90),
.B(n_175),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_744),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_742),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_SL g832 ( 
.A(n_767),
.B(n_25),
.C(n_26),
.Y(n_832)
);

INVx5_ASAP7_75t_L g833 ( 
.A(n_756),
.Y(n_833)
);

OAI21x1_ASAP7_75t_L g834 ( 
.A1(n_780),
.A2(n_102),
.B(n_173),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_795),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_746),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_787),
.B(n_788),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_741),
.B(n_29),
.Y(n_838)
);

AO21x2_ASAP7_75t_L g839 ( 
.A1(n_747),
.A2(n_105),
.B(n_172),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_747),
.Y(n_840)
);

AO21x2_ASAP7_75t_L g841 ( 
.A1(n_751),
.A2(n_78),
.B(n_171),
.Y(n_841)
);

NOR2xp67_ASAP7_75t_SL g842 ( 
.A(n_794),
.B(n_30),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_781),
.B(n_31),
.Y(n_843)
);

AOI21x1_ASAP7_75t_L g844 ( 
.A1(n_793),
.A2(n_106),
.B(n_169),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_792),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_743),
.B(n_35),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_800),
.Y(n_847)
);

AO21x2_ASAP7_75t_L g848 ( 
.A1(n_761),
.A2(n_108),
.B(n_168),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_781),
.B(n_36),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_788),
.A2(n_786),
.B1(n_801),
.B2(n_774),
.Y(n_850)
);

OA21x2_ASAP7_75t_L g851 ( 
.A1(n_784),
.A2(n_77),
.B(n_166),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_800),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_772),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_783),
.Y(n_854)
);

NOR2x1_ASAP7_75t_R g855 ( 
.A(n_785),
.B(n_37),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_775),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_813),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_811),
.Y(n_858)
);

AOI21xp33_ASAP7_75t_L g859 ( 
.A1(n_842),
.A2(n_794),
.B(n_777),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_813),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_840),
.B(n_761),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_823),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_805),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_823),
.Y(n_864)
);

NOR2x1_ASAP7_75t_R g865 ( 
.A(n_827),
.B(n_755),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_826),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_827),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_854),
.B(n_783),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_805),
.A2(n_765),
.B(n_782),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_826),
.Y(n_870)
);

AO21x2_ASAP7_75t_L g871 ( 
.A1(n_854),
.A2(n_773),
.B(n_795),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_815),
.A2(n_776),
.B1(n_771),
.B2(n_778),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_845),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_845),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_836),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_840),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_806),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_812),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_812),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_811),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_847),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_852),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_852),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_831),
.Y(n_885)
);

HB1xp67_ASAP7_75t_L g886 ( 
.A(n_816),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_816),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_831),
.B(n_777),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_837),
.B(n_753),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_839),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_811),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_843),
.B(n_783),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_839),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_839),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_817),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_848),
.Y(n_896)
);

HB1xp67_ASAP7_75t_L g897 ( 
.A(n_816),
.Y(n_897)
);

AO21x1_ASAP7_75t_SL g898 ( 
.A1(n_804),
.A2(n_796),
.B(n_797),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_848),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_843),
.B(n_37),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_848),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_816),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_841),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_841),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_841),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_819),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_806),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_809),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_878),
.Y(n_909)
);

XNOR2xp5_ASAP7_75t_L g910 ( 
.A(n_900),
.B(n_850),
.Y(n_910)
);

NAND2xp33_ASAP7_75t_R g911 ( 
.A(n_900),
.B(n_832),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_SL g912 ( 
.A(n_886),
.B(n_842),
.Y(n_912)
);

BUFx12f_ASAP7_75t_L g913 ( 
.A(n_900),
.Y(n_913)
);

XNOR2xp5_ASAP7_75t_L g914 ( 
.A(n_872),
.B(n_822),
.Y(n_914)
);

NAND2xp33_ASAP7_75t_R g915 ( 
.A(n_892),
.B(n_846),
.Y(n_915)
);

XNOR2xp5_ASAP7_75t_L g916 ( 
.A(n_872),
.B(n_822),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_878),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_R g918 ( 
.A(n_867),
.B(n_824),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_879),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_R g920 ( 
.A(n_867),
.B(n_824),
.Y(n_920)
);

XNOR2xp5_ASAP7_75t_L g921 ( 
.A(n_892),
.B(n_818),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_863),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_879),
.B(n_849),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_883),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_SL g925 ( 
.A(n_886),
.B(n_849),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_880),
.Y(n_926)
);

INVxp67_ASAP7_75t_L g927 ( 
.A(n_883),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_887),
.B(n_810),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_R g929 ( 
.A(n_887),
.B(n_750),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_885),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_876),
.B(n_833),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_877),
.B(n_833),
.Y(n_932)
);

NAND2xp33_ASAP7_75t_R g933 ( 
.A(n_892),
.B(n_851),
.Y(n_933)
);

NOR2x1_ASAP7_75t_L g934 ( 
.A(n_882),
.B(n_803),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_880),
.B(n_833),
.Y(n_935)
);

NAND2xp33_ASAP7_75t_R g936 ( 
.A(n_868),
.B(n_851),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_882),
.Y(n_937)
);

CKINVDCx8_ASAP7_75t_R g938 ( 
.A(n_863),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_907),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_884),
.B(n_833),
.Y(n_940)
);

BUFx10_ASAP7_75t_L g941 ( 
.A(n_884),
.Y(n_941)
);

INVxp67_ASAP7_75t_L g942 ( 
.A(n_907),
.Y(n_942)
);

XOR2xp5_ASAP7_75t_L g943 ( 
.A(n_885),
.B(n_818),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_R g944 ( 
.A(n_887),
.B(n_810),
.Y(n_944)
);

NAND2xp33_ASAP7_75t_R g945 ( 
.A(n_868),
.B(n_851),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_876),
.B(n_856),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_919),
.B(n_862),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_930),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_924),
.B(n_927),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_946),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_922),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_922),
.B(n_877),
.Y(n_952)
);

AOI22xp33_ASAP7_75t_L g953 ( 
.A1(n_921),
.A2(n_833),
.B1(n_859),
.B2(n_861),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_909),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_938),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_922),
.B(n_858),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_917),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_926),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_923),
.B(n_862),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_923),
.B(n_868),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_937),
.Y(n_961)
);

OR2x2_ASAP7_75t_L g962 ( 
.A(n_931),
.B(n_857),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_858),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_941),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_940),
.B(n_858),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_939),
.B(n_890),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_931),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_942),
.B(n_857),
.Y(n_968)
);

INVxp67_ASAP7_75t_SL g969 ( 
.A(n_936),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_941),
.B(n_906),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_944),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_934),
.B(n_871),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_932),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_945),
.Y(n_974)
);

OAI221xp5_ASAP7_75t_SL g975 ( 
.A1(n_910),
.A2(n_835),
.B1(n_830),
.B2(n_855),
.C(n_838),
.Y(n_975)
);

OR2x2_ASAP7_75t_L g976 ( 
.A(n_925),
.B(n_860),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_943),
.B(n_897),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_918),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_920),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_928),
.B(n_897),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_932),
.Y(n_981)
);

NAND2x1p5_ASAP7_75t_L g982 ( 
.A(n_933),
.B(n_877),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_SL g983 ( 
.A1(n_914),
.A2(n_859),
.B(n_888),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_912),
.B(n_902),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_913),
.B(n_906),
.Y(n_985)
);

OAI222xp33_ASAP7_75t_L g986 ( 
.A1(n_916),
.A2(n_833),
.B1(n_888),
.B2(n_861),
.C1(n_806),
.C2(n_889),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_957),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_967),
.B(n_902),
.Y(n_988)
);

INVx1_ASAP7_75t_SL g989 ( 
.A(n_949),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_957),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_969),
.B(n_863),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_982),
.B(n_877),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_969),
.B(n_963),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_963),
.B(n_863),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_978),
.B(n_979),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_960),
.B(n_871),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_948),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_971),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_971),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_963),
.B(n_863),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_955),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_967),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_959),
.B(n_871),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_955),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_957),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_950),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_958),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_959),
.B(n_871),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_958),
.Y(n_1009)
);

NOR3xp33_ASAP7_75t_L g1010 ( 
.A(n_975),
.B(n_855),
.C(n_821),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_958),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_993),
.B(n_974),
.Y(n_1012)
);

AND2x4_ASAP7_75t_SL g1013 ( 
.A(n_1006),
.B(n_973),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_987),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_992),
.B(n_974),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1002),
.B(n_950),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_998),
.B(n_973),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_987),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1002),
.B(n_949),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_990),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_998),
.B(n_999),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_989),
.B(n_960),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_997),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_989),
.B(n_962),
.Y(n_1024)
);

OR2x2_ASAP7_75t_L g1025 ( 
.A(n_996),
.B(n_962),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_990),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_996),
.B(n_1003),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_1003),
.B(n_947),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_999),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_1001),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_1008),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1005),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1016),
.B(n_993),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1012),
.A2(n_983),
.B1(n_1010),
.B2(n_915),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1012),
.B(n_1001),
.Y(n_1035)
);

OAI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1015),
.A2(n_983),
.B1(n_982),
.B2(n_992),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1021),
.B(n_1001),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_1015),
.A2(n_1010),
.B1(n_911),
.B2(n_982),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1019),
.B(n_1024),
.Y(n_1039)
);

OAI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_1015),
.A2(n_982),
.B1(n_992),
.B2(n_1008),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_1015),
.A2(n_985),
.B1(n_972),
.B2(n_992),
.Y(n_1041)
);

AO221x2_ASAP7_75t_L g1042 ( 
.A1(n_1021),
.A2(n_977),
.B1(n_986),
.B2(n_984),
.C(n_988),
.Y(n_1042)
);

INVx3_ASAP7_75t_SL g1043 ( 
.A(n_1021),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1039),
.B(n_1028),
.Y(n_1044)
);

NAND2xp33_ASAP7_75t_L g1045 ( 
.A(n_1034),
.B(n_978),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1033),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1035),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_1043),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1037),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1042),
.B(n_1029),
.Y(n_1050)
);

XNOR2xp5_ASAP7_75t_L g1051 ( 
.A(n_1048),
.B(n_1038),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_1045),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1044),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1053),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1054),
.B(n_1049),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1052),
.B(n_1050),
.Y(n_1057)
);

INVx1_ASAP7_75t_SL g1058 ( 
.A(n_1051),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1051),
.A2(n_1042),
.B1(n_1045),
.B2(n_1036),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1053),
.B(n_1031),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1053),
.Y(n_1061)
);

INVx2_ASAP7_75t_SL g1062 ( 
.A(n_1051),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_1053),
.B(n_1028),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1052),
.B(n_1030),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_1053),
.B(n_995),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1063),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1055),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1061),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1060),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1060),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1056),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1065),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1065),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1064),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_1062),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1058),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1058),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_1057),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1059),
.Y(n_1079)
);

INVxp33_ASAP7_75t_SL g1080 ( 
.A(n_1058),
.Y(n_1080)
);

INVxp33_ASAP7_75t_SL g1081 ( 
.A(n_1058),
.Y(n_1081)
);

NAND4xp25_ASAP7_75t_L g1082 ( 
.A(n_1074),
.B(n_975),
.C(n_979),
.D(n_1041),
.Y(n_1082)
);

OAI211xp5_ASAP7_75t_L g1083 ( 
.A1(n_1075),
.A2(n_984),
.B(n_988),
.C(n_1004),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1080),
.A2(n_1031),
.B(n_1040),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_1081),
.B(n_1027),
.Y(n_1085)
);

NAND4xp25_ASAP7_75t_L g1086 ( 
.A(n_1075),
.B(n_1017),
.C(n_1004),
.D(n_964),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1077),
.B(n_1025),
.Y(n_1087)
);

NAND4xp25_ASAP7_75t_L g1088 ( 
.A(n_1072),
.B(n_1017),
.C(n_1004),
.D(n_964),
.Y(n_1088)
);

AOI211xp5_ASAP7_75t_L g1089 ( 
.A1(n_1078),
.A2(n_985),
.B(n_991),
.C(n_977),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1076),
.B(n_1017),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1077),
.Y(n_1091)
);

AND3x2_ASAP7_75t_L g1092 ( 
.A(n_1073),
.B(n_1068),
.C(n_1067),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1066),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_SL g1094 ( 
.A1(n_1071),
.A2(n_1013),
.B(n_985),
.Y(n_1094)
);

NOR3xp33_ASAP7_75t_L g1095 ( 
.A(n_1069),
.B(n_1022),
.C(n_808),
.Y(n_1095)
);

OAI21xp33_ASAP7_75t_L g1096 ( 
.A1(n_1070),
.A2(n_1013),
.B(n_991),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1079),
.B(n_1014),
.Y(n_1097)
);

AOI211xp5_ASAP7_75t_L g1098 ( 
.A1(n_1078),
.A2(n_972),
.B(n_986),
.C(n_814),
.Y(n_1098)
);

AOI221xp5_ASAP7_75t_L g1099 ( 
.A1(n_1080),
.A2(n_953),
.B1(n_1026),
.B2(n_1020),
.C(n_1018),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1080),
.B(n_964),
.Y(n_1100)
);

OAI22xp33_ASAP7_75t_R g1101 ( 
.A1(n_1091),
.A2(n_951),
.B1(n_947),
.B2(n_976),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_851),
.B(n_976),
.C(n_1032),
.Y(n_1102)
);

OAI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1084),
.A2(n_1023),
.B1(n_992),
.B2(n_951),
.C(n_955),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1092),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1090),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1085),
.A2(n_1100),
.B(n_1087),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_1097),
.A2(n_1023),
.B(n_951),
.C(n_966),
.Y(n_1107)
);

OAI211xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1094),
.A2(n_980),
.B(n_39),
.C(n_41),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1086),
.Y(n_1109)
);

NAND3xp33_ASAP7_75t_SL g1110 ( 
.A(n_1089),
.B(n_929),
.C(n_762),
.Y(n_1110)
);

NOR4xp25_ASAP7_75t_L g1111 ( 
.A(n_1083),
.B(n_954),
.C(n_38),
.D(n_980),
.Y(n_1111)
);

OAI211xp5_ASAP7_75t_L g1112 ( 
.A1(n_1088),
.A2(n_1000),
.B(n_994),
.C(n_887),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_L g1113 ( 
.A1(n_1095),
.A2(n_871),
.B1(n_769),
.B2(n_893),
.C(n_894),
.Y(n_1113)
);

OAI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1082),
.A2(n_970),
.B(n_1000),
.Y(n_1114)
);

AOI221xp5_ASAP7_75t_L g1115 ( 
.A1(n_1099),
.A2(n_894),
.B1(n_893),
.B2(n_890),
.C(n_904),
.Y(n_1115)
);

AOI221xp5_ASAP7_75t_L g1116 ( 
.A1(n_1098),
.A2(n_1096),
.B1(n_903),
.B2(n_904),
.C(n_889),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1092),
.B(n_994),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_1104),
.B(n_38),
.Y(n_1118)
);

AOI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1101),
.A2(n_1011),
.B1(n_1009),
.B2(n_1007),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_SL g1120 ( 
.A(n_1105),
.B(n_810),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1106),
.Y(n_1121)
);

NOR2x1_ASAP7_75t_L g1122 ( 
.A(n_1108),
.B(n_803),
.Y(n_1122)
);

XNOR2xp5_ASAP7_75t_L g1123 ( 
.A(n_1111),
.B(n_966),
.Y(n_1123)
);

NOR2x1p5_ASAP7_75t_L g1124 ( 
.A(n_1109),
.B(n_1117),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_1109),
.B(n_970),
.Y(n_1125)
);

NAND4xp75_ASAP7_75t_L g1126 ( 
.A(n_1116),
.B(n_970),
.C(n_802),
.D(n_799),
.Y(n_1126)
);

NAND4xp75_ASAP7_75t_L g1127 ( 
.A(n_1113),
.B(n_754),
.C(n_1009),
.D(n_1007),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1110),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1103),
.Y(n_1129)
);

XOR2xp5_ASAP7_75t_L g1130 ( 
.A(n_1114),
.B(n_981),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1112),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1107),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1102),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1115),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1104),
.Y(n_1135)
);

NAND4xp75_ASAP7_75t_L g1136 ( 
.A(n_1106),
.B(n_1011),
.C(n_1005),
.D(n_956),
.Y(n_1136)
);

NOR2x1_ASAP7_75t_L g1137 ( 
.A(n_1104),
.B(n_803),
.Y(n_1137)
);

NAND2x1p5_ASAP7_75t_L g1138 ( 
.A(n_1104),
.B(n_803),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1104),
.Y(n_1139)
);

XNOR2x1_ASAP7_75t_L g1140 ( 
.A(n_1104),
.B(n_807),
.Y(n_1140)
);

NOR2x1_ASAP7_75t_L g1141 ( 
.A(n_1104),
.B(n_808),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1135),
.B(n_954),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_R g1143 ( 
.A(n_1121),
.B(n_808),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1139),
.B(n_961),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1118),
.B(n_961),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_R g1146 ( 
.A(n_1128),
.B(n_808),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1137),
.B(n_1138),
.Y(n_1147)
);

NAND2xp33_ASAP7_75t_L g1148 ( 
.A(n_1124),
.B(n_887),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_1120),
.B(n_853),
.C(n_968),
.Y(n_1149)
);

NAND2xp33_ASAP7_75t_SL g1150 ( 
.A(n_1124),
.B(n_968),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1122),
.B(n_961),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_SL g1152 ( 
.A(n_1131),
.B(n_853),
.Y(n_1152)
);

NAND2xp33_ASAP7_75t_SL g1153 ( 
.A(n_1131),
.B(n_853),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_R g1154 ( 
.A(n_1133),
.B(n_44),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_R g1155 ( 
.A(n_1123),
.B(n_45),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1141),
.B(n_853),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_1141),
.B(n_853),
.C(n_807),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1132),
.B(n_807),
.C(n_863),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_1122),
.B(n_863),
.Y(n_1159)
);

NAND2xp33_ASAP7_75t_SL g1160 ( 
.A(n_1125),
.B(n_973),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_1129),
.B(n_807),
.C(n_863),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_R g1162 ( 
.A(n_1134),
.B(n_1140),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_R g1163 ( 
.A(n_1127),
.B(n_1126),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1119),
.B(n_973),
.Y(n_1164)
);

NAND2xp33_ASAP7_75t_SL g1165 ( 
.A(n_1136),
.B(n_956),
.Y(n_1165)
);

AOI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1150),
.A2(n_1130),
.B1(n_952),
.B2(n_903),
.Y(n_1166)
);

NAND5xp2_ASAP7_75t_L g1167 ( 
.A(n_1142),
.B(n_844),
.C(n_828),
.D(n_956),
.E(n_965),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1147),
.Y(n_1168)
);

XOR2xp5_ASAP7_75t_L g1169 ( 
.A(n_1144),
.B(n_46),
.Y(n_1169)
);

XNOR2xp5_ASAP7_75t_L g1170 ( 
.A(n_1145),
.B(n_952),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_1148),
.B(n_997),
.C(n_952),
.Y(n_1171)
);

XNOR2x1_ASAP7_75t_L g1172 ( 
.A(n_1161),
.B(n_834),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_1155),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_SL g1174 ( 
.A1(n_1163),
.A2(n_952),
.B1(n_981),
.B2(n_898),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_1162),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1156),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1154),
.B(n_997),
.Y(n_1177)
);

NAND4xp25_ASAP7_75t_L g1178 ( 
.A(n_1160),
.B(n_965),
.C(n_981),
.D(n_908),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1152),
.B(n_965),
.C(n_908),
.Y(n_1179)
);

INVx5_ASAP7_75t_L g1180 ( 
.A(n_1146),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1164),
.B(n_869),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1151),
.Y(n_1182)
);

XNOR2xp5_ASAP7_75t_L g1183 ( 
.A(n_1153),
.B(n_828),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1159),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1165),
.A2(n_905),
.B1(n_899),
.B2(n_901),
.Y(n_1185)
);

AOI211xp5_ASAP7_75t_L g1186 ( 
.A1(n_1143),
.A2(n_869),
.B(n_865),
.C(n_834),
.Y(n_1186)
);

XNOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1158),
.B(n_844),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1175),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1180),
.B(n_1168),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1180),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1173),
.Y(n_1191)
);

AOI222xp33_ASAP7_75t_L g1192 ( 
.A1(n_1182),
.A2(n_1149),
.B1(n_1157),
.B2(n_905),
.C1(n_901),
.C2(n_899),
.Y(n_1192)
);

AND2x2_ASAP7_75t_SL g1193 ( 
.A(n_1176),
.B(n_908),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1184),
.A2(n_869),
.B(n_829),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1169),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1170),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1172),
.A2(n_905),
.B1(n_901),
.B2(n_899),
.Y(n_1197)
);

AOI32xp33_ASAP7_75t_L g1198 ( 
.A1(n_1186),
.A2(n_899),
.A3(n_901),
.B1(n_905),
.B2(n_896),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1174),
.A2(n_829),
.B(n_820),
.Y(n_1199)
);

OA22x2_ASAP7_75t_L g1200 ( 
.A1(n_1166),
.A2(n_820),
.B1(n_908),
.B2(n_809),
.Y(n_1200)
);

OAI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1178),
.A2(n_896),
.B1(n_948),
.B2(n_873),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1181),
.B(n_819),
.Y(n_1202)
);

OA22x2_ASAP7_75t_L g1203 ( 
.A1(n_1188),
.A2(n_1177),
.B1(n_1183),
.B2(n_1185),
.Y(n_1203)
);

OAI22x1_ASAP7_75t_L g1204 ( 
.A1(n_1189),
.A2(n_1190),
.B1(n_1196),
.B2(n_1191),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1195),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1193),
.B(n_1187),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1197),
.A2(n_1179),
.B1(n_1171),
.B2(n_1167),
.Y(n_1207)
);

AOI22x1_ASAP7_75t_L g1208 ( 
.A1(n_1199),
.A2(n_51),
.B1(n_53),
.B2(n_60),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_1200),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1198),
.B(n_62),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1202),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1192),
.B(n_1201),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_L g1213 ( 
.A1(n_1194),
.A2(n_874),
.B(n_873),
.Y(n_1213)
);

OAI22x1_ASAP7_75t_L g1214 ( 
.A1(n_1188),
.A2(n_948),
.B1(n_896),
.B2(n_898),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_1188),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1188),
.Y(n_1216)
);

AO22x1_ASAP7_75t_L g1217 ( 
.A1(n_1188),
.A2(n_898),
.B1(n_874),
.B2(n_873),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1209),
.A2(n_870),
.B1(n_866),
.B2(n_873),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1206),
.A2(n_870),
.B1(n_866),
.B2(n_873),
.Y(n_1219)
);

AOI31xp33_ASAP7_75t_L g1220 ( 
.A1(n_1215),
.A2(n_865),
.A3(n_65),
.B(n_67),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1207),
.A2(n_874),
.B1(n_860),
.B2(n_864),
.Y(n_1221)
);

AOI31xp33_ASAP7_75t_L g1222 ( 
.A1(n_1216),
.A2(n_63),
.A3(n_69),
.B(n_70),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1203),
.A2(n_1212),
.B1(n_1210),
.B2(n_1205),
.Y(n_1223)
);

AOI31xp33_ASAP7_75t_L g1224 ( 
.A1(n_1211),
.A2(n_75),
.A3(n_112),
.B(n_113),
.Y(n_1224)
);

AOI31xp33_ASAP7_75t_L g1225 ( 
.A1(n_1204),
.A2(n_123),
.A3(n_126),
.B(n_128),
.Y(n_1225)
);

AOI31xp33_ASAP7_75t_L g1226 ( 
.A1(n_1208),
.A2(n_133),
.A3(n_134),
.B(n_137),
.Y(n_1226)
);

AOI31xp33_ASAP7_75t_L g1227 ( 
.A1(n_1213),
.A2(n_138),
.A3(n_140),
.B(n_141),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1223),
.A2(n_1214),
.B1(n_1217),
.B2(n_874),
.Y(n_1228)
);

AOI211xp5_ASAP7_75t_L g1229 ( 
.A1(n_1225),
.A2(n_825),
.B(n_150),
.C(n_151),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1218),
.A2(n_874),
.B1(n_825),
.B2(n_864),
.Y(n_1230)
);

AOI221x1_ASAP7_75t_L g1231 ( 
.A1(n_1227),
.A2(n_146),
.B1(n_163),
.B2(n_184),
.C(n_895),
.Y(n_1231)
);

AO22x2_ASAP7_75t_L g1232 ( 
.A1(n_1226),
.A2(n_1222),
.B1(n_1224),
.B2(n_1220),
.Y(n_1232)
);

AOI211xp5_ASAP7_75t_L g1233 ( 
.A1(n_1221),
.A2(n_895),
.B(n_891),
.C(n_881),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1232),
.Y(n_1234)
);

OAI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1231),
.A2(n_1219),
.B1(n_891),
.B2(n_881),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1229),
.A2(n_891),
.B(n_881),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1228),
.A2(n_1230),
.B1(n_1233),
.B2(n_895),
.Y(n_1237)
);

XNOR2xp5_ASAP7_75t_L g1238 ( 
.A(n_1234),
.B(n_875),
.Y(n_1238)
);

OAI221xp5_ASAP7_75t_L g1239 ( 
.A1(n_1238),
.A2(n_1237),
.B1(n_1236),
.B2(n_1235),
.C(n_895),
.Y(n_1239)
);

AOI211xp5_ASAP7_75t_L g1240 ( 
.A1(n_1239),
.A2(n_895),
.B(n_891),
.C(n_881),
.Y(n_1240)
);


endmodule