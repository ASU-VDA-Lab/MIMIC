module fake_jpeg_816_n_175 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_175);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_175;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_1),
.B(n_40),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_67),
.Y(n_72)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_46),
.Y(n_66)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_21),
.B1(n_43),
.B2(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2x1_ASAP7_75t_SL g73 ( 
.A(n_68),
.B(n_46),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_60),
.B1(n_66),
.B2(n_56),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_79),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_50),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_72),
.A2(n_57),
.B1(n_60),
.B2(n_54),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_47),
.B1(n_46),
.B2(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_54),
.B1(n_56),
.B2(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_59),
.B1(n_69),
.B2(n_6),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_45),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_61),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_91),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_109),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_115),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_55),
.B(n_53),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_9),
.B(n_10),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_75),
.B1(n_59),
.B2(n_47),
.Y(n_102)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_110),
.B(n_26),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_95),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_114),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_69),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_59),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_94),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_96),
.B1(n_94),
.B2(n_83),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_100),
.B1(n_14),
.B2(n_15),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_8),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_125),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_123),
.Y(n_136)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_95),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_8),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_9),
.Y(n_127)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_132),
.B(n_13),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_27),
.C(n_38),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_30),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g132 ( 
.A(n_107),
.B(n_10),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_28),
.Y(n_133)
);

OAI321xp33_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_31),
.A3(n_35),
.B1(n_18),
.B2(n_19),
.C(n_23),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_11),
.B(n_12),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_100),
.B(n_105),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_135),
.A2(n_16),
.B1(n_29),
.B2(n_32),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_143),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_135),
.B1(n_129),
.B2(n_132),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_147),
.B(n_149),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_15),
.B(n_16),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_148),
.A2(n_133),
.B(n_34),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_130),
.B1(n_121),
.B2(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_158),
.B(n_146),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_33),
.B(n_44),
.C(n_139),
.D(n_142),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_148),
.B(n_137),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_154),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_155),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_163),
.A2(n_164),
.B(n_138),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_162),
.Y(n_169)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_159),
.B(n_153),
.C(n_152),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_160),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_170),
.B(n_169),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_168),
.B(n_158),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_149),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_157),
.B(n_150),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_144),
.Y(n_175)
);


endmodule