module fake_jpeg_16261_n_86 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_86);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_86;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_24),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

CKINVDCx11_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_1),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_3),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_29),
.Y(n_44)
);

AOI32xp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_39),
.A2(n_33),
.B1(n_32),
.B2(n_30),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_47),
.Y(n_57)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_52),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_3),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_55),
.B(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_60),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_4),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_7),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_63),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_64),
.B(n_65),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_13),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_49),
.A2(n_14),
.B1(n_15),
.B2(n_17),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_20),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_21),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g68 ( 
.A(n_58),
.Y(n_68)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

CKINVDCx10_ASAP7_75t_R g71 ( 
.A(n_55),
.Y(n_71)
);

INVxp33_ASAP7_75t_SL g76 ( 
.A(n_71),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_73),
.A2(n_74),
.B1(n_57),
.B2(n_25),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_77),
.B(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_75),
.B(n_70),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_72),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_81),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_82),
.B(n_76),
.Y(n_83)
);

OAI211xp5_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_76),
.B(n_79),
.C(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_23),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g86 ( 
.A(n_85),
.Y(n_86)
);


endmodule