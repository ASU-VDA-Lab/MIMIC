module fake_jpeg_20808_n_271 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_271);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_271;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_18),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_40),
.B(n_23),
.Y(n_46)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_42),
.B(n_31),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_48),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_47),
.B(n_55),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_19),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_50),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_20),
.B1(n_34),
.B2(n_29),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g84 ( 
.A(n_58),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_25),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_63),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_56),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_27),
.B1(n_29),
.B2(n_34),
.Y(n_64)
);

OAI22x1_ASAP7_75t_L g97 ( 
.A1(n_64),
.A2(n_37),
.B1(n_36),
.B2(n_41),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_46),
.B(n_40),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_41),
.Y(n_115)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_78),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_28),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_79),
.Y(n_109)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_47),
.A2(n_20),
.B1(n_29),
.B2(n_42),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_90),
.B1(n_72),
.B2(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_83),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_40),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g118 ( 
.A(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_39),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_39),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_94),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_91),
.Y(n_117)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_32),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_41),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_58),
.B1(n_84),
.B2(n_75),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_24),
.B(n_22),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_104),
.B(n_115),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_38),
.A3(n_24),
.B1(n_27),
.B2(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_108),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_41),
.B(n_38),
.Y(n_104)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_113),
.Y(n_134)
);

AO22x2_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_41),
.B1(n_38),
.B2(n_49),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_119),
.B1(n_58),
.B2(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_36),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_81),
.A2(n_94),
.B(n_61),
.C(n_70),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_67),
.B(n_36),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_27),
.B1(n_38),
.B2(n_22),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_30),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_60),
.C(n_23),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_122),
.B(n_123),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_112),
.A2(n_61),
.B(n_87),
.C(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_131),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_129),
.A2(n_138),
.B1(n_147),
.B2(n_74),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_139),
.C(n_145),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_132),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_60),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_38),
.B1(n_85),
.B2(n_92),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_108),
.B1(n_76),
.B2(n_68),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_120),
.B(n_110),
.C(n_113),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_115),
.C(n_110),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_15),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g145 ( 
.A1(n_101),
.A2(n_30),
.B(n_13),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g146 ( 
.A(n_95),
.B(n_23),
.C(n_17),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_146),
.B(n_23),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_104),
.A2(n_75),
.B1(n_58),
.B2(n_91),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_114),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_95),
.B(n_30),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_149),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_150),
.B(n_151),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_127),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_161),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_159),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_140),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_164),
.B(n_173),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_115),
.B(n_99),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_112),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_52),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_99),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_133),
.B1(n_128),
.B2(n_137),
.C(n_135),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g204 ( 
.A1(n_181),
.A2(n_193),
.B(n_194),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_160),
.B1(n_159),
.B2(n_154),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_133),
.B(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_188),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_131),
.B(n_141),
.Y(n_188)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_146),
.CI(n_17),
.CON(n_190),
.SN(n_190)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_12),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_172),
.B(n_157),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_13),
.C(n_2),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_199),
.B1(n_154),
.B2(n_171),
.Y(n_215)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_150),
.B1(n_169),
.B2(n_160),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_148),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_162),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_202),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_168),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_206),
.Y(n_223)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_158),
.B(n_165),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_158),
.C(n_179),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_217),
.C(n_33),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_179),
.B(n_167),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_159),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_216),
.C(n_186),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_185),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_211),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_152),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_187),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_17),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_153),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_153),
.C(n_107),
.Y(n_217)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

OAI211xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_188),
.B(n_197),
.C(n_178),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_1),
.B(n_2),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_227),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_26),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_232),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_182),
.B1(n_187),
.B2(n_197),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_229),
.B1(n_89),
.B2(n_44),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_196),
.C(n_182),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_178),
.C(n_114),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_26),
.C(n_33),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_232),
.B(n_217),
.C(n_205),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_234),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_210),
.C(n_208),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_203),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_44),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_221),
.A2(n_218),
.B1(n_225),
.B2(n_204),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_1),
.B(n_5),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_37),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_1),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_242),
.A2(n_223),
.B(n_44),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_249),
.B1(n_239),
.B2(n_233),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_252),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_234),
.A2(n_26),
.B1(n_37),
.B2(n_3),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_248),
.Y(n_255)
);

AOI21x1_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_5),
.B(n_7),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_259),
.Y(n_264)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_260),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_235),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_254),
.B(n_247),
.C(n_235),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_248),
.B(n_236),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_246),
.C(n_258),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

AOI322xp5_ASAP7_75t_L g268 ( 
.A1(n_262),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_264),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_265),
.B1(n_10),
.B2(n_11),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_269),
.Y(n_271)
);


endmodule