module fake_jpeg_27740_n_24 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_24);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_24;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_9),
.B1(n_8),
.B2(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_16),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

NAND4xp25_ASAP7_75t_SL g18 ( 
.A(n_16),
.B(n_12),
.C(n_11),
.D(n_5),
.Y(n_18)
);

AO221x1_ASAP7_75t_L g20 ( 
.A1(n_18),
.A2(n_12),
.B1(n_4),
.B2(n_6),
.C(n_3),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_21),
.C(n_17),
.Y(n_22)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_15),
.B(n_14),
.C(n_6),
.D(n_4),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_23),
.A2(n_18),
.B(n_17),
.Y(n_24)
);


endmodule