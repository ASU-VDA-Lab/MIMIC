module fake_jpeg_11122_n_95 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_1),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_38),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_33),
.A2(n_17),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_50),
.Y(n_56)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_53),
.B(n_57),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_39),
.B1(n_42),
.B2(n_34),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_54),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_7),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_43),
.B1(n_35),
.B2(n_36),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_45),
.B1(n_35),
.B2(n_34),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_61),
.A2(n_20),
.B(n_23),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_1),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_71),
.Y(n_75)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_45),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_67),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_65),
.Y(n_76)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_3),
.C(n_6),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_70),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_19),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_79),
.A2(n_83),
.B(n_26),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_24),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_29),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_87),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_85),
.C(n_86),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_73),
.B(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_89),
.Y(n_92)
);

BUFx12f_ASAP7_75t_SL g93 ( 
.A(n_92),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_80),
.C(n_75),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_78),
.Y(n_95)
);


endmodule