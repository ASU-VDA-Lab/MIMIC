module real_jpeg_7729_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_1),
.A2(n_31),
.B1(n_34),
.B2(n_54),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_2),
.A2(n_31),
.B1(n_34),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_2),
.A2(n_25),
.B1(n_38),
.B2(n_71),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_71),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_3),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_4),
.A2(n_25),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_40),
.B1(n_48),
.B2(n_49),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_4),
.A2(n_31),
.B1(n_34),
.B2(n_40),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_31),
.B1(n_34),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_5),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_5),
.A2(n_48),
.B1(n_49),
.B2(n_75),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx6f_ASAP7_75t_SL g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_11),
.B(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_11),
.A2(n_25),
.B(n_59),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_11),
.A2(n_80),
.B1(n_93),
.B2(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_11),
.A2(n_34),
.B(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_11),
.B(n_34),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_45),
.B1(n_85),
.B2(n_146),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_13),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_14),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_25),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_15),
.A2(n_37),
.B1(n_93),
.B2(n_116),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_15),
.A2(n_31),
.B1(n_34),
.B2(n_37),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_15),
.A2(n_37),
.B1(n_48),
.B2(n_49),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_87),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_19),
.B(n_87),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_64),
.C(n_76),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_20),
.A2(n_21),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_42),
.B1(n_43),
.B2(n_63),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_35),
.B1(n_39),
.B2(n_41),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_23),
.A2(n_39),
.B1(n_41),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_24),
.A2(n_30),
.B1(n_36),
.B2(n_79),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_25),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_25),
.B(n_80),
.CON(n_79),
.SN(n_79)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_27),
.B(n_34),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_29),
.A2(n_31),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_66),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_41),
.B(n_80),
.Y(n_157)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_44),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_52),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_45),
.A2(n_47),
.B1(n_85),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_45),
.A2(n_85),
.B1(n_128),
.B2(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_45),
.B(n_80),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_53),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_46),
.A2(n_55),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_46),
.B(n_84),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_49),
.B1(n_66),
.B2(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_48),
.B(n_69),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_48),
.B(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_49),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_137)
);

BUFx24_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_55),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_56),
.B(n_61),
.C(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_57),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_111)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_58),
.A2(n_60),
.B(n_93),
.C(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_80),
.B(n_92),
.C(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_60),
.B(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_64),
.A2(n_76),
.B1(n_77),
.B2(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_64),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_70),
.B(n_72),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_65),
.A2(n_68),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_65),
.A2(n_68),
.B1(n_136),
.B2(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_65),
.A2(n_68),
.B1(n_70),
.B2(n_159),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_68),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_68),
.B(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_78),
.B(n_82),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_85),
.A2(n_130),
.B(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_93),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_111),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_108),
.B2(n_109),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_174),
.B(n_180),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_163),
.B(n_173),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_153),
.B(n_162),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_142),
.B(n_152),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_126),
.B(n_131),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_141),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_141),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_135),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_137),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_147),
.B(n_151),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_145),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_155),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_156),
.B(n_164),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.CI(n_160),
.CON(n_156),
.SN(n_156)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_171),
.B2(n_172),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_167),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_168),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_175),
.B(n_176),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);


endmodule