module fake_jpeg_13589_n_262 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_35),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_33),
.C(n_35),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_22),
.C(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_59),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_55),
.Y(n_100)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_34),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_62),
.Y(n_85)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_44),
.A2(n_24),
.B1(n_17),
.B2(n_20),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_40),
.B1(n_17),
.B2(n_39),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_17),
.B(n_26),
.C(n_25),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_17),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_75),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_25),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_31),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_78),
.A2(n_70),
.B1(n_17),
.B2(n_47),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_21),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_43),
.B1(n_24),
.B2(n_36),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_83),
.A2(n_20),
.B1(n_23),
.B2(n_32),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_21),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_24),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_94),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_89),
.A2(n_32),
.B1(n_30),
.B2(n_28),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_47),
.B(n_21),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_27),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_46),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_101),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_64),
.A2(n_39),
.B1(n_36),
.B2(n_40),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_98),
.A2(n_66),
.B1(n_36),
.B2(n_39),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_58),
.B(n_46),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_127),
.B1(n_91),
.B2(n_92),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_80),
.C(n_72),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_52),
.CI(n_90),
.CON(n_133),
.SN(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_100),
.Y(n_141)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_119),
.B1(n_120),
.B2(n_125),
.Y(n_134)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_116),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_20),
.B(n_52),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_117),
.A2(n_86),
.B(n_71),
.Y(n_147)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_16),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_16),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_94),
.A2(n_75),
.B1(n_88),
.B2(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_95),
.A2(n_23),
.B1(n_28),
.B2(n_32),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_92),
.B1(n_30),
.B2(n_91),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_30),
.B1(n_28),
.B2(n_55),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_85),
.A2(n_30),
.B1(n_28),
.B2(n_55),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_111),
.B(n_85),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_136),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_114),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_SL g172 ( 
.A(n_131),
.B(n_137),
.C(n_141),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_29),
.C(n_5),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_135),
.A2(n_126),
.B1(n_106),
.B2(n_122),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_111),
.B(n_90),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_138),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_100),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_97),
.B(n_96),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_143),
.A2(n_147),
.B(n_149),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_99),
.B(n_96),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_155),
.B1(n_102),
.B2(n_125),
.Y(n_158)
);

INVx8_ASAP7_75t_L g151 ( 
.A(n_106),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_153),
.Y(n_177)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_110),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_71),
.B1(n_99),
.B2(n_27),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_123),
.B1(n_118),
.B2(n_119),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_158),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_115),
.B(n_103),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_175),
.B(n_145),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_141),
.A2(n_127),
.B1(n_120),
.B2(n_115),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_155),
.B1(n_148),
.B2(n_131),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_145),
.B(n_129),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_145),
.B1(n_151),
.B2(n_139),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_146),
.A2(n_126),
.B1(n_113),
.B2(n_108),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_113),
.B1(n_29),
.B2(n_2),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_174),
.B1(n_176),
.B2(n_178),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_0),
.B(n_1),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_29),
.B1(n_1),
.B2(n_3),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_133),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_178),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_130),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_164),
.B(n_133),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_154),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_188),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_183),
.A2(n_191),
.B1(n_200),
.B2(n_176),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_157),
.B(n_168),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_194),
.C(n_199),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_177),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_196),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_197),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_169),
.A2(n_145),
.B1(n_142),
.B2(n_129),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_162),
.B(n_169),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_173),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_153),
.C(n_152),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_185),
.A2(n_171),
.B1(n_161),
.B2(n_174),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_204),
.A2(n_192),
.B1(n_191),
.B2(n_190),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_192),
.A2(n_167),
.B1(n_158),
.B2(n_160),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_170),
.C(n_166),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_209),
.C(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_166),
.C(n_156),
.Y(n_209)
);

AOI321xp33_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_172),
.A3(n_156),
.B1(n_159),
.B2(n_175),
.C(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_211),
.B(n_215),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_197),
.Y(n_227)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_156),
.C(n_15),
.Y(n_217)
);

INVx13_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_218),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_227),
.B1(n_211),
.B2(n_210),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_199),
.C(n_193),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_203),
.C(n_13),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_225),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_193),
.B(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_208),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_193),
.B1(n_15),
.B2(n_12),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_230),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_9),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_205),
.B1(n_204),
.B2(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_236),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_235),
.B(n_225),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_14),
.B(n_11),
.Y(n_240)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_240),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_229),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_242),
.B(n_246),
.Y(n_249)
);

BUFx12f_ASAP7_75t_SL g243 ( 
.A(n_234),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_233),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_220),
.C(n_222),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_251),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_220),
.C(n_235),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_252),
.B(n_240),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g258 ( 
.A1(n_253),
.A2(n_254),
.B(n_226),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_241),
.C(n_228),
.Y(n_254)
);

OAI221xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_243),
.B1(n_227),
.B2(n_245),
.C(n_240),
.Y(n_257)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_257),
.A2(n_258),
.A3(n_256),
.B1(n_238),
.B2(n_218),
.C1(n_226),
.C2(n_232),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_14),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

AO21x2_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_11),
.B(n_13),
.Y(n_262)
);


endmodule