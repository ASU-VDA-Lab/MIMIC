module fake_jpeg_26163_n_79 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_39),
.B(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_44),
.Y(n_58)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_45),
.B(n_46),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_57)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_14),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_15),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_57),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_44),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_68),
.B1(n_38),
.B2(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_35),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_34),
.C(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_36),
.C(n_64),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_56),
.C(n_55),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_72),
.A2(n_52),
.B1(n_20),
.B2(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_75),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_54),
.B1(n_57),
.B2(n_61),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_59),
.B(n_53),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);


endmodule