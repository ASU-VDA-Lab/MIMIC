module fake_ariane_227_n_851 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_851);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_851;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_176;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_481;
wire n_433;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_455;
wire n_429;
wire n_365;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_772;
wire n_741;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_37),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_121),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_90),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_106),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_48),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_52),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_143),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_85),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_6),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_8),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_28),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_23),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_30),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_69),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_22),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_0),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_5),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_163),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_119),
.Y(n_201)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_47),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_124),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_32),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_41),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_64),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_116),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_20),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_138),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_12),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_70),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_44),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_152),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_22),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_89),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_13),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_33),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_76),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_165),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_122),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_131),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_1),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_92),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_133),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_153),
.Y(n_239)
);

BUFx8_ASAP7_75t_SL g240 ( 
.A(n_91),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_36),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_8),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_197),
.Y(n_244)
);

BUFx2_ASAP7_75t_SL g245 ( 
.A(n_187),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_0),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_181),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_1),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_181),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_194),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_237),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_203),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_198),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_203),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_216),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g266 ( 
.A(n_188),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_237),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_207),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_207),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_L g270 ( 
.A(n_217),
.B(n_2),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_240),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_187),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_187),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_188),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_189),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_189),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_210),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_210),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_192),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_211),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_190),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_231),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_193),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_199),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_235),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_201),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_242),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_214),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_215),
.Y(n_293)
);

NAND2x1_ASAP7_75t_L g294 ( 
.A(n_257),
.B(n_218),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g298 ( 
.A(n_262),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_225),
.B(n_219),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_258),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_228),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_257),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_241),
.B(n_232),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_248),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_253),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_282),
.Y(n_307)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_257),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_272),
.B(n_202),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_258),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_251),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_271),
.Y(n_315)
);

CKINVDCx8_ASAP7_75t_R g316 ( 
.A(n_271),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_252),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_283),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_251),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_264),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_276),
.B(n_278),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_176),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_247),
.Y(n_326)
);

NAND2x1p5_ASAP7_75t_L g327 ( 
.A(n_270),
.B(n_177),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_281),
.B(n_179),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_272),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_245),
.B(n_180),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_257),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_277),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_284),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_256),
.B(n_182),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_274),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_290),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_254),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_255),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_277),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_285),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_285),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_249),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_332),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_273),
.Y(n_347)
);

BUFx10_ASAP7_75t_L g348 ( 
.A(n_329),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_311),
.Y(n_349)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_308),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_280),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_325),
.B(n_246),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_303),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_326),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_323),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_324),
.B(n_286),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_305),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_286),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_282),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx4_ASAP7_75t_SL g366 ( 
.A(n_331),
.Y(n_366)
);

NAND3xp33_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_250),
.C(n_291),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_324),
.B(n_261),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_327),
.B(n_183),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_324),
.B(n_263),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_307),
.Y(n_372)
);

BUFx8_ASAP7_75t_SL g373 ( 
.A(n_307),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_265),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_306),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_320),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_326),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_336),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

OAI22xp33_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_291),
.B1(n_269),
.B2(n_268),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_339),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_318),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_342),
.Y(n_388)
);

AO22x2_ASAP7_75t_L g389 ( 
.A1(n_301),
.A2(n_269),
.B1(n_268),
.B2(n_259),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_320),
.B(n_186),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_249),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_313),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_319),
.Y(n_394)
);

INVx4_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g396 ( 
.A(n_309),
.B(n_259),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_334),
.B(n_191),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_335),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_338),
.B(n_2),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_299),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_294),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_299),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_304),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_304),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_297),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_327),
.B(n_333),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_327),
.B(n_195),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_344),
.B(n_3),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_314),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_297),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_310),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_310),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_344),
.B(n_4),
.Y(n_413)
);

XOR2x2_ASAP7_75t_SL g414 ( 
.A(n_345),
.B(n_4),
.Y(n_414)
);

NAND2x1p5_ASAP7_75t_L g415 ( 
.A(n_314),
.B(n_321),
.Y(n_415)
);

OAI221xp5_ASAP7_75t_L g416 ( 
.A1(n_333),
.A2(n_341),
.B1(n_316),
.B2(n_205),
.C(n_206),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_353),
.A2(n_341),
.B(n_300),
.C(n_315),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_353),
.B(n_316),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_362),
.B(n_300),
.Y(n_419)
);

AOI22x1_ASAP7_75t_L g420 ( 
.A1(n_356),
.A2(n_315),
.B1(n_312),
.B2(n_321),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_406),
.B(n_312),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_358),
.Y(n_422)
);

O2A1O1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_354),
.A2(n_314),
.B(n_6),
.C(n_7),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_322),
.B1(n_318),
.B2(n_345),
.Y(n_424)
);

OR2x6_ASAP7_75t_L g425 ( 
.A(n_346),
.B(n_387),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_204),
.B(n_200),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_322),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_362),
.B(n_208),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_374),
.B(n_212),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_380),
.B(n_213),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_399),
.A2(n_230),
.B1(n_239),
.B2(n_238),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_351),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_399),
.A2(n_227),
.B1(n_236),
.B2(n_234),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_369),
.A2(n_233),
.B1(n_229),
.B2(n_224),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_394),
.B(n_220),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g440 ( 
.A(n_416),
.B(n_221),
.C(n_222),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_394),
.B(n_297),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_347),
.B(n_5),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_394),
.B(n_297),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_367),
.B(n_7),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_361),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_9),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_356),
.A2(n_83),
.B(n_170),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

BUFx8_ASAP7_75t_L g449 ( 
.A(n_391),
.Y(n_449)
);

AOI22xp33_ASAP7_75t_L g450 ( 
.A1(n_368),
.A2(n_370),
.B1(n_408),
.B2(n_413),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_392),
.B(n_9),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_10),
.Y(n_453)
);

OAI22xp33_ASAP7_75t_L g454 ( 
.A1(n_360),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_11),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_369),
.B(n_13),
.Y(n_456)
);

AND3x1_ASAP7_75t_L g457 ( 
.A(n_364),
.B(n_14),
.C(n_15),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_408),
.B(n_15),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_397),
.B(n_16),
.Y(n_459)
);

AND2x2_ASAP7_75t_SL g460 ( 
.A(n_408),
.B(n_16),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_368),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_350),
.Y(n_463)
);

NAND2x1_ASAP7_75t_L g464 ( 
.A(n_350),
.B(n_34),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_397),
.B(n_17),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_372),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_384),
.B(n_386),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_388),
.B(n_18),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_373),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_413),
.B(n_19),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_407),
.B(n_20),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_359),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_368),
.B(n_21),
.Y(n_474)
);

O2A1O1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_407),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_378),
.Y(n_477)
);

A2O1A1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_402),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_370),
.B(n_25),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_378),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_348),
.B(n_26),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_370),
.B(n_27),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_401),
.B(n_175),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_403),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_348),
.B(n_29),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g486 ( 
.A1(n_400),
.A2(n_98),
.B(n_167),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_356),
.B(n_30),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_383),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_383),
.Y(n_489)
);

NOR3xp33_ASAP7_75t_SL g490 ( 
.A(n_417),
.B(n_382),
.C(n_414),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_466),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_428),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_438),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_445),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

CKINVDCx8_ASAP7_75t_R g496 ( 
.A(n_425),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_418),
.B(n_348),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_418),
.B(n_375),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_425),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_442),
.B(n_375),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_448),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_442),
.B(n_375),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_L g504 ( 
.A1(n_460),
.A2(n_444),
.B1(n_472),
.B2(n_456),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_489),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_460),
.A2(n_396),
.B1(n_389),
.B2(n_381),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_448),
.Y(n_507)
);

NOR3xp33_ASAP7_75t_SL g508 ( 
.A(n_481),
.B(n_414),
.C(n_409),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_477),
.B(n_385),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_422),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_R g511 ( 
.A(n_449),
.B(n_385),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_462),
.B(n_404),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_431),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_385),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_435),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_462),
.Y(n_517)
);

AND3x2_ASAP7_75t_SL g518 ( 
.A(n_457),
.B(n_389),
.C(n_363),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_419),
.B(n_377),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_421),
.B(n_390),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_455),
.B(n_377),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_470),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_421),
.B(n_377),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_430),
.B(n_390),
.Y(n_525)
);

NOR2x1p5_ASAP7_75t_L g526 ( 
.A(n_439),
.B(n_389),
.Y(n_526)
);

INVx8_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

NOR3xp33_ASAP7_75t_SL g528 ( 
.A(n_485),
.B(n_31),
.C(n_415),
.Y(n_528)
);

NOR3xp33_ASAP7_75t_SL g529 ( 
.A(n_458),
.B(n_31),
.C(n_415),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_480),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_424),
.B(n_363),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_468),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_400),
.Y(n_533)
);

NOR3xp33_ASAP7_75t_SL g534 ( 
.A(n_471),
.B(n_366),
.C(n_405),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_422),
.B(n_404),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_451),
.B(n_411),
.Y(n_536)
);

INVx4_ASAP7_75t_L g537 ( 
.A(n_463),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_464),
.Y(n_538)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_424),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_451),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_473),
.B(n_411),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_473),
.Y(n_543)
);

AND3x1_ASAP7_75t_SL g544 ( 
.A(n_461),
.B(n_35),
.C(n_38),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_510),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g546 ( 
.A1(n_521),
.A2(n_487),
.B(n_426),
.Y(n_546)
);

OAI21x1_ASAP7_75t_L g547 ( 
.A1(n_535),
.A2(n_486),
.B(n_447),
.Y(n_547)
);

OAI21x1_ASAP7_75t_L g548 ( 
.A1(n_535),
.A2(n_483),
.B(n_427),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_492),
.Y(n_549)
);

OAI21xp33_ASAP7_75t_L g550 ( 
.A1(n_504),
.A2(n_465),
.B(n_459),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_533),
.A2(n_441),
.B(n_443),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_533),
.A2(n_446),
.B(n_469),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_499),
.B(n_456),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_536),
.A2(n_453),
.B(n_452),
.Y(n_554)
);

OAI21xp33_ASAP7_75t_L g555 ( 
.A1(n_490),
.A2(n_444),
.B(n_472),
.Y(n_555)
);

A2O1A1Ixp33_ASAP7_75t_L g556 ( 
.A1(n_524),
.A2(n_461),
.B(n_475),
.C(n_423),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g557 ( 
.A1(n_501),
.A2(n_412),
.B(n_433),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_536),
.A2(n_412),
.B(n_482),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_499),
.B(n_450),
.Y(n_559)
);

AOI221xp5_ASAP7_75t_SL g560 ( 
.A1(n_540),
.A2(n_454),
.B1(n_474),
.B2(n_479),
.C(n_436),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_542),
.A2(n_420),
.B(n_432),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_493),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_513),
.Y(n_563)
);

AO32x2_ASAP7_75t_L g564 ( 
.A1(n_518),
.A2(n_434),
.A3(n_395),
.B1(n_410),
.B2(n_405),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_494),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_513),
.Y(n_566)
);

OAI21xp5_ASAP7_75t_L g567 ( 
.A1(n_501),
.A2(n_440),
.B(n_437),
.Y(n_567)
);

AO31x2_ASAP7_75t_L g568 ( 
.A1(n_503),
.A2(n_484),
.A3(n_478),
.B(n_395),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_539),
.A2(n_450),
.B1(n_476),
.B2(n_410),
.Y(n_569)
);

NOR4xp25_ASAP7_75t_L g570 ( 
.A(n_531),
.B(n_366),
.C(n_405),
.D(n_395),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

AO31x2_ASAP7_75t_L g572 ( 
.A1(n_503),
.A2(n_410),
.A3(n_393),
.B(n_379),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_497),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_L g575 ( 
.A1(n_525),
.A2(n_366),
.B(n_393),
.C(n_371),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_527),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_520),
.Y(n_577)
);

NOR2xp67_ASAP7_75t_L g578 ( 
.A(n_491),
.B(n_498),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_542),
.A2(n_393),
.B(n_379),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_495),
.B(n_357),
.Y(n_580)
);

BUFx5_ASAP7_75t_L g581 ( 
.A(n_513),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_512),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_519),
.B(n_522),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_514),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_508),
.B(n_357),
.Y(n_585)
);

AO31x2_ASAP7_75t_L g586 ( 
.A1(n_543),
.A2(n_393),
.A3(n_379),
.B(n_371),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_527),
.Y(n_587)
);

OAI21x1_ASAP7_75t_L g588 ( 
.A1(n_509),
.A2(n_379),
.B(n_371),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_577),
.Y(n_589)
);

OAI22x1_ASAP7_75t_L g590 ( 
.A1(n_569),
.A2(n_526),
.B1(n_518),
.B2(n_500),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_571),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_582),
.Y(n_592)
);

BUFx12f_ASAP7_75t_L g593 ( 
.A(n_587),
.Y(n_593)
);

OR2x6_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_527),
.Y(n_594)
);

AO31x2_ASAP7_75t_L g595 ( 
.A1(n_556),
.A2(n_509),
.A3(n_515),
.B(n_516),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_556),
.A2(n_522),
.B(n_515),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_571),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_577),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_563),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_550),
.B(n_528),
.C(n_529),
.Y(n_600)
);

AO31x2_ASAP7_75t_L g601 ( 
.A1(n_545),
.A2(n_544),
.A3(n_537),
.B(n_513),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_563),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_548),
.A2(n_506),
.B(n_534),
.Y(n_603)
);

OAI21x1_ASAP7_75t_L g604 ( 
.A1(n_558),
.A2(n_507),
.B(n_502),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_563),
.B(n_541),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_545),
.Y(n_606)
);

OA21x2_ASAP7_75t_L g607 ( 
.A1(n_552),
.A2(n_517),
.B(n_513),
.Y(n_607)
);

NAND2x1p5_ASAP7_75t_L g608 ( 
.A(n_566),
.B(n_541),
.Y(n_608)
);

OAI21x1_ASAP7_75t_L g609 ( 
.A1(n_579),
.A2(n_502),
.B(n_507),
.Y(n_609)
);

AOI21xp33_ASAP7_75t_SL g610 ( 
.A1(n_555),
.A2(n_532),
.B(n_511),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_549),
.B(n_541),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_566),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_541),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g614 ( 
.A(n_559),
.B(n_523),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_559),
.A2(n_578),
.B1(n_583),
.B2(n_560),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_583),
.A2(n_537),
.B1(n_496),
.B2(n_538),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

CKINVDCx6p67_ASAP7_75t_R g618 ( 
.A(n_587),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_573),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_561),
.A2(n_538),
.B(n_371),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_567),
.A2(n_538),
.B1(n_365),
.B2(n_357),
.Y(n_621)
);

OAI221xp5_ASAP7_75t_L g622 ( 
.A1(n_546),
.A2(n_365),
.B1(n_40),
.B2(n_43),
.C(n_45),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_574),
.Y(n_623)
);

O2A1O1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_553),
.A2(n_365),
.B(n_46),
.C(n_49),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_575),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_588),
.A2(n_365),
.B(n_50),
.Y(n_626)
);

OAI21x1_ASAP7_75t_L g627 ( 
.A1(n_547),
.A2(n_39),
.B(n_51),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

BUFx4f_ASAP7_75t_SL g629 ( 
.A(n_584),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_566),
.Y(n_630)
);

AOI221xp5_ASAP7_75t_L g631 ( 
.A1(n_600),
.A2(n_553),
.B1(n_570),
.B2(n_585),
.C(n_580),
.Y(n_631)
);

AOI221xp5_ASAP7_75t_L g632 ( 
.A1(n_600),
.A2(n_580),
.B1(n_575),
.B2(n_568),
.C(n_564),
.Y(n_632)
);

OR2x2_ASAP7_75t_L g633 ( 
.A(n_619),
.B(n_572),
.Y(n_633)
);

AOI21xp33_ASAP7_75t_L g634 ( 
.A1(n_590),
.A2(n_554),
.B(n_551),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_605),
.B(n_576),
.Y(n_635)
);

AOI22x1_ASAP7_75t_L g636 ( 
.A1(n_596),
.A2(n_576),
.B1(n_568),
.B2(n_564),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_615),
.A2(n_557),
.B1(n_564),
.B2(n_568),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_619),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_L g639 ( 
.A1(n_590),
.A2(n_581),
.B1(n_564),
.B2(n_568),
.Y(n_639)
);

OAI211xp5_ASAP7_75t_SL g640 ( 
.A1(n_615),
.A2(n_572),
.B(n_586),
.C(n_581),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_605),
.B(n_586),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_614),
.A2(n_629),
.B1(n_622),
.B2(n_625),
.Y(n_642)
);

AOI22xp33_ASAP7_75t_L g643 ( 
.A1(n_614),
.A2(n_581),
.B1(n_572),
.B2(n_586),
.Y(n_643)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_623),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_616),
.A2(n_581),
.B1(n_572),
.B2(n_55),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_598),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_592),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_628),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_594),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_628),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_591),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_SL g652 ( 
.A1(n_603),
.A2(n_581),
.B1(n_54),
.B2(n_56),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_589),
.Y(n_653)
);

OR2x6_ASAP7_75t_L g654 ( 
.A(n_594),
.B(n_581),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_621),
.A2(n_53),
.B(n_57),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_611),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_656)
);

BUFx12f_ASAP7_75t_L g657 ( 
.A(n_589),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_SL g658 ( 
.A1(n_603),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_598),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_610),
.A2(n_67),
.B1(n_68),
.B2(n_71),
.Y(n_660)
);

AOI31xp33_ASAP7_75t_SL g661 ( 
.A1(n_610),
.A2(n_72),
.A3(n_73),
.B(n_74),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_591),
.B(n_75),
.Y(n_662)
);

AO221x2_ASAP7_75t_L g663 ( 
.A1(n_601),
.A2(n_595),
.B1(n_597),
.B2(n_627),
.C(n_606),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_597),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_606),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_611),
.B(n_169),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_593),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_613),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_613),
.B(n_77),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_594),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_670)
);

CKINVDCx11_ASAP7_75t_R g671 ( 
.A(n_593),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_624),
.A2(n_81),
.B(n_82),
.C(n_84),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_595),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_594),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_603),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_675)
);

NAND2x1p5_ASAP7_75t_L g676 ( 
.A(n_605),
.B(n_96),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_595),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_603),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_618),
.B(n_617),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_605),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_594),
.B(n_105),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_642),
.A2(n_599),
.B1(n_602),
.B2(n_617),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_661),
.A2(n_630),
.B(n_612),
.C(n_602),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_638),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_642),
.A2(n_660),
.B1(n_674),
.B2(n_656),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_679),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_660),
.A2(n_602),
.B1(n_617),
.B2(n_599),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_647),
.A2(n_630),
.B1(n_612),
.B2(n_599),
.Y(n_688)
);

OAI21xp5_ASAP7_75t_L g689 ( 
.A1(n_672),
.A2(n_627),
.B(n_604),
.Y(n_689)
);

BUFx12f_ASAP7_75t_L g690 ( 
.A(n_671),
.Y(n_690)
);

AOI221xp5_ASAP7_75t_L g691 ( 
.A1(n_637),
.A2(n_595),
.B1(n_601),
.B2(n_608),
.C(n_607),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_646),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_647),
.A2(n_618),
.B1(n_608),
.B2(n_607),
.Y(n_693)
);

OAI21x1_ASAP7_75t_SL g694 ( 
.A1(n_631),
.A2(n_607),
.B(n_601),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_668),
.A2(n_607),
.B1(n_608),
.B2(n_604),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_644),
.B(n_601),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_636),
.A2(n_626),
.B1(n_609),
.B2(n_620),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_655),
.A2(n_609),
.B1(n_626),
.B2(n_620),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_641),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_639),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_648),
.Y(n_701)
);

AO31x2_ASAP7_75t_L g702 ( 
.A1(n_637),
.A2(n_110),
.A3(n_112),
.B(n_113),
.Y(n_702)
);

OAI211xp5_ASAP7_75t_L g703 ( 
.A1(n_632),
.A2(n_114),
.B(n_118),
.C(n_120),
.Y(n_703)
);

AOI21xp33_ASAP7_75t_L g704 ( 
.A1(n_655),
.A2(n_125),
.B(n_127),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_675),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_705)
);

OAI211xp5_ASAP7_75t_SL g706 ( 
.A1(n_634),
.A2(n_134),
.B(n_135),
.C(n_136),
.Y(n_706)
);

AO21x2_ASAP7_75t_L g707 ( 
.A1(n_640),
.A2(n_137),
.B(n_140),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_650),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_633),
.B(n_651),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g710 ( 
.A1(n_645),
.A2(n_141),
.B(n_145),
.Y(n_710)
);

AOI222xp33_ASAP7_75t_L g711 ( 
.A1(n_681),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.C1(n_149),
.C2(n_150),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_678),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_641),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_664),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_681),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_L g716 ( 
.A1(n_658),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_635),
.B(n_162),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_657),
.Y(n_718)
);

AO21x1_ASAP7_75t_SL g719 ( 
.A1(n_673),
.A2(n_166),
.B(n_677),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_663),
.B(n_652),
.C(n_680),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_670),
.A2(n_649),
.B1(n_635),
.B2(n_669),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_686),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_701),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_708),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_714),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_709),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_696),
.B(n_663),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_684),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_686),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_691),
.B(n_643),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_707),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_685),
.A2(n_676),
.B1(n_654),
.B2(n_661),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_695),
.B(n_665),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_694),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_699),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_693),
.B(n_649),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_699),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_713),
.B(n_654),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_713),
.B(n_702),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_692),
.B(n_659),
.Y(n_740)
);

INVx4_ASAP7_75t_R g741 ( 
.A(n_717),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_702),
.B(n_654),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_702),
.B(n_666),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_707),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_689),
.Y(n_745)
);

BUFx2_ASAP7_75t_SL g746 ( 
.A(n_721),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_689),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_697),
.B(n_676),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_710),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_710),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_688),
.Y(n_751)
);

OAI21x1_ASAP7_75t_SL g752 ( 
.A1(n_731),
.A2(n_683),
.B(n_704),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_732),
.A2(n_720),
.B(n_711),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_740),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_SL g755 ( 
.A1(n_730),
.A2(n_720),
.B1(n_703),
.B2(n_716),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_727),
.B(n_719),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_730),
.A2(n_711),
.B1(n_716),
.B2(n_712),
.Y(n_757)
);

AOI33xp33_ASAP7_75t_L g758 ( 
.A1(n_727),
.A2(n_725),
.A3(n_730),
.B1(n_751),
.B2(n_726),
.B3(n_734),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_724),
.Y(n_759)
);

AO21x2_ASAP7_75t_L g760 ( 
.A1(n_744),
.A2(n_698),
.B(n_682),
.Y(n_760)
);

NOR4xp25_ASAP7_75t_SL g761 ( 
.A(n_745),
.B(n_653),
.C(n_667),
.D(n_706),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_SL g762 ( 
.A1(n_742),
.A2(n_705),
.B1(n_712),
.B2(n_690),
.Y(n_762)
);

AOI221xp5_ASAP7_75t_L g763 ( 
.A1(n_745),
.A2(n_705),
.B1(n_700),
.B2(n_687),
.C(n_715),
.Y(n_763)
);

AOI33xp33_ASAP7_75t_L g764 ( 
.A1(n_727),
.A2(n_662),
.A3(n_718),
.B1(n_725),
.B2(n_751),
.B3(n_726),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_722),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_747),
.B(n_718),
.Y(n_766)
);

NOR2x1_ASAP7_75t_SL g767 ( 
.A(n_746),
.B(n_739),
.Y(n_767)
);

OAI221xp5_ASAP7_75t_L g768 ( 
.A1(n_743),
.A2(n_747),
.B1(n_746),
.B2(n_749),
.C(n_750),
.Y(n_768)
);

OAI31xp33_ASAP7_75t_L g769 ( 
.A1(n_743),
.A2(n_748),
.A3(n_742),
.B(n_739),
.Y(n_769)
);

AND2x4_ASAP7_75t_L g770 ( 
.A(n_735),
.B(n_722),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_742),
.A2(n_748),
.B1(n_750),
.B2(n_749),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_748),
.B(n_734),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_749),
.A2(n_750),
.B1(n_736),
.B2(n_733),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_756),
.B(n_772),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_756),
.B(n_735),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_759),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_772),
.B(n_735),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_759),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_772),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_772),
.B(n_734),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_758),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_770),
.B(n_731),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_769),
.B(n_724),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_770),
.B(n_767),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_767),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_764),
.B(n_733),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_770),
.B(n_737),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_766),
.B(n_737),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_786),
.B(n_769),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_778),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_774),
.B(n_754),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_778),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_781),
.B(n_765),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_781),
.B(n_783),
.Y(n_794)
);

NOR2x1p5_ASAP7_75t_L g795 ( 
.A(n_774),
.B(n_722),
.Y(n_795)
);

AOI31xp33_ASAP7_75t_L g796 ( 
.A1(n_794),
.A2(n_753),
.A3(n_755),
.B(n_762),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_793),
.Y(n_797)
);

NAND4xp75_ASAP7_75t_L g798 ( 
.A(n_791),
.B(n_763),
.C(n_784),
.D(n_779),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_790),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_789),
.A2(n_757),
.B(n_752),
.Y(n_800)
);

OAI22xp33_ASAP7_75t_L g801 ( 
.A1(n_796),
.A2(n_783),
.B1(n_768),
.B2(n_731),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_800),
.B(n_792),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_797),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_798),
.A2(n_771),
.B1(n_760),
.B2(n_773),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_803),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_802),
.B(n_796),
.Y(n_806)
);

NAND3xp33_ASAP7_75t_L g807 ( 
.A(n_806),
.B(n_804),
.C(n_801),
.Y(n_807)
);

BUFx2_ASAP7_75t_L g808 ( 
.A(n_805),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_805),
.Y(n_809)
);

NOR4xp25_ASAP7_75t_L g810 ( 
.A(n_807),
.B(n_799),
.C(n_785),
.D(n_788),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_808),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_809),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_808),
.B(n_785),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_807),
.B(n_731),
.C(n_761),
.Y(n_814)
);

INVxp33_ASAP7_75t_L g815 ( 
.A(n_811),
.Y(n_815)
);

INVxp33_ASAP7_75t_SL g816 ( 
.A(n_812),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_SL g817 ( 
.A1(n_814),
.A2(n_813),
.B(n_810),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_811),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_811),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_819),
.Y(n_820)
);

NOR3xp33_ASAP7_75t_L g821 ( 
.A(n_817),
.B(n_818),
.C(n_816),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_SL g822 ( 
.A1(n_815),
.A2(n_784),
.B(n_782),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_818),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_817),
.A2(n_752),
.B(n_761),
.Y(n_824)
);

NAND4xp25_ASAP7_75t_L g825 ( 
.A(n_821),
.B(n_775),
.C(n_788),
.D(n_729),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_823),
.A2(n_795),
.B1(n_782),
.B2(n_775),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_820),
.B(n_824),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_822),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_823),
.B(n_777),
.Y(n_829)
);

NAND5xp2_ASAP7_75t_L g830 ( 
.A(n_821),
.B(n_782),
.C(n_777),
.D(n_741),
.E(n_787),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_823),
.B(n_787),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_829),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_831),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_828),
.B(n_722),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_827),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_825),
.Y(n_836)
);

OR3x1_ASAP7_75t_L g837 ( 
.A(n_830),
.B(n_741),
.C(n_729),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_832),
.Y(n_838)
);

CKINVDCx16_ASAP7_75t_R g839 ( 
.A(n_833),
.Y(n_839)
);

NAND4xp25_ASAP7_75t_L g840 ( 
.A(n_835),
.B(n_826),
.C(n_729),
.D(n_780),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_836),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_SL g842 ( 
.A(n_836),
.B(n_736),
.C(n_776),
.Y(n_842)
);

OAI222xp33_ASAP7_75t_L g843 ( 
.A1(n_834),
.A2(n_779),
.B1(n_780),
.B2(n_744),
.C1(n_724),
.C2(n_733),
.Y(n_843)
);

AO21x1_ASAP7_75t_L g844 ( 
.A1(n_838),
.A2(n_839),
.B(n_841),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_844),
.A2(n_837),
.B1(n_842),
.B2(n_840),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_845),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_846),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_SL g848 ( 
.A1(n_847),
.A2(n_843),
.B1(n_744),
.B2(n_780),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_848),
.Y(n_849)
);

AOI221xp5_ASAP7_75t_L g850 ( 
.A1(n_849),
.A2(n_760),
.B1(n_728),
.B2(n_729),
.C(n_723),
.Y(n_850)
);

AOI211xp5_ASAP7_75t_L g851 ( 
.A1(n_850),
.A2(n_738),
.B(n_728),
.C(n_723),
.Y(n_851)
);


endmodule