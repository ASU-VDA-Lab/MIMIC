module fake_jpeg_21310_n_202 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx4f_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx4f_ASAP7_75t_SL g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_35),
.Y(n_41)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_21),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_18),
.B1(n_23),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_50),
.B1(n_23),
.B2(n_16),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_19),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_30),
.B(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_55),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_18),
.B1(n_32),
.B2(n_34),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_56),
.B(n_60),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_34),
.C(n_39),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_66),
.C(n_74),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_77),
.B1(n_75),
.B2(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_16),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_21),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_64),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_27),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_35),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_67),
.Y(n_97)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_45),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_72),
.A2(n_76),
.B1(n_57),
.B2(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_28),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_31),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_39),
.B1(n_30),
.B2(n_46),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_31),
.B1(n_39),
.B2(n_30),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_22),
.Y(n_78)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_39),
.B1(n_30),
.B2(n_38),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_92),
.B1(n_56),
.B2(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_77),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_46),
.B(n_26),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_94),
.B(n_100),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_46),
.B(n_26),
.C(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_59),
.B1(n_24),
.B2(n_3),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_60),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_102),
.A2(n_103),
.B1(n_106),
.B2(n_107),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_81),
.A2(n_68),
.B1(n_71),
.B2(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_115),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_67),
.B1(n_73),
.B2(n_52),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_119),
.B1(n_1),
.B2(n_2),
.Y(n_142)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_26),
.B(n_53),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_92),
.B(n_89),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_88),
.B(n_13),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_109),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_101),
.B(n_12),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_12),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_26),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_118),
.C(n_79),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_20),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_26),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_113),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_94),
.B(n_87),
.C(n_79),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_123),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_124),
.A2(n_86),
.B1(n_90),
.B2(n_59),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_122),
.A2(n_97),
.B1(n_100),
.B2(n_87),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_100),
.B(n_91),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_132),
.B(n_143),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_123),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_102),
.A2(n_82),
.B1(n_98),
.B2(n_85),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_106),
.A2(n_92),
.B1(n_84),
.B2(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_124),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_130),
.B1(n_129),
.B2(n_112),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_118),
.A2(n_24),
.B(n_4),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_156),
.B(n_158),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_107),
.B1(n_117),
.B2(n_104),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_105),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_121),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_158),
.B1(n_145),
.B2(n_148),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_110),
.C(n_4),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_143),
.C(n_140),
.Y(n_163)
);

OAI322xp33_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_1),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_8),
.C2(n_10),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_136),
.Y(n_158)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_126),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_163),
.B(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_144),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_135),
.B1(n_138),
.B2(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

AOI321xp33_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_132),
.A3(n_141),
.B1(n_138),
.B2(n_127),
.C(n_6),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_161),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_165),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_155),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_177),
.C(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_152),
.C(n_154),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_141),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_168),
.Y(n_184)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_166),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_7),
.B(n_8),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_183),
.Y(n_190)
);

OAI31xp33_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_169),
.A3(n_162),
.B(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_168),
.C(n_157),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_7),
.C(n_8),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_185),
.B(n_10),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_175),
.B1(n_172),
.B2(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_189),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_11),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_188),
.A2(n_181),
.B1(n_171),
.B2(n_11),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_192),
.B(n_193),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_171),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_195),
.A2(n_181),
.B1(n_190),
.B2(n_11),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_196),
.A2(n_194),
.B(n_192),
.Y(n_198)
);

INVxp33_ASAP7_75t_SL g200 ( 
.A(n_198),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_193),
.C(n_196),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_200),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule