module fake_jpeg_18754_n_274 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_14;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_7),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_13),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_33),
.Y(n_42)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_26),
.Y(n_49)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_50),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_26),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_51),
.A2(n_55),
.B1(n_40),
.B2(n_38),
.Y(n_67)
);

OR2x4_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_23),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_43),
.Y(n_66)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_13),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_60),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_28),
.B1(n_27),
.B2(n_18),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_41),
.C(n_35),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_63),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_78),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_70),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_60),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_16),
.B1(n_13),
.B2(n_18),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_57),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_56),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_79),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_33),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_94),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_64),
.B(n_65),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_72),
.Y(n_103)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_25),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_97),
.Y(n_104)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_25),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_85),
.B1(n_70),
.B2(n_95),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_101),
.B1(n_114),
.B2(n_91),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_77),
.B1(n_62),
.B2(n_54),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_77),
.B(n_72),
.C(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_103),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_68),
.B1(n_71),
.B2(n_35),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_33),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_109),
.C(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_88),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_112),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_41),
.C(n_46),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_33),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_74),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_84),
.A2(n_86),
.B1(n_97),
.B2(n_92),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_118),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_80),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_18),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_80),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_91),
.B(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_127),
.B(n_22),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g122 ( 
.A(n_113),
.B(n_89),
.C(n_94),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_129),
.B1(n_40),
.B2(n_29),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_109),
.A2(n_91),
.B1(n_15),
.B2(n_11),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_61),
.B1(n_74),
.B2(n_54),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_98),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_136),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_89),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_138),
.B(n_144),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_141),
.Y(n_162)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_142),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_104),
.Y(n_141)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_102),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_145),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_147),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_61),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_168),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_11),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_11),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_160),
.A2(n_170),
.B(n_127),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_11),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_163),
.B(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_141),
.B(n_12),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_58),
.C(n_47),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_129),
.C(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_12),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_15),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_147),
.B(n_124),
.C(n_120),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_187),
.C(n_188),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_145),
.B(n_121),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_134),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_160),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_121),
.B1(n_139),
.B2(n_132),
.Y(n_180)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_150),
.A2(n_128),
.B(n_130),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_45),
.C(n_47),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_58),
.C(n_45),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_142),
.C(n_140),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_192),
.Y(n_203)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_40),
.B1(n_15),
.B2(n_14),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_194),
.A2(n_154),
.B1(n_151),
.B2(n_172),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_170),
.B1(n_171),
.B2(n_156),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_195),
.A2(n_174),
.B1(n_187),
.B2(n_178),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_196),
.B(n_208),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_206),
.A3(n_212),
.B1(n_178),
.B2(n_183),
.C1(n_34),
.C2(n_23),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_153),
.B(n_169),
.C(n_158),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_201),
.A2(n_211),
.B(n_7),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_193),
.A2(n_153),
.B1(n_149),
.B2(n_158),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_19),
.Y(n_208)
);

NOR2xp67_ASAP7_75t_SL g211 ( 
.A(n_189),
.B(n_5),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_185),
.B1(n_182),
.B2(n_175),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_184),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_217),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_198),
.B(n_183),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_221),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_209),
.A2(n_12),
.B(n_22),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_225),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_202),
.A2(n_14),
.B1(n_29),
.B2(n_20),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_29),
.B1(n_14),
.B2(n_20),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_9),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_14),
.B1(n_20),
.B2(n_23),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_200),
.B(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_210),
.C(n_200),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_232),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_225),
.B(n_222),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_238),
.C(n_32),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_208),
.C(n_195),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_6),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_235),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_6),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_32),
.C(n_30),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_237),
.B(n_9),
.Y(n_240)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_240),
.Y(n_250)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_9),
.Y(n_241)
);

AOI31xp67_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_249),
.A3(n_8),
.B(n_16),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_245),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_8),
.Y(n_244)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_244),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_21),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_246),
.B(n_248),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_236),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_234),
.A2(n_236),
.B1(n_238),
.B2(n_16),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_243),
.A2(n_13),
.B(n_16),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_252),
.B(n_254),
.Y(n_259)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_239),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_8),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_257),
.B(n_258),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_21),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_249),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

A2O1A1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_19),
.B(n_1),
.C(n_2),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_263),
.B(n_264),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g264 ( 
.A1(n_256),
.A2(n_34),
.A3(n_30),
.B1(n_31),
.B2(n_19),
.C1(n_4),
.C2(n_3),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_258),
.B(n_251),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_266),
.A2(n_262),
.B(n_34),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_269),
.B(n_267),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_265),
.A2(n_262),
.B(n_31),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_19),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_271),
.A2(n_34),
.B(n_1),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_272),
.A2(n_0),
.B(n_1),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_3),
.B(n_4),
.Y(n_274)
);


endmodule