module fake_ariane_3103_n_460 (n_8, n_56, n_60, n_64, n_38, n_47, n_18, n_75, n_67, n_34, n_69, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_49, n_20, n_17, n_50, n_62, n_51, n_76, n_79, n_26, n_3, n_46, n_0, n_36, n_72, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_6, n_48, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_23, n_61, n_22, n_43, n_1, n_81, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_14, n_68, n_78, n_39, n_59, n_63, n_16, n_5, n_35, n_54, n_25, n_460);

input n_8;
input n_56;
input n_60;
input n_64;
input n_38;
input n_47;
input n_18;
input n_75;
input n_67;
input n_34;
input n_69;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_49;
input n_20;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_36;
input n_72;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_6;
input n_48;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_61;
input n_22;
input n_43;
input n_1;
input n_81;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_14;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_460;

wire n_295;
wire n_356;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_373;
wire n_299;
wire n_133;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_319;
wire n_416;
wire n_283;
wire n_187;
wire n_367;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_424;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_85;
wire n_130;
wire n_349;
wire n_391;
wire n_346;
wire n_214;
wire n_348;
wire n_410;
wire n_379;
wire n_445;
wire n_162;
wire n_138;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_441;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_87;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_167;
wire n_90;
wire n_422;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_95;
wire n_446;
wire n_143;
wire n_152;
wire n_405;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_115;
wire n_331;
wire n_401;
wire n_267;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_200;
wire n_166;
wire n_253;
wire n_218;
wire n_271;
wire n_247;
wire n_91;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_420;
wire n_439;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_301;
wire n_248;
wire n_277;
wire n_432;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_427;
wire n_108;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_88;
wire n_141;
wire n_390;
wire n_104;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_459;
wire n_221;
wire n_321;
wire n_86;
wire n_361;
wire n_458;
wire n_89;
wire n_149;
wire n_383;
wire n_237;
wire n_175;
wire n_453;
wire n_181;
wire n_260;
wire n_362;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_84;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_452;
wire n_178;
wire n_308;
wire n_417;
wire n_201;
wire n_343;
wire n_414;
wire n_287;
wire n_302;
wire n_380;
wire n_94;
wire n_284;
wire n_448;
wire n_249;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_278;
wire n_255;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_135;
wire n_409;
wire n_171;
wire n_384;
wire n_102;
wire n_182;
wire n_316;
wire n_196;
wire n_125;
wire n_407;
wire n_254;
wire n_219;
wire n_231;
wire n_366;
wire n_234;
wire n_280;
wire n_252;
wire n_215;
wire n_161;
wire n_454;
wire n_298;
wire n_415;
wire n_99;
wire n_216;
wire n_418;
wire n_223;
wire n_403;
wire n_83;
wire n_389;
wire n_288;
wire n_179;
wire n_395;
wire n_195;
wire n_213;
wire n_110;
wire n_304;
wire n_306;
wire n_313;
wire n_92;
wire n_430;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_268;
wire n_266;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_121;
wire n_118;
wire n_411;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_211;
wire n_97;
wire n_408;
wire n_322;
wire n_251;
wire n_116;
wire n_397;
wire n_351;
wire n_393;
wire n_359;
wire n_155;
wire n_127;

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_9),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_17),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g92 ( 
.A(n_61),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_11),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_9),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_26),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_60),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_32),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_36),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_29),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_1),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_45),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_5),
.Y(n_119)
);

INVxp33_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_12),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_54),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_6),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_15),
.Y(n_126)
);

NOR2xp67_ASAP7_75t_L g127 ( 
.A(n_14),
.B(n_31),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_12),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_19),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_27),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_66),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_40),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_39),
.Y(n_135)
);

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_69),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_33),
.Y(n_138)
);

NOR2xp67_ASAP7_75t_L g139 ( 
.A(n_8),
.B(n_62),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_4),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_73),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_41),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_18),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_46),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_16),
.B(n_34),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_10),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_44),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_8),
.Y(n_152)
);

NOR2xp67_ASAP7_75t_L g153 ( 
.A(n_43),
.B(n_56),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_25),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_3),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_64),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_75),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_51),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_0),
.Y(n_161)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_109),
.B(n_0),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_90),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_4),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_6),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_83),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_117),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_85),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

OAI21x1_ASAP7_75t_L g184 ( 
.A1(n_88),
.A2(n_22),
.B(n_23),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_98),
.B(n_24),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_102),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_101),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_146),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_91),
.B(n_30),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

OAI21x1_ASAP7_75t_L g200 ( 
.A1(n_94),
.A2(n_38),
.B(n_48),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_120),
.B(n_57),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_137),
.B(n_93),
.Y(n_202)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_103),
.A2(n_63),
.B(n_71),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g204 ( 
.A(n_93),
.B(n_84),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_97),
.B(n_76),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_81),
.B1(n_118),
.B2(n_108),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_143),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

AOI22x1_ASAP7_75t_SL g216 ( 
.A1(n_87),
.A2(n_128),
.B1(n_152),
.B2(n_130),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_113),
.A2(n_120),
.B1(n_107),
.B2(n_122),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_148),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_131),
.Y(n_219)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_149),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_149),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_99),
.A2(n_124),
.B1(n_113),
.B2(n_127),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_149),
.B(n_154),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_134),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g227 ( 
.A(n_96),
.B(n_116),
.Y(n_227)
);

OR2x6_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_147),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_227),
.B(n_116),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_163),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_96),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_168),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_157),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g234 ( 
.A(n_186),
.B(n_106),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_151),
.Y(n_235)
);

OR2x6_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_139),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_162),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_168),
.B(n_145),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_174),
.B(n_144),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_201),
.B(n_138),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_163),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_177),
.Y(n_242)
);

AO21x2_ASAP7_75t_L g243 ( 
.A1(n_198),
.A2(n_141),
.B(n_153),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_178),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

OR2x6_ASAP7_75t_L g246 ( 
.A(n_190),
.B(n_100),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_221),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_205),
.A2(n_154),
.B1(n_92),
.B2(n_95),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_187),
.B(n_89),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_177),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_187),
.B(n_105),
.Y(n_252)
);

AND3x2_ASAP7_75t_L g253 ( 
.A(n_208),
.B(n_167),
.C(n_210),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_111),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_165),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_166),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_178),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

INVxp33_ASAP7_75t_SL g260 ( 
.A(n_207),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_166),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_205),
.A2(n_123),
.B1(n_133),
.B2(n_136),
.Y(n_262)
);

AND2x6_ASAP7_75t_L g263 ( 
.A(n_205),
.B(n_142),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_181),
.B(n_156),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g265 ( 
.A1(n_205),
.A2(n_192),
.B1(n_222),
.B2(n_219),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_185),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_208),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_220),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_167),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_193),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_202),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_265),
.B(n_202),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_202),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_192),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_192),
.B1(n_164),
.B2(n_171),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_224),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_251),
.B(n_224),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_235),
.A2(n_172),
.B1(n_222),
.B2(n_219),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_206),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_186),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_229),
.A2(n_176),
.B1(n_207),
.B2(n_213),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_176),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_231),
.A2(n_203),
.B(n_200),
.C(n_184),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_226),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_234),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_258),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_209),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_239),
.B(n_218),
.Y(n_295)
);

AND2x6_ASAP7_75t_SL g296 ( 
.A(n_228),
.B(n_196),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_239),
.B(n_218),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_232),
.B(n_246),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_199),
.B1(n_193),
.B2(n_211),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_263),
.A2(n_216),
.B1(n_211),
.B2(n_214),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_240),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

BUFx3_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_254),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_254),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_240),
.A2(n_200),
.B(n_184),
.C(n_203),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_292),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_228),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_274),
.A2(n_260),
.B1(n_263),
.B2(n_243),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_273),
.B(n_243),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_283),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_276),
.A2(n_280),
.B(n_284),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_286),
.A2(n_297),
.B(n_295),
.C(n_275),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_244),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_282),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_195),
.B(n_194),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g321 ( 
.A1(n_278),
.A2(n_236),
.B(n_214),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_280),
.A2(n_188),
.B1(n_189),
.B2(n_170),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_253),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_288),
.A2(n_261),
.B(n_230),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_281),
.A2(n_261),
.B(n_241),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_281),
.A2(n_257),
.B(n_241),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_173),
.B1(n_170),
.B2(n_169),
.Y(n_329)
);

OAI22x1_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_216),
.B1(n_215),
.B2(n_212),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_173),
.B(n_179),
.C(n_180),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_289),
.B(n_215),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_307),
.B(n_294),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_279),
.B(n_215),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_298),
.B(n_212),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_301),
.A2(n_257),
.B(n_221),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_R g338 ( 
.A(n_285),
.B(n_212),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_279),
.B(n_266),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_304),
.A2(n_221),
.B(n_248),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_293),
.B(n_175),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_182),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_309),
.A2(n_182),
.B1(n_183),
.B2(n_191),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_309),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_274),
.A2(n_182),
.B1(n_183),
.B2(n_191),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_273),
.B(n_183),
.Y(n_348)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_284),
.A2(n_183),
.B1(n_191),
.B2(n_197),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

AO31x2_ASAP7_75t_L g351 ( 
.A1(n_320),
.A2(n_223),
.A3(n_332),
.B(n_339),
.Y(n_351)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_325),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_311),
.Y(n_353)
);

CKINVDCx6p67_ASAP7_75t_R g354 ( 
.A(n_331),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_324),
.A2(n_327),
.B(n_326),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_346),
.Y(n_358)
);

OAI21x1_ASAP7_75t_L g359 ( 
.A1(n_341),
.A2(n_345),
.B(n_337),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_323),
.Y(n_360)
);

O2A1O1Ixp33_ASAP7_75t_L g361 ( 
.A1(n_321),
.A2(n_333),
.B(n_336),
.C(n_322),
.Y(n_361)
);

INVx3_ASAP7_75t_SL g362 ( 
.A(n_342),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_338),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_330),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_313),
.B(n_349),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_344),
.A2(n_334),
.B(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx4_ASAP7_75t_L g369 ( 
.A(n_311),
.Y(n_369)
);

AO31x2_ASAP7_75t_L g370 ( 
.A1(n_320),
.A2(n_310),
.A3(n_287),
.B(n_314),
.Y(n_370)
);

AO31x2_ASAP7_75t_L g371 ( 
.A1(n_320),
.A2(n_310),
.A3(n_287),
.B(n_314),
.Y(n_371)
);

AO32x2_ASAP7_75t_L g372 ( 
.A1(n_322),
.A2(n_329),
.A3(n_299),
.B1(n_349),
.B2(n_316),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_316),
.A2(n_276),
.B1(n_273),
.B2(n_265),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_334),
.A2(n_317),
.B(n_348),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_334),
.A2(n_317),
.B(n_348),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_311),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_315),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_319),
.B(n_282),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_316),
.A2(n_276),
.B1(n_273),
.B2(n_265),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_316),
.A2(n_276),
.B(n_317),
.C(n_277),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_273),
.Y(n_382)
);

A2O1A1Ixp33_ASAP7_75t_L g383 ( 
.A1(n_316),
.A2(n_276),
.B(n_317),
.C(n_277),
.Y(n_383)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_312),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

NAND2x1p5_ASAP7_75t_L g386 ( 
.A(n_384),
.B(n_358),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_367),
.A2(n_382),
.B(n_383),
.Y(n_387)
);

A2O1A1Ixp33_ASAP7_75t_L g388 ( 
.A1(n_381),
.A2(n_373),
.B(n_380),
.C(n_361),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_378),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_350),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_368),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_365),
.B(n_384),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_365),
.B(n_384),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_359),
.B(n_366),
.Y(n_396)
);

NOR2x1_ASAP7_75t_R g397 ( 
.A(n_369),
.B(n_363),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_360),
.B(n_385),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_379),
.B(n_354),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_364),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_356),
.Y(n_401)
);

BUFx2_ASAP7_75t_R g402 ( 
.A(n_362),
.Y(n_402)
);

OR2x6_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_358),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_372),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_351),
.B(n_370),
.Y(n_406)
);

OA21x2_ASAP7_75t_L g407 ( 
.A1(n_370),
.A2(n_371),
.B(n_372),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_375),
.B(n_374),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_353),
.A2(n_318),
.B1(n_316),
.B2(n_260),
.Y(n_409)
);

INVx2_ASAP7_75t_SL g410 ( 
.A(n_376),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

AO21x2_ASAP7_75t_L g412 ( 
.A1(n_408),
.A2(n_387),
.B(n_388),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_411),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_409),
.B(n_390),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_393),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_401),
.Y(n_416)
);

INVx8_ASAP7_75t_L g417 ( 
.A(n_403),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_391),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_391),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_407),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_406),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_399),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_400),
.B(n_404),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_418),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_420),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_419),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_405),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_396),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_423),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_413),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_412),
.Y(n_432)
);

BUFx2_ASAP7_75t_SL g433 ( 
.A(n_424),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_429),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_426),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_429),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_434),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_435),
.B(n_427),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_436),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_433),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_432),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_438),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_443),
.Y(n_445)
);

NAND3xp33_ASAP7_75t_L g446 ( 
.A(n_443),
.B(n_441),
.C(n_437),
.Y(n_446)
);

AOI322xp5_ASAP7_75t_L g447 ( 
.A1(n_442),
.A2(n_414),
.A3(n_432),
.B1(n_431),
.B2(n_439),
.C1(n_425),
.C2(n_427),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_446),
.A2(n_441),
.B(n_444),
.Y(n_448)
);

AOI221xp5_ASAP7_75t_L g449 ( 
.A1(n_448),
.A2(n_445),
.B1(n_442),
.B2(n_422),
.C(n_447),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_449),
.Y(n_450)
);

NOR3xp33_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_389),
.C(n_410),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_389),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_403),
.C(n_415),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_452),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_454),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_455),
.A2(n_453),
.B1(n_433),
.B2(n_402),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_456),
.Y(n_457)
);

OA21x2_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_397),
.B(n_394),
.Y(n_458)
);

OR2x6_ASAP7_75t_L g459 ( 
.A(n_458),
.B(n_417),
.Y(n_459)
);

AOI21xp33_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_386),
.B(n_395),
.Y(n_460)
);


endmodule