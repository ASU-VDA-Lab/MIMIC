module real_jpeg_28019_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_150;
wire n_32;
wire n_20;
wire n_228;
wire n_80;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_0),
.A2(n_23),
.B1(n_24),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_0),
.A2(n_43),
.B1(n_47),
.B2(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_0),
.A2(n_49),
.B1(n_51),
.B2(n_66),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_1),
.B(n_51),
.Y(n_83)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_1),
.B(n_213),
.Y(n_218)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_1),
.Y(n_229)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_4),
.A2(n_6),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_30),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_4),
.A2(n_30),
.B1(n_43),
.B2(n_47),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_4),
.A2(n_30),
.B1(n_49),
.B2(n_51),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_5),
.A2(n_29),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_5),
.B(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_43),
.B1(n_47),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_5),
.A2(n_49),
.B1(n_51),
.B2(n_55),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_55),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_20),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_SL g179 ( 
.A1(n_5),
.A2(n_10),
.B(n_43),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_7),
.B(n_49),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_5),
.B(n_63),
.Y(n_208)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_6),
.A2(n_8),
.B1(n_29),
.B2(n_115),
.Y(n_114)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_8),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_115),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_8),
.A2(n_43),
.B1(n_47),
.B2(n_115),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_8),
.A2(n_49),
.B1(n_51),
.B2(n_115),
.Y(n_213)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_11),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_123),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_121),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_91),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_15),
.B(n_91),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_15),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_70),
.CI(n_78),
.CON(n_15),
.SN(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_37),
.B2(n_38),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_19),
.B(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_20),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_22),
.B(n_29),
.C(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_21),
.A2(n_33),
.B(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_23),
.B(n_26),
.Y(n_155)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_24),
.A2(n_58),
.B(n_59),
.C(n_63),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_24),
.B(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_24),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g178 ( 
.A1(n_24),
.A2(n_55),
.B(n_60),
.C(n_179),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_28),
.B(n_33),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_32),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_34),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_35),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_36),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_56),
.Y(n_38)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_39),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_39),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_52),
.B(n_53),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_41),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_41),
.B(n_54),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_41),
.B(n_186),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_47),
.B1(n_61),
.B2(n_62),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_43),
.A2(n_45),
.B(n_55),
.C(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_45),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_48),
.B(n_77),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_48),
.B(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_51),
.B(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_52),
.A2(n_76),
.B(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_52),
.B(n_55),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_55),
.B(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_64),
.B(n_67),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_57),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_57),
.B(n_142),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_57),
.Y(n_261)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_63),
.B(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_68),
.B(n_152),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_70),
.A2(n_71),
.B(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_72),
.B(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_72),
.A2(n_150),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_73),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_75),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_76),
.B(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_82),
.B(n_90),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_80),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_82),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_81),
.A2(n_82),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_81),
.A2(n_82),
.B1(n_87),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_82),
.B(n_178),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_86),
.Y(n_82)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_83),
.B(n_86),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_83),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_84),
.B(n_100),
.Y(n_132)
);

INVx11_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_87),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_89),
.B(n_195),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_116),
.C(n_117),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_92),
.A2(n_93),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_103),
.C(n_107),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_94),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_102),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_95),
.B(n_102),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_96),
.B(n_212),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_97),
.A2(n_131),
.B(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_98),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVxp33_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_103),
.A2(n_107),
.B1(n_108),
.B2(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_103),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_105),
.B(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_116),
.B(n_117),
.Y(n_282)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_278),
.B(n_283),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_265),
.B(n_277),
.Y(n_124)
);

O2A1O1Ixp33_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_172),
.B(n_247),
.C(n_264),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_160),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_127),
.B(n_160),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_143),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_129),
.B(n_135),
.C(n_143),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_130),
.B(n_133),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_132),
.B(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_134),
.B(n_185),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_138),
.C(n_139),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_137),
.B(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_145),
.B(n_148),
.C(n_153),
.Y(n_262)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_158),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_166),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_162),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.C(n_170),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_171),
.B(n_218),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_246),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_239),
.B(n_245),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_197),
.B(n_238),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_187),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_176),
.B(n_187),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_183),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_188),
.B(n_194),
.C(n_196),
.Y(n_240)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_233),
.B(n_237),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_214),
.B(n_232),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_205),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_203),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_211),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_210),
.C(n_211),
.Y(n_234)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_221),
.B(n_231),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_225),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_224),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_235),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_248),
.B(n_249),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_262),
.B2(n_263),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_253),
.C(n_263),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_257),
.C(n_259),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_266),
.B(n_267),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_276),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_274),
.C(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_279),
.B(n_280),
.Y(n_283)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);


endmodule