module real_aes_7299_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g276 ( .A(n_0), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g284 ( .A1(n_1), .A2(n_31), .B1(n_231), .B2(n_285), .Y(n_284) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_2), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_3), .B(n_256), .Y(n_265) );
INVx1_ASAP7_75t_L g212 ( .A(n_4), .Y(n_212) );
AND2x6_ASAP7_75t_L g249 ( .A(n_4), .B(n_210), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_4), .B(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_5), .A2(n_35), .B1(n_148), .B2(n_152), .Y(n_147) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_6), .A2(n_27), .B1(n_93), .B2(n_94), .Y(n_92) );
INVx1_ASAP7_75t_L g227 ( .A(n_7), .Y(n_227) );
INVx1_ASAP7_75t_L g269 ( .A(n_8), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_9), .B(n_235), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_10), .B(n_223), .Y(n_340) );
AO32x2_ASAP7_75t_L g282 ( .A1(n_11), .A2(n_222), .A3(n_248), .B1(n_256), .B2(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g308 ( .A(n_12), .B(n_231), .Y(n_308) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_13), .A2(n_29), .B1(n_93), .B2(n_97), .Y(n_96) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_14), .B(n_223), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_15), .A2(n_41), .B1(n_231), .B2(n_285), .Y(n_286) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_16), .A2(n_62), .B1(n_231), .B2(n_235), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_17), .B(n_231), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_18), .A2(n_50), .B1(n_169), .B2(n_171), .Y(n_168) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_19), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_20), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_21), .B(n_127), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_22), .A2(n_188), .B1(n_195), .B2(n_196), .Y(n_187) );
INVx1_ASAP7_75t_L g195 ( .A(n_22), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_23), .A2(n_81), .B1(n_82), .B2(n_536), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_23), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_24), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_25), .B(n_251), .Y(n_299) );
INVx2_ASAP7_75t_L g233 ( .A(n_26), .Y(n_233) );
OAI22xp5_ASAP7_75t_SL g197 ( .A1(n_28), .A2(n_43), .B1(n_198), .B2(n_199), .Y(n_197) );
INVx1_ASAP7_75t_L g199 ( .A(n_28), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_28), .B(n_231), .Y(n_230) );
OAI221xp5_ASAP7_75t_L g203 ( .A1(n_29), .A2(n_45), .B1(n_56), .B2(n_204), .C(n_205), .Y(n_203) );
INVxp67_ASAP7_75t_L g206 ( .A(n_29), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_30), .B(n_251), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_32), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g190 ( .A1(n_33), .A2(n_191), .B1(n_192), .B2(n_193), .Y(n_190) );
INVx1_ASAP7_75t_L g192 ( .A(n_33), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_34), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_36), .B(n_231), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_37), .A2(n_69), .B1(n_285), .B2(n_323), .Y(n_322) );
AOI22xp5_ASAP7_75t_SL g525 ( .A1(n_37), .A2(n_81), .B1(n_185), .B2(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_37), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_38), .B(n_231), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_39), .B(n_231), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_40), .B(n_243), .Y(n_263) );
AOI22xp33_ASAP7_75t_SL g338 ( .A1(n_42), .A2(n_46), .B1(n_231), .B2(n_235), .Y(n_338) );
INVx1_ASAP7_75t_L g198 ( .A(n_43), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_43), .B(n_231), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_44), .B(n_231), .Y(n_245) );
AO22x2_ASAP7_75t_L g102 ( .A1(n_45), .A2(n_65), .B1(n_93), .B2(n_97), .Y(n_102) );
INVxp67_ASAP7_75t_L g207 ( .A(n_45), .Y(n_207) );
INVx1_ASAP7_75t_L g210 ( .A(n_47), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_48), .B(n_231), .Y(n_277) );
INVx1_ASAP7_75t_L g226 ( .A(n_49), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_51), .Y(n_204) );
AO32x2_ASAP7_75t_L g320 ( .A1(n_52), .A2(n_248), .A3(n_256), .B1(n_321), .B2(n_325), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_53), .Y(n_86) );
INVx1_ASAP7_75t_L g241 ( .A(n_54), .Y(n_241) );
INVx1_ASAP7_75t_L g294 ( .A(n_55), .Y(n_294) );
AO22x2_ASAP7_75t_L g100 ( .A1(n_56), .A2(n_71), .B1(n_93), .B2(n_94), .Y(n_100) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_57), .A2(n_76), .B1(n_175), .B2(n_179), .Y(n_174) );
INVxp67_ASAP7_75t_L g191 ( .A(n_58), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_59), .B(n_235), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_60), .A2(n_81), .B1(n_184), .B2(n_185), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_60), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_61), .A2(n_67), .B1(n_157), .B2(n_162), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_63), .B(n_285), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_64), .B(n_235), .Y(n_298) );
INVx2_ASAP7_75t_L g224 ( .A(n_66), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_68), .B(n_235), .Y(n_260) );
INVx1_ASAP7_75t_L g534 ( .A(n_69), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_70), .A2(n_77), .B1(n_235), .B2(n_236), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_72), .A2(n_189), .B1(n_190), .B2(n_194), .Y(n_188) );
INVx1_ASAP7_75t_L g194 ( .A(n_72), .Y(n_194) );
INVx1_ASAP7_75t_L g93 ( .A(n_73), .Y(n_93) );
INVx1_ASAP7_75t_L g95 ( .A(n_73), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_74), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_75), .B(n_235), .Y(n_234) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_200), .B1(n_213), .B2(n_518), .C(n_524), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_186), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_81), .Y(n_185) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_145), .Y(n_83) );
NOR3xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_109), .C(n_131), .Y(n_84) );
OAI22xp5_ASAP7_75t_L g85 ( .A1(n_86), .A2(n_87), .B1(n_103), .B2(n_104), .Y(n_85) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
OR2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_98), .Y(n_89) );
INVx2_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
OR2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_96), .Y(n_90) );
AND2x2_ASAP7_75t_L g108 ( .A(n_91), .B(n_96), .Y(n_108) );
AND2x2_ASAP7_75t_L g151 ( .A(n_91), .B(n_123), .Y(n_151) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g114 ( .A(n_92), .B(n_96), .Y(n_114) );
AND2x2_ASAP7_75t_L g124 ( .A(n_92), .B(n_102), .Y(n_124) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx1_ASAP7_75t_L g97 ( .A(n_95), .Y(n_97) );
INVx2_ASAP7_75t_L g123 ( .A(n_96), .Y(n_123) );
INVx1_ASAP7_75t_L g165 ( .A(n_96), .Y(n_165) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
NAND2x1p5_ASAP7_75t_L g107 ( .A(n_99), .B(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g178 ( .A(n_99), .B(n_151), .Y(n_178) );
AND2x2_ASAP7_75t_L g99 ( .A(n_100), .B(n_101), .Y(n_99) );
INVx1_ASAP7_75t_L g116 ( .A(n_100), .Y(n_116) );
INVx1_ASAP7_75t_L g122 ( .A(n_100), .Y(n_122) );
INVx1_ASAP7_75t_L g144 ( .A(n_100), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_100), .B(n_102), .Y(n_166) );
AND2x2_ASAP7_75t_L g115 ( .A(n_101), .B(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g161 ( .A(n_102), .B(n_144), .Y(n_161) );
INVx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g160 ( .A(n_108), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g170 ( .A(n_108), .B(n_115), .Y(n_170) );
OAI221xp5_ASAP7_75t_SL g109 ( .A1(n_110), .A2(n_117), .B1(n_118), .B2(n_125), .C(n_126), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx4_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx4_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
INVx1_ASAP7_75t_L g141 ( .A(n_114), .Y(n_141) );
AND2x2_ASAP7_75t_L g150 ( .A(n_115), .B(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g154 ( .A(n_115), .B(n_155), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
INVx1_ASAP7_75t_L g130 ( .A(n_122), .Y(n_130) );
INVx1_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
AND2x4_ASAP7_75t_L g129 ( .A(n_124), .B(n_130), .Y(n_129) );
NAND2x1p5_ASAP7_75t_L g135 ( .A(n_124), .B(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B1(n_137), .B2(n_138), .Y(n_131) );
INVx3_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
CKINVDCx16_ASAP7_75t_R g139 ( .A(n_140), .Y(n_139) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_167), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_147), .B(n_156), .Y(n_146) );
BUFx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g173 ( .A(n_151), .B(n_161), .Y(n_173) );
AND2x4_ASAP7_75t_L g182 ( .A(n_151), .B(n_183), .Y(n_182) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx11_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx8_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx6_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
OR2x6_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_174), .Y(n_167) );
BUFx3_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
XNOR2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_197), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_188), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g193 ( .A(n_191), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
AND3x1_ASAP7_75t_SL g202 ( .A(n_203), .B(n_208), .C(n_211), .Y(n_202) );
INVxp67_ASAP7_75t_L g530 ( .A(n_203), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_208), .A2(n_520), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g540 ( .A(n_208), .Y(n_540) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OAI322xp33_ASAP7_75t_L g524 ( .A1(n_209), .A2(n_525), .A3(n_527), .B1(n_531), .B2(n_534), .C1(n_535), .C2(n_537), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_209), .B(n_212), .Y(n_533) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
OR2x2_ASAP7_75t_SL g539 ( .A(n_211), .B(n_540), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OR3x1_ASAP7_75t_L g215 ( .A(n_216), .B(n_446), .C(n_495), .Y(n_215) );
NAND5xp2_ASAP7_75t_L g216 ( .A(n_217), .B(n_361), .C(n_389), .D(n_419), .E(n_433), .Y(n_216) );
AOI221xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_279), .B1(n_311), .B2(n_316), .C(n_327), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_252), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_219), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g341 ( .A(n_220), .Y(n_341) );
AND2x2_ASAP7_75t_L g349 ( .A(n_220), .B(n_255), .Y(n_349) );
AND2x2_ASAP7_75t_L g372 ( .A(n_220), .B(n_254), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_220), .B(n_266), .Y(n_387) );
OR2x2_ASAP7_75t_L g396 ( .A(n_220), .B(n_334), .Y(n_396) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_220), .Y(n_399) );
AND2x2_ASAP7_75t_L g507 ( .A(n_220), .B(n_334), .Y(n_507) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_228), .B(n_250), .Y(n_220) );
OA21x2_ASAP7_75t_L g266 ( .A1(n_221), .A2(n_267), .B(n_278), .Y(n_266) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
AND2x2_ASAP7_75t_SL g251 ( .A(n_224), .B(n_225), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_240), .B(n_248), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_234), .B(n_237), .Y(n_229) );
INVx3_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
BUFx3_ASAP7_75t_L g323 ( .A(n_232), .Y(n_323) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g236 ( .A(n_233), .Y(n_236) );
INVx1_ASAP7_75t_L g244 ( .A(n_233), .Y(n_244) );
INVx2_ASAP7_75t_L g270 ( .A(n_235), .Y(n_270) );
INVx3_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
O2A1O1Ixp5_ASAP7_75t_SL g292 ( .A1(n_237), .A2(n_293), .B(n_294), .C(n_295), .Y(n_292) );
INVx5_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g321 ( .A1(n_238), .A2(n_247), .B1(n_322), .B2(n_324), .Y(n_321) );
INVx3_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_239), .Y(n_247) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_239), .Y(n_274) );
INVx1_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
O2A1O1Ixp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_245), .C(n_246), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_242), .A2(n_264), .B(n_276), .C(n_277), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_242), .B(n_521), .Y(n_520) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_246), .A2(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_247), .A2(n_264), .B1(n_284), .B2(n_286), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_247), .A2(n_264), .B1(n_337), .B2(n_338), .Y(n_336) );
NAND3xp33_ASAP7_75t_L g360 ( .A(n_248), .B(n_335), .C(n_336), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_248), .B(n_520), .Y(n_519) );
BUFx3_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_249), .A2(n_258), .B(n_261), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_268), .B(n_275), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g291 ( .A1(n_249), .A2(n_292), .B(n_296), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g301 ( .A1(n_249), .A2(n_302), .B(n_307), .Y(n_301) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_251), .A2(n_291), .B(n_299), .Y(n_290) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_251), .A2(n_301), .B(n_310), .Y(n_300) );
INVx2_ASAP7_75t_L g325 ( .A(n_251), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_252), .B(n_399), .Y(n_455) );
INVx2_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OAI311xp33_ASAP7_75t_L g397 ( .A1(n_253), .A2(n_398), .A3(n_399), .B1(n_400), .C1(n_415), .Y(n_397) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_266), .Y(n_253) );
AND2x2_ASAP7_75t_L g358 ( .A(n_254), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g365 ( .A(n_254), .Y(n_365) );
AND2x2_ASAP7_75t_L g486 ( .A(n_254), .B(n_315), .Y(n_486) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_255), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g342 ( .A(n_255), .B(n_266), .Y(n_342) );
AND2x2_ASAP7_75t_L g394 ( .A(n_255), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g408 ( .A(n_255), .B(n_341), .Y(n_408) );
OA21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_265), .Y(n_255) );
INVx4_ASAP7_75t_L g335 ( .A(n_256), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_264), .Y(n_261) );
INVx2_ASAP7_75t_L g315 ( .A(n_266), .Y(n_315) );
AND2x2_ASAP7_75t_L g357 ( .A(n_266), .B(n_341), .Y(n_357) );
O2A1O1Ixp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_270), .B(n_271), .C(n_272), .Y(n_268) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_273), .A2(n_297), .B(n_298), .Y(n_296) );
INVx4_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g523 ( .A(n_274), .Y(n_523) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_287), .Y(n_279) );
OR2x2_ASAP7_75t_L g452 ( .A(n_280), .B(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_280), .B(n_458), .Y(n_469) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_281), .B(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
AND2x2_ASAP7_75t_L g393 ( .A(n_282), .B(n_320), .Y(n_393) );
AND2x2_ASAP7_75t_L g404 ( .A(n_282), .B(n_300), .Y(n_404) );
AND2x2_ASAP7_75t_L g413 ( .A(n_282), .B(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_287), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_287), .B(n_354), .Y(n_398) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
OR2x2_ASAP7_75t_L g385 ( .A(n_288), .B(n_344), .Y(n_385) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_300), .Y(n_288) );
INVx2_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
AND2x2_ASAP7_75t_L g412 ( .A(n_289), .B(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
OR2x2_ASAP7_75t_L g429 ( .A(n_290), .B(n_430), .Y(n_429) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_290), .Y(n_492) );
AND2x2_ASAP7_75t_L g331 ( .A(n_300), .B(n_326), .Y(n_331) );
INVx1_ASAP7_75t_L g352 ( .A(n_300), .Y(n_352) );
AND2x2_ASAP7_75t_L g373 ( .A(n_300), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g414 ( .A(n_300), .Y(n_414) );
INVx1_ASAP7_75t_L g430 ( .A(n_300), .Y(n_430) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_300), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_313), .B(n_418), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_313), .A2(n_403), .B1(n_452), .B2(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
OAI211xp5_ASAP7_75t_SL g495 ( .A1(n_314), .A2(n_496), .B(n_498), .C(n_516), .Y(n_495) );
INVx2_ASAP7_75t_L g348 ( .A(n_315), .Y(n_348) );
AND2x2_ASAP7_75t_L g406 ( .A(n_315), .B(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g417 ( .A(n_315), .B(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_316), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x2_ASAP7_75t_L g390 ( .A(n_317), .B(n_354), .Y(n_390) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g422 ( .A(n_318), .B(n_413), .Y(n_422) );
AND2x2_ASAP7_75t_L g441 ( .A(n_318), .B(n_355), .Y(n_441) );
AND2x4_ASAP7_75t_L g377 ( .A(n_319), .B(n_351), .Y(n_377) );
AND2x2_ASAP7_75t_L g515 ( .A(n_319), .B(n_491), .Y(n_515) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_326), .Y(n_319) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_320), .Y(n_344) );
INVx1_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
INVx1_ASAP7_75t_L g454 ( .A(n_320), .Y(n_454) );
OR2x2_ASAP7_75t_L g345 ( .A(n_326), .B(n_330), .Y(n_345) );
AND2x2_ASAP7_75t_L g354 ( .A(n_326), .B(n_355), .Y(n_354) );
NOR2xp67_ASAP7_75t_L g374 ( .A(n_326), .B(n_375), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_332), .B1(n_343), .B2(n_346), .C(n_350), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_329), .A2(n_351), .B(n_353), .C(n_356), .Y(n_350) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_330), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_SL g458 ( .A(n_330), .B(n_352), .Y(n_458) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_330), .Y(n_465) );
AND2x2_ASAP7_75t_L g383 ( .A(n_331), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g420 ( .A(n_331), .B(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_342), .Y(n_332) );
INVx2_ASAP7_75t_L g411 ( .A(n_333), .Y(n_411) );
AOI222xp33_ASAP7_75t_L g460 ( .A1(n_333), .A2(n_344), .B1(n_461), .B2(n_463), .C1(n_464), .C2(n_466), .Y(n_460) );
AND2x2_ASAP7_75t_L g517 ( .A(n_333), .B(n_486), .Y(n_517) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_341), .Y(n_333) );
INVx1_ASAP7_75t_L g407 ( .A(n_334), .Y(n_407) );
AO21x1_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B(n_339), .Y(n_334) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g359 ( .A(n_340), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g445 ( .A(n_342), .B(n_379), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g456 ( .A1(n_343), .A2(n_457), .B(n_459), .Y(n_456) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx2_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_344), .B(n_351), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_344), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx3_ASAP7_75t_L g410 ( .A(n_348), .Y(n_410) );
OR2x2_ASAP7_75t_L g462 ( .A(n_348), .B(n_384), .Y(n_462) );
AND2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g416 ( .A(n_349), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_349), .B(n_410), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_349), .B(n_406), .Y(n_432) );
AND2x2_ASAP7_75t_L g436 ( .A(n_349), .B(n_418), .Y(n_436) );
INVxp67_ASAP7_75t_L g368 ( .A(n_351), .Y(n_368) );
BUFx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_353), .A2(n_426), .B1(n_431), .B2(n_432), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_353), .B(n_458), .Y(n_488) );
INVx1_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g474 ( .A(n_354), .B(n_465), .Y(n_474) );
AND2x2_ASAP7_75t_L g503 ( .A(n_354), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g508 ( .A(n_354), .B(n_458), .Y(n_508) );
INVx1_ASAP7_75t_L g421 ( .A(n_355), .Y(n_421) );
BUFx2_ASAP7_75t_L g427 ( .A(n_355), .Y(n_427) );
INVx1_ASAP7_75t_L g512 ( .A(n_356), .Y(n_512) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g363 ( .A(n_357), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g388 ( .A(n_358), .Y(n_388) );
NOR2x1_ASAP7_75t_L g364 ( .A(n_359), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g371 ( .A(n_359), .B(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g380 ( .A(n_359), .Y(n_380) );
INVx3_ASAP7_75t_L g418 ( .A(n_359), .Y(n_418) );
OR2x2_ASAP7_75t_L g484 ( .A(n_359), .B(n_485), .Y(n_484) );
AOI211xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_366), .B(n_369), .C(n_381), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_362), .A2(n_499), .B1(n_506), .B2(n_508), .C(n_509), .Y(n_498) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_370), .B(n_376), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_371), .B(n_373), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_372), .B(n_410), .Y(n_424) );
AND2x2_ASAP7_75t_L g466 ( .A(n_372), .B(n_406), .Y(n_466) );
INVx1_ASAP7_75t_SL g479 ( .A(n_373), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_373), .B(n_427), .Y(n_482) );
INVx1_ASAP7_75t_L g500 ( .A(n_374), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_378), .A2(n_468), .B1(n_470), .B2(n_474), .C(n_475), .Y(n_467) );
AND2x2_ASAP7_75t_L g494 ( .A(n_379), .B(n_486), .Y(n_494) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g478 ( .A(n_380), .Y(n_478) );
AOI21xp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_385), .B(n_386), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g449 ( .A(n_384), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g435 ( .A(n_385), .Y(n_435) );
INVx1_ASAP7_75t_L g463 ( .A(n_386), .Y(n_463) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
O2A1O1Ixp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_394), .C(n_397), .Y(n_389) );
OAI31xp33_ASAP7_75t_L g516 ( .A1(n_390), .A2(n_428), .A3(n_515), .B(n_517), .Y(n_516) );
INVxp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g490 ( .A(n_393), .B(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g511 ( .A(n_393), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_395), .B(n_410), .Y(n_438) );
INVx1_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g513 ( .A(n_396), .B(n_410), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_405), .B1(n_409), .B2(n_412), .Y(n_400) );
NAND2xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_403), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_404), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g440 ( .A(n_404), .B(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g443 ( .A(n_404), .B(n_427), .Y(n_443) );
AND2x2_ASAP7_75t_L g497 ( .A(n_404), .B(n_492), .Y(n_497) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx1_ASAP7_75t_L g472 ( .A(n_408), .Y(n_472) );
NOR2xp67_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
OAI32xp33_ASAP7_75t_L g475 ( .A1(n_410), .A2(n_444), .A3(n_476), .B1(n_478), .B2(n_479), .Y(n_475) );
INVx1_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_413), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g473 ( .A(n_417), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_423), .C(n_425), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_421), .B(n_458), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_422), .A2(n_434), .B1(n_435), .B2(n_436), .C(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_428), .Y(n_426) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g434 ( .A(n_432), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B1(n_442), .B2(n_444), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND4xp25_ASAP7_75t_SL g499 ( .A(n_442), .B(n_500), .C(n_501), .D(n_502), .Y(n_499) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
NAND4xp25_ASAP7_75t_SL g446 ( .A(n_447), .B(n_460), .C(n_467), .D(n_480), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_451), .B(n_455), .C(n_456), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_SL g477 ( .A(n_453), .Y(n_477) );
INVx2_ASAP7_75t_L g501 ( .A(n_458), .Y(n_501) );
OR2x2_ASAP7_75t_L g510 ( .A(n_465), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B(n_487), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g506 ( .A(n_486), .B(n_507), .Y(n_506) );
AOI21xp33_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_489), .B(n_493), .Y(n_487) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_509) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
CKINVDCx16_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_538), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
endmodule