module fake_jpeg_12437_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_40),
.Y(n_52)
);

CKINVDCx11_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_46),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_33),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_26),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_16),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_8),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_0),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_65),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_81),
.Y(n_89)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_1),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx6_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_56),
.A2(n_21),
.B(n_49),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_84),
.A2(n_61),
.B(n_71),
.C(n_57),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_74),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_91),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_3),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_72),
.B1(n_57),
.B2(n_67),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_97),
.B1(n_51),
.B2(n_53),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_64),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_69),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_75),
.A2(n_61),
.B1(n_55),
.B2(n_64),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_63),
.B(n_59),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_115),
.Y(n_119)
);

AO22x2_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_66),
.B1(n_62),
.B2(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_111),
.B1(n_113),
.B2(n_23),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_106),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_107),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_58),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_108),
.B(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_68),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_1),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_22),
.B1(n_48),
.B2(n_44),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_2),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_116),
.B(n_117),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_3),
.Y(n_117)
);

OAI211xp5_ASAP7_75t_L g118 ( 
.A1(n_98),
.A2(n_19),
.B(n_42),
.C(n_39),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_15),
.Y(n_127)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_120),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_102),
.B(n_106),
.C(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_5),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_6),
.Y(n_129)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_130),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_131),
.A2(n_133),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_50),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_134),
.B(n_9),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_7),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_10),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_127),
.B1(n_124),
.B2(n_126),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_25),
.C(n_37),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_140),
.B(n_141),
.C(n_144),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_13),
.C(n_31),
.Y(n_141)
);

AND2x6_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_119),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_142),
.B(n_146),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_27),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_29),
.B(n_38),
.C(n_11),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_145),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_125),
.B(n_131),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_121),
.B(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_146),
.C(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_156),
.B(n_152),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_149),
.B(n_153),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_158),
.A2(n_159),
.B(n_155),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_136),
.B1(n_143),
.B2(n_145),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_145),
.C(n_148),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_12),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_12),
.Y(n_164)
);


endmodule