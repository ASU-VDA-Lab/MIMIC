module fake_netlist_6_4442_n_2031 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_2031);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2031;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_683;
wire n_811;
wire n_474;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1650;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_2001;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_173),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_127),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_28),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_64),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_158),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_107),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_17),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_85),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_128),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_5),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_82),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_21),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_181),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_86),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_171),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_30),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_73),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_27),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_39),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_108),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_83),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_172),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_167),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_0),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_101),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_180),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_110),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_109),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_97),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_3),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_79),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_24),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_74),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_139),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_41),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_136),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_26),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

BUFx2_ASAP7_75t_SL g242 ( 
.A(n_81),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_119),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_73),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_45),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_135),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_124),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_61),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_138),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_36),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_142),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_41),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_9),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_57),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_17),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_129),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_43),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_178),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_161),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_112),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_165),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_100),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_102),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_104),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_47),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_37),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_48),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_76),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_164),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_56),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_90),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_123),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_168),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_114),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_34),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_137),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_13),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_77),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_71),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_186),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_34),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_53),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_152),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_48),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_130),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_36),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_117),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_159),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_4),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_20),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_13),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_113),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_126),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_59),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_68),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_143),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_103),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_170),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_51),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_27),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_10),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_118),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_105),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_29),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_7),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_21),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_174),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_94),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_23),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_68),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_166),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_51),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_49),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_69),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_6),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_67),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_1),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_52),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_35),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_151),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_16),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_59),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_6),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_71),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_50),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_0),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_80),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_15),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_92),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_106),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_19),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_38),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_93),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_78),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_31),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_3),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_185),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_179),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_95),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_39),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_62),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_133),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_145),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_20),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_1),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_125),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_54),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_89),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_19),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_99),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_91),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_148),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_60),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_188),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_24),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_156),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_25),
.Y(n_363)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_190),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_61),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_11),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_45),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_72),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_54),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_44),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_65),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_32),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_98),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_70),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_70),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_60),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_42),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_141),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_9),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_37),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_272),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_301),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_232),
.B(n_2),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_191),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_216),
.B(n_5),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_192),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_272),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_197),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_272),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_272),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_285),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_196),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_272),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_272),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_272),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_200),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_201),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_272),
.B(n_8),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_364),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_343),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_293),
.B(n_10),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_204),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_358),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_328),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_272),
.Y(n_406)
);

NOR2xp67_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_11),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_312),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_206),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_285),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_265),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_211),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_232),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_312),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_221),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_364),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_218),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_221),
.B(n_12),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_265),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_222),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_223),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_208),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_224),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_221),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_225),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_235),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_226),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_229),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_235),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_236),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_237),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_237),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_245),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_334),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_245),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_293),
.B(n_14),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_238),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_194),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_246),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_247),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_251),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_250),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_250),
.Y(n_445)
);

NOR2xp67_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_14),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_258),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_260),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_262),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_334),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_253),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_253),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_255),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_264),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_208),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_278),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_195),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_337),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_255),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_279),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_266),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_266),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_326),
.B(n_15),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_270),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_282),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_198),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_284),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_270),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_326),
.B(n_16),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_208),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_310),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_286),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_289),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_310),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_315),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_381),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_431),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_419),
.B(n_227),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_434),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_382),
.B(n_217),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_381),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_SL g485 ( 
.A(n_419),
.B(n_377),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_417),
.B(n_291),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_386),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_391),
.A2(n_287),
.B1(n_374),
.B2(n_305),
.Y(n_489)
);

NAND2xp33_ASAP7_75t_R g490 ( 
.A(n_440),
.B(n_385),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_382),
.B(n_217),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_393),
.B(n_199),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_416),
.B(n_227),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_387),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_416),
.B(n_227),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_393),
.B(n_199),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_388),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_389),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_425),
.B(n_340),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_389),
.Y(n_500)
);

INVx1_ASAP7_75t_SL g501 ( 
.A(n_411),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_390),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_390),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_393),
.B(n_400),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_434),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_400),
.B(n_294),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_402),
.B(n_243),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_394),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_437),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_399),
.B(n_377),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_400),
.B(n_298),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_394),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_438),
.B(n_299),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_405),
.A2(n_316),
.B1(n_327),
.B2(n_288),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_395),
.B(n_219),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_427),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_463),
.B(n_302),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_444),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_444),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_396),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_469),
.B(n_303),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_425),
.B(n_304),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_445),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_396),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_406),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_451),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_398),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_406),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_452),
.Y(n_534)
);

OAI21x1_ASAP7_75t_L g535 ( 
.A1(n_423),
.A2(n_357),
.B(n_219),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_423),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_423),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_408),
.B(n_340),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_455),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_455),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_470),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_470),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_408),
.B(n_340),
.Y(n_547)
);

BUFx8_ASAP7_75t_L g548 ( 
.A(n_383),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_414),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_453),
.B(n_314),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_414),
.B(n_193),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_410),
.B(n_249),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_453),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_450),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_538),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_477),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_477),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_481),
.A2(n_407),
.B1(n_446),
.B2(n_383),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_477),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_477),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_477),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_403),
.Y(n_562)
);

OAI22xp33_ASAP7_75t_L g563 ( 
.A1(n_490),
.A2(n_436),
.B1(n_405),
.B2(n_205),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_487),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_507),
.B(n_409),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_486),
.B(n_412),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_504),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_552),
.B(n_418),
.Y(n_568)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_489),
.B(n_436),
.C(n_254),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_498),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_481),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_552),
.A2(n_439),
.B1(n_447),
.B2(n_430),
.Y(n_573)
);

OR2x6_ASAP7_75t_L g574 ( 
.A(n_504),
.B(n_242),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_540),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_554),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_506),
.B(n_421),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_538),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_492),
.B(n_193),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_488),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_506),
.B(n_422),
.Y(n_582)
);

INVx4_ASAP7_75t_L g583 ( 
.A(n_540),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_486),
.B(n_424),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_515),
.B(n_426),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_498),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_512),
.B(n_429),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_540),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_515),
.B(n_432),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_497),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_540),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_492),
.B(n_496),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_532),
.B(n_441),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_520),
.B(n_442),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_484),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_498),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_492),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_548),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_511),
.B(n_446),
.C(n_407),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_484),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_512),
.B(n_443),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_498),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_520),
.B(n_456),
.Y(n_603)
);

AND2x2_ASAP7_75t_SL g604 ( 
.A(n_481),
.B(n_357),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_525),
.B(n_465),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_540),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_525),
.B(n_467),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_L g608 ( 
.A1(n_490),
.A2(n_311),
.B1(n_252),
.B2(n_281),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_508),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_493),
.B(n_415),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_484),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_548),
.B(n_472),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_485),
.A2(n_361),
.B1(n_315),
.B2(n_318),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_484),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_508),
.Y(n_616)
);

BUFx2_ASAP7_75t_L g617 ( 
.A(n_548),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_508),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_548),
.B(n_473),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_548),
.B(n_448),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_502),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_501),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_492),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_529),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_542),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_529),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_526),
.B(n_458),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_529),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_485),
.A2(n_274),
.B1(n_367),
.B2(n_292),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_483),
.B(n_449),
.Y(n_633)
);

OR2x6_ASAP7_75t_L g634 ( 
.A(n_483),
.B(n_242),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_526),
.B(n_457),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_492),
.Y(n_636)
);

NOR3xp33_ASAP7_75t_L g637 ( 
.A(n_489),
.B(n_466),
.C(n_428),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_550),
.B(n_275),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_529),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_491),
.A2(n_454),
.B1(n_460),
.B2(n_329),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_496),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_487),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_508),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_554),
.B(n_384),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_508),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_517),
.B(n_435),
.C(n_413),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_496),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_550),
.B(n_392),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_487),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_524),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_397),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_524),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_501),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_519),
.B(n_401),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_519),
.B(n_404),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_496),
.B(n_333),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_541),
.Y(n_658)
);

BUFx4f_ASAP7_75t_L g659 ( 
.A(n_487),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_517),
.A2(n_337),
.B1(n_233),
.B2(n_217),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_496),
.B(n_217),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_510),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_524),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_476),
.B(n_471),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_524),
.Y(n_665)
);

BUFx4f_ASAP7_75t_L g666 ( 
.A(n_487),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_541),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_542),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_524),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_487),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_493),
.B(n_202),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_511),
.B(n_207),
.C(n_202),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_541),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_518),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_510),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_542),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_518),
.B(n_233),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_518),
.A2(n_330),
.B1(n_318),
.B2(n_321),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_536),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_528),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_518),
.Y(n_682)
);

BUFx10_ASAP7_75t_L g683 ( 
.A(n_518),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_476),
.B(n_233),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_510),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_493),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_528),
.B(n_335),
.Y(n_688)
);

INVxp33_ASAP7_75t_SL g689 ( 
.A(n_495),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_R g690 ( 
.A(n_495),
.B(n_203),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_478),
.B(n_209),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_495),
.A2(n_499),
.B1(n_551),
.B2(n_547),
.Y(n_693)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_499),
.B(n_212),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_478),
.B(n_233),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_533),
.B(n_336),
.Y(n_696)
);

INVx4_ASAP7_75t_SL g697 ( 
.A(n_487),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_533),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_533),
.B(n_542),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_499),
.A2(n_321),
.B1(n_324),
.B2(n_330),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_551),
.B(n_415),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_536),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_551),
.B(n_207),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_533),
.B(n_345),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_479),
.B(n_349),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_487),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_542),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_576),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_562),
.B(n_213),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_604),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_565),
.B(n_215),
.C(n_214),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_604),
.B(n_494),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_597),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_597),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_689),
.A2(n_354),
.B1(n_356),
.B2(n_360),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_589),
.B(n_228),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_605),
.B(n_230),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_571),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_604),
.A2(n_533),
.B1(n_210),
.B2(n_373),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_578),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_588),
.B(n_275),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_567),
.B(n_494),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_566),
.B(n_231),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_578),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_636),
.Y(n_726)
);

A2O1A1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_572),
.A2(n_324),
.B(n_371),
.C(n_338),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_572),
.B(n_494),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_689),
.A2(n_378),
.B1(n_220),
.B2(n_234),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_588),
.B(n_494),
.Y(n_730)
);

AND2x4_ASAP7_75t_SL g731 ( 
.A(n_590),
.B(n_337),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_588),
.B(n_494),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_584),
.B(n_240),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_581),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_693),
.B(n_494),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_636),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_655),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_603),
.B(n_244),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_574),
.Y(n_739)
);

AOI22xp33_ASAP7_75t_L g740 ( 
.A1(n_687),
.A2(n_703),
.B1(n_634),
.B2(n_579),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_641),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_641),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_607),
.B(n_248),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_687),
.B(n_539),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_591),
.B(n_606),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_577),
.B(n_256),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_648),
.A2(n_378),
.B1(n_220),
.B2(n_234),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_591),
.B(n_494),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_592),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_558),
.A2(n_372),
.B(n_361),
.C(n_371),
.Y(n_751)
);

AND2x6_ASAP7_75t_SL g752 ( 
.A(n_656),
.B(n_338),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_664),
.B(n_479),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_592),
.Y(n_754)
);

INVx2_ASAP7_75t_SL g755 ( 
.A(n_592),
.Y(n_755)
);

BUFx6f_ASAP7_75t_SL g756 ( 
.A(n_590),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_591),
.B(n_494),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_674),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_703),
.A2(n_210),
.B1(n_352),
.B2(n_362),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_634),
.A2(n_239),
.B1(n_373),
.B2(n_241),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_674),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_598),
.B(n_239),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_606),
.B(n_500),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_635),
.A2(n_553),
.B(n_505),
.C(n_509),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_581),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_682),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_574),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_606),
.B(n_500),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_628),
.B(n_500),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_582),
.B(n_259),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_628),
.B(n_500),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_682),
.Y(n_772)
);

NOR2x1p5_ASAP7_75t_L g773 ( 
.A(n_630),
.B(n_263),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_628),
.B(n_500),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_694),
.B(n_480),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_694),
.B(n_480),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_707),
.B(n_500),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_611),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_595),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_634),
.A2(n_241),
.B1(n_362),
.B2(n_257),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_611),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_707),
.B(n_500),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_699),
.A2(n_535),
.B(n_503),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_707),
.B(n_500),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_587),
.B(n_269),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_647),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_647),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_575),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_575),
.B(n_503),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_595),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_601),
.B(n_271),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_600),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_L g794 ( 
.A1(n_703),
.A2(n_257),
.B1(n_352),
.B2(n_348),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_555),
.B(n_586),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_701),
.Y(n_796)
);

INVx8_ASAP7_75t_L g797 ( 
.A(n_574),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_574),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_634),
.A2(n_348),
.B1(n_267),
.B2(n_268),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_573),
.B(n_482),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_644),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_701),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_556),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_574),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_600),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_556),
.Y(n_806)
);

NOR2xp67_ASAP7_75t_L g807 ( 
.A(n_580),
.B(n_482),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_555),
.B(n_503),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_557),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_555),
.B(n_703),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_612),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_568),
.B(n_273),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_557),
.B(n_503),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_590),
.B(n_505),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_688),
.A2(n_535),
.B(n_514),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_559),
.B(n_503),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_634),
.A2(n_585),
.B1(n_594),
.B2(n_690),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_559),
.B(n_503),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_575),
.B(n_503),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_612),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_615),
.Y(n_821)
);

NAND2xp33_ASAP7_75t_L g822 ( 
.A(n_560),
.B(n_275),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_696),
.A2(n_535),
.B(n_514),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_560),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_691),
.B(n_509),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_583),
.B(n_503),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_583),
.B(n_514),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_561),
.B(n_514),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_561),
.B(n_275),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_570),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_626),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_570),
.B(n_514),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_SL g833 ( 
.A(n_563),
.B(n_283),
.C(n_276),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_583),
.B(n_514),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_596),
.B(n_514),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_668),
.B(n_514),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_615),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_671),
.Y(n_838)
);

AND2x2_ASAP7_75t_SL g839 ( 
.A(n_569),
.B(n_275),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_596),
.B(n_516),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_602),
.B(n_516),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_L g842 ( 
.A(n_602),
.B(n_275),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_609),
.B(n_516),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_626),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_609),
.B(n_516),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_618),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_593),
.B(n_290),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_610),
.B(n_516),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_640),
.B(n_295),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_610),
.B(n_516),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_671),
.B(n_579),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_608),
.B(n_296),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_616),
.Y(n_853)
);

NOR2x1p5_ASAP7_75t_L g854 ( 
.A(n_580),
.B(n_297),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_579),
.A2(n_280),
.B1(n_261),
.B2(n_267),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_616),
.B(n_516),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_618),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_619),
.B(n_516),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_620),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_668),
.B(n_545),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_619),
.B(n_539),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_643),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_705),
.B(n_300),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_625),
.B(n_513),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_668),
.B(n_545),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_643),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_579),
.B(n_513),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_645),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_684),
.B(n_306),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_672),
.A2(n_368),
.B(n_372),
.C(n_539),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_620),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_695),
.B(n_307),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_623),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_623),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_638),
.A2(n_553),
.B(n_521),
.C(n_544),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_625),
.B(n_521),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_671),
.B(n_522),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_645),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_650),
.B(n_547),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_671),
.Y(n_880)
);

BUFx3_ASAP7_75t_L g881 ( 
.A(n_713),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_716),
.A2(n_651),
.B(n_599),
.C(n_632),
.Y(n_882)
);

AOI21xp33_ASAP7_75t_L g883 ( 
.A1(n_724),
.A2(n_733),
.B(n_717),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_718),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_710),
.A2(n_599),
.B(n_632),
.C(n_672),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_814),
.B(n_654),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_825),
.B(n_671),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_709),
.B(n_650),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_744),
.B(n_654),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_722),
.A2(n_677),
.B(n_659),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_722),
.A2(n_677),
.B(n_659),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_803),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_710),
.B(n_677),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_738),
.B(n_653),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_746),
.A2(n_659),
.B(n_564),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_743),
.B(n_653),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_747),
.B(n_663),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_817),
.B(n_683),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_806),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_712),
.A2(n_704),
.B(n_665),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_744),
.B(n_637),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_740),
.A2(n_720),
.B1(n_735),
.B2(n_838),
.Y(n_902)
);

OAI21xp5_ASAP7_75t_L g903 ( 
.A1(n_712),
.A2(n_665),
.B(n_663),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_770),
.B(n_669),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_809),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_723),
.A2(n_666),
.B(n_564),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_786),
.B(n_669),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_792),
.B(n_675),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_753),
.B(n_675),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_839),
.A2(n_802),
.B1(n_796),
.B2(n_778),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_SL g911 ( 
.A(n_756),
.B(n_662),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_737),
.B(n_646),
.Y(n_912)
);

NOR2x1_ASAP7_75t_R g913 ( 
.A(n_877),
.B(n_662),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_757),
.A2(n_666),
.B(n_564),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_824),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_718),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_711),
.B(n_613),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_719),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_763),
.A2(n_666),
.B(n_657),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_782),
.B(n_681),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_830),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_838),
.A2(n_598),
.B1(n_617),
.B2(n_621),
.Y(n_922)
);

NOR2x1p5_ASAP7_75t_L g923 ( 
.A(n_775),
.B(n_676),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_853),
.Y(n_924)
);

INVx4_ASAP7_75t_L g925 ( 
.A(n_781),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_862),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_867),
.B(n_681),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_867),
.B(n_685),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_781),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_769),
.A2(n_777),
.B(n_771),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_877),
.B(n_617),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_751),
.A2(n_870),
.B(n_799),
.C(n_727),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_866),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_867),
.B(n_787),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_810),
.A2(n_692),
.B(n_685),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_864),
.B(n_633),
.Y(n_936)
);

NAND2x1_ASAP7_75t_L g937 ( 
.A(n_789),
.B(n_692),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_877),
.B(n_713),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_784),
.A2(n_698),
.B(n_627),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_781),
.B(n_683),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_868),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_876),
.B(n_676),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_878),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_788),
.B(n_698),
.Y(n_944)
);

O2A1O1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_751),
.A2(n_678),
.B(n_661),
.C(n_622),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_849),
.A2(n_660),
.B(n_614),
.C(n_700),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_781),
.B(n_683),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_766),
.B(n_624),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_831),
.B(n_642),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_783),
.A2(n_785),
.B(n_732),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_708),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_766),
.B(n_624),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_745),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_L g954 ( 
.A(n_831),
.B(n_642),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_852),
.A2(n_679),
.B(n_368),
.C(n_309),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_831),
.B(n_706),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_851),
.B(n_261),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_730),
.A2(n_649),
.B(n_642),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_772),
.B(n_627),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_839),
.A2(n_313),
.B1(n_277),
.B2(n_280),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_860),
.A2(n_631),
.B(n_629),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_754),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_730),
.A2(n_649),
.B(n_642),
.Y(n_963)
);

AND2x2_ASAP7_75t_SL g964 ( 
.A(n_760),
.B(n_268),
.Y(n_964)
);

AO21x1_ASAP7_75t_L g965 ( 
.A1(n_780),
.A2(n_317),
.B(n_308),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_851),
.B(n_277),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_880),
.B(n_308),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_772),
.Y(n_968)
);

AOI21xp33_ASAP7_75t_L g969 ( 
.A1(n_812),
.A2(n_686),
.B(n_313),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_732),
.A2(n_706),
.B(n_642),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_749),
.A2(n_774),
.B(n_768),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_795),
.B(n_629),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_807),
.B(n_686),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_749),
.A2(n_706),
.B(n_649),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_768),
.A2(n_706),
.B(n_649),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_831),
.B(n_706),
.Y(n_976)
);

OAI21x1_ASAP7_75t_L g977 ( 
.A1(n_815),
.A2(n_631),
.B(n_639),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_776),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_758),
.B(n_639),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_761),
.B(n_714),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_726),
.B(n_649),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_800),
.B(n_522),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_736),
.B(n_670),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_801),
.B(n_670),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_750),
.A2(n_670),
.B1(n_702),
.B2(n_680),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_741),
.B(n_670),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_774),
.A2(n_819),
.B(n_790),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_756),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_847),
.B(n_523),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_742),
.B(n_670),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_731),
.B(n_523),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_750),
.B(n_697),
.Y(n_992)
);

AOI21xp33_ASAP7_75t_L g993 ( 
.A1(n_863),
.A2(n_309),
.B(n_317),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_860),
.A2(n_865),
.B(n_819),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_728),
.B(n_680),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_755),
.B(n_702),
.Y(n_996)
);

BUFx2_ASAP7_75t_L g997 ( 
.A(n_762),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_880),
.B(n_339),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_731),
.B(n_527),
.Y(n_999)
);

AND2x6_ASAP7_75t_L g1000 ( 
.A(n_844),
.B(n_339),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_767),
.A2(n_344),
.B1(n_545),
.B2(n_530),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_755),
.B(n_652),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_764),
.B(n_652),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_779),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_715),
.B(n_319),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_869),
.B(n_320),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_872),
.B(n_322),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_789),
.B(n_658),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_790),
.A2(n_546),
.B(n_536),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_719),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_844),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_789),
.B(n_697),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_826),
.A2(n_834),
.B(n_827),
.Y(n_1013)
);

INVx3_ASAP7_75t_L g1014 ( 
.A(n_721),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_823),
.A2(n_673),
.B(n_667),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_826),
.A2(n_546),
.B(n_536),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_L g1017 ( 
.A1(n_865),
.A2(n_673),
.B(n_667),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_767),
.B(n_344),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_861),
.B(n_658),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_808),
.A2(n_547),
.B(n_545),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_827),
.A2(n_836),
.B(n_834),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_879),
.A2(n_836),
.B(n_816),
.Y(n_1022)
);

AOI21x1_ASAP7_75t_L g1023 ( 
.A1(n_813),
.A2(n_546),
.B(n_527),
.Y(n_1023)
);

OAI21xp33_ASAP7_75t_L g1024 ( 
.A1(n_748),
.A2(n_365),
.B(n_363),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_798),
.B(n_323),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_756),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_739),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_818),
.A2(n_832),
.B(n_828),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_721),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_798),
.B(n_697),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_835),
.A2(n_546),
.B(n_536),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_779),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_840),
.A2(n_545),
.B(n_537),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_759),
.B(n_697),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_804),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_804),
.B(n_325),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_794),
.B(n_530),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_725),
.B(n_531),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_729),
.B(n_531),
.Y(n_1039)
);

BUFx4f_ASAP7_75t_L g1040 ( 
.A(n_762),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_739),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_841),
.A2(n_543),
.B(n_537),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_791),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_791),
.Y(n_1044)
);

OAI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_843),
.A2(n_534),
.B(n_544),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_773),
.A2(n_534),
.B1(n_549),
.B2(n_370),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_845),
.A2(n_543),
.B(n_537),
.Y(n_1047)
);

BUFx3_ASAP7_75t_L g1048 ( 
.A(n_739),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_725),
.B(n_549),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_734),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_734),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_765),
.B(n_537),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_854),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_833),
.B(n_337),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_765),
.B(n_549),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_793),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_870),
.A2(n_475),
.B(n_474),
.C(n_468),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_762),
.B(n_331),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_848),
.A2(n_543),
.B(n_537),
.Y(n_1059)
);

OAI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_850),
.A2(n_459),
.B(n_461),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_855),
.B(n_549),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_762),
.B(n_459),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_856),
.A2(n_543),
.B(n_537),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_793),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_805),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_727),
.B(n_461),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_805),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_739),
.A2(n_549),
.B1(n_369),
.B2(n_366),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_811),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_811),
.Y(n_1070)
);

OAI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_858),
.A2(n_462),
.B(n_464),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_820),
.B(n_549),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_752),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_797),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_938),
.B(n_820),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_890),
.A2(n_891),
.B(n_954),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_951),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_925),
.Y(n_1078)
);

NAND2x1p5_ASAP7_75t_L g1079 ( 
.A(n_925),
.B(n_821),
.Y(n_1079)
);

BUFx8_ASAP7_75t_SL g1080 ( 
.A(n_988),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_SL g1081 ( 
.A1(n_883),
.A2(n_859),
.B(n_874),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_887),
.A2(n_797),
.B1(n_874),
.B2(n_873),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_882),
.A2(n_822),
.B(n_829),
.C(n_842),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_892),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_982),
.B(n_821),
.Y(n_1085)
);

AND2x4_ASAP7_75t_L g1086 ( 
.A(n_938),
.B(n_837),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_954),
.A2(n_797),
.B(n_822),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_882),
.A2(n_797),
.B(n_875),
.C(n_871),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_884),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_969),
.A2(n_829),
.B(n_842),
.C(n_859),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_978),
.B(n_837),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_906),
.A2(n_873),
.B(n_871),
.Y(n_1092)
);

BUFx3_ASAP7_75t_L g1093 ( 
.A(n_1053),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_901),
.B(n_846),
.Y(n_1094)
);

NAND2x1p5_ASAP7_75t_L g1095 ( 
.A(n_925),
.B(n_846),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1013),
.A2(n_857),
.B(n_462),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1021),
.A2(n_857),
.B(n_543),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1006),
.A2(n_1007),
.B(n_946),
.C(n_1005),
.Y(n_1098)
);

INVx1_ASAP7_75t_SL g1099 ( 
.A(n_889),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_886),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1006),
.B(n_332),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_898),
.A2(n_543),
.B(n_537),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_929),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1007),
.B(n_341),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_909),
.B(n_342),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_938),
.B(n_464),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_942),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_960),
.A2(n_468),
.B1(n_474),
.B2(n_475),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_884),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_988),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_987),
.A2(n_359),
.B(n_347),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_946),
.B(n_380),
.C(n_379),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_899),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_912),
.B(n_346),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_973),
.B(n_931),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1005),
.A2(n_355),
.B(n_351),
.C(n_353),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_898),
.A2(n_543),
.B(n_537),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_989),
.B(n_375),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_931),
.Y(n_1119)
);

INVx3_ASAP7_75t_L g1120 ( 
.A(n_929),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_930),
.A2(n_543),
.B(n_549),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_916),
.Y(n_1122)
);

AOI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_936),
.A2(n_350),
.B1(n_549),
.B2(n_183),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1058),
.B(n_18),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_893),
.A2(n_176),
.B(n_175),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_931),
.B(n_1011),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_984),
.B(n_18),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_893),
.A2(n_169),
.B(n_162),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_993),
.A2(n_157),
.B(n_155),
.C(n_153),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1008),
.A2(n_150),
.B(n_147),
.Y(n_1130)
);

O2A1O1Ixp5_ASAP7_75t_L g1131 ( 
.A1(n_888),
.A2(n_144),
.B(n_140),
.C(n_134),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_984),
.B(n_960),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1062),
.B(n_22),
.Y(n_1133)
);

NOR3xp33_ASAP7_75t_SL g1134 ( 
.A(n_1058),
.B(n_22),
.C(n_23),
.Y(n_1134)
);

NAND2x1p5_ASAP7_75t_L g1135 ( 
.A(n_1027),
.B(n_131),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_929),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_895),
.A2(n_122),
.B(n_120),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_917),
.A2(n_116),
.B1(n_115),
.B2(n_111),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_934),
.B(n_25),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_1011),
.B(n_96),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_R g1141 ( 
.A(n_1026),
.B(n_88),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_919),
.A2(n_87),
.B(n_84),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_929),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_914),
.A2(n_896),
.B(n_894),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_905),
.B(n_26),
.Y(n_1145)
);

BUFx2_ASAP7_75t_SL g1146 ( 
.A(n_1011),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_910),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_SL g1148 ( 
.A(n_945),
.B(n_32),
.C(n_33),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_916),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_910),
.A2(n_33),
.B1(n_38),
.B2(n_40),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_885),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1027),
.B(n_44),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_915),
.B(n_46),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_SL g1154 ( 
.A1(n_1073),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_885),
.A2(n_50),
.B(n_52),
.C(n_53),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1026),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_897),
.A2(n_76),
.B(n_58),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_955),
.A2(n_55),
.B(n_58),
.C(n_62),
.Y(n_1158)
);

O2A1O1Ixp33_ASAP7_75t_SL g1159 ( 
.A1(n_1030),
.A2(n_63),
.B(n_64),
.C(n_65),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_881),
.B(n_63),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_921),
.B(n_66),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_1074),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_902),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_922),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_904),
.A2(n_908),
.B(n_907),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_924),
.B(n_926),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1011),
.Y(n_1167)
);

INVx4_ASAP7_75t_L g1168 ( 
.A(n_1074),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1027),
.B(n_1074),
.Y(n_1169)
);

NOR2xp67_ASAP7_75t_L g1170 ( 
.A(n_1046),
.B(n_1068),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1040),
.B(n_991),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_950),
.A2(n_1022),
.B(n_1019),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_933),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_927),
.A2(n_928),
.B1(n_881),
.B2(n_941),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_999),
.A2(n_1036),
.B1(n_1025),
.B2(n_966),
.Y(n_1175)
);

OAI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_943),
.A2(n_1035),
.B1(n_1040),
.B2(n_1041),
.Y(n_1176)
);

INVx2_ASAP7_75t_SL g1177 ( 
.A(n_923),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_953),
.B(n_962),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1074),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_972),
.A2(n_976),
.B(n_956),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1041),
.B(n_1048),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1024),
.A2(n_1036),
.B(n_1025),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_920),
.B(n_957),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_955),
.A2(n_980),
.B(n_1054),
.C(n_1039),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1035),
.A2(n_1048),
.B1(n_971),
.B2(n_968),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_R g1186 ( 
.A(n_911),
.B(n_968),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_964),
.A2(n_1066),
.B1(n_965),
.B2(n_957),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_949),
.A2(n_976),
.B(n_956),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_957),
.B(n_966),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_940),
.B(n_947),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_949),
.A2(n_1028),
.B(n_935),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_966),
.B(n_997),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_961),
.A2(n_1017),
.B(n_1015),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_964),
.A2(n_1018),
.B1(n_967),
.B2(n_998),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_937),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_967),
.B(n_998),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_967),
.B(n_998),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_932),
.A2(n_1037),
.B(n_1018),
.C(n_903),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1018),
.B(n_918),
.Y(n_1199)
);

NAND2x1_ASAP7_75t_L g1200 ( 
.A(n_1056),
.B(n_1069),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1004),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_913),
.B(n_944),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_995),
.A2(n_1020),
.B(n_939),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1038),
.B(n_1051),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1014),
.B(n_1051),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1000),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1000),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1056),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_918),
.A2(n_1050),
.B1(n_1010),
.B2(n_1029),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1010),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1014),
.B(n_1069),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1029),
.A2(n_1050),
.B1(n_1070),
.B2(n_1032),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1064),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1002),
.A2(n_952),
.B(n_959),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1064),
.B(n_1065),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1043),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1044),
.Y(n_1217)
);

AND2x6_ASAP7_75t_L g1218 ( 
.A(n_1034),
.B(n_1065),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_940),
.A2(n_947),
.B(n_1012),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1012),
.A2(n_996),
.B(n_958),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_994),
.B(n_1030),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1045),
.B(n_1060),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1000),
.Y(n_1223)
);

OA22x2_ASAP7_75t_L g1224 ( 
.A1(n_992),
.A2(n_1001),
.B1(n_1003),
.B2(n_1067),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_985),
.A2(n_990),
.B1(n_981),
.B2(n_986),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1071),
.B(n_1000),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_979),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1000),
.B(n_990),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_948),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_983),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_992),
.B(n_1057),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1072),
.Y(n_1232)
);

HB1xp67_ASAP7_75t_L g1233 ( 
.A(n_900),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_963),
.A2(n_970),
.B(n_974),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1061),
.B(n_1052),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_R g1236 ( 
.A(n_1023),
.B(n_1049),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1052),
.B(n_1055),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1033),
.B(n_1031),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_977),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_975),
.B(n_1016),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1098),
.B(n_1009),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1076),
.A2(n_1144),
.B(n_1165),
.Y(n_1242)
);

OAI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1124),
.A2(n_977),
.B1(n_1015),
.B2(n_1042),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1101),
.A2(n_1047),
.B(n_1059),
.C(n_1063),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1193),
.A2(n_1092),
.B(n_1097),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1239),
.A2(n_1088),
.A3(n_1191),
.B(n_1172),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1194),
.A2(n_1132),
.B1(n_1187),
.B2(n_1170),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1093),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1203),
.A2(n_1222),
.B(n_1087),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1221),
.A2(n_1198),
.A3(n_1082),
.B(n_1225),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1099),
.B(n_1175),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1238),
.A2(n_1083),
.B(n_1180),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_SL g1253 ( 
.A(n_1107),
.B(n_1100),
.Y(n_1253)
);

NAND3x1_ASAP7_75t_L g1254 ( 
.A(n_1164),
.B(n_1202),
.C(n_1160),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1234),
.A2(n_1235),
.A3(n_1220),
.B(n_1219),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1121),
.A2(n_1117),
.B(n_1102),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_SL g1257 ( 
.A1(n_1184),
.A2(n_1151),
.B(n_1128),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1112),
.A2(n_1081),
.B(n_1224),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1182),
.A2(n_1104),
.B(n_1112),
.C(n_1114),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1084),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1113),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1240),
.A2(n_1188),
.B(n_1096),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1235),
.A2(n_1237),
.A3(n_1226),
.B(n_1185),
.Y(n_1263)
);

OA21x2_ASAP7_75t_L g1264 ( 
.A1(n_1131),
.A2(n_1233),
.B(n_1214),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1224),
.A2(n_1090),
.B(n_1094),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1077),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1228),
.A2(n_1183),
.B(n_1085),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1100),
.B(n_1202),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1189),
.A2(n_1197),
.B(n_1196),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1094),
.B(n_1227),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1116),
.A2(n_1148),
.B(n_1163),
.C(n_1147),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1131),
.A2(n_1127),
.B(n_1148),
.Y(n_1272)
);

AO32x2_ASAP7_75t_L g1273 ( 
.A1(n_1150),
.A2(n_1174),
.A3(n_1176),
.B1(n_1156),
.B2(n_1154),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1186),
.B(n_1091),
.Y(n_1274)
);

CKINVDCx16_ASAP7_75t_R g1275 ( 
.A(n_1141),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1137),
.A2(n_1142),
.B(n_1190),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1190),
.A2(n_1095),
.B(n_1079),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1133),
.B(n_1106),
.Y(n_1278)
);

AOI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1115),
.A2(n_1171),
.B1(n_1192),
.B2(n_1177),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1232),
.A2(n_1139),
.A3(n_1157),
.B(n_1230),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1194),
.A2(n_1187),
.B1(n_1166),
.B2(n_1178),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1089),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1109),
.Y(n_1283)
);

CKINVDCx9p33_ASAP7_75t_R g1284 ( 
.A(n_1192),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1229),
.A2(n_1204),
.B(n_1233),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1139),
.A2(n_1218),
.B(n_1111),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_SL g1287 ( 
.A(n_1110),
.B(n_1168),
.Y(n_1287)
);

NAND3x1_ASAP7_75t_L g1288 ( 
.A(n_1091),
.B(n_1161),
.C(n_1145),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1129),
.A2(n_1140),
.B(n_1153),
.C(n_1211),
.Y(n_1289)
);

BUFx4f_ASAP7_75t_SL g1290 ( 
.A(n_1167),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_L g1291 ( 
.A(n_1119),
.B(n_1105),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1218),
.A2(n_1123),
.B(n_1215),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1106),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1119),
.B(n_1173),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1213),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1199),
.B(n_1213),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1212),
.A2(n_1209),
.B1(n_1108),
.B2(n_1216),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1118),
.B(n_1075),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1122),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1126),
.A2(n_1078),
.B(n_1231),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1136),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1075),
.B(n_1086),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1086),
.B(n_1181),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1079),
.A2(n_1095),
.B(n_1169),
.Y(n_1304)
);

INVx5_ASAP7_75t_L g1305 ( 
.A(n_1136),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1125),
.A2(n_1130),
.A3(n_1201),
.B(n_1217),
.Y(n_1306)
);

INVx5_ASAP7_75t_L g1307 ( 
.A(n_1136),
.Y(n_1307)
);

AND2x2_ASAP7_75t_SL g1308 ( 
.A(n_1223),
.B(n_1138),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1205),
.A2(n_1200),
.B(n_1158),
.C(n_1208),
.Y(n_1309)
);

NAND2xp33_ASAP7_75t_SL g1310 ( 
.A(n_1134),
.B(n_1181),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1169),
.A2(n_1209),
.B(n_1212),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1208),
.B(n_1146),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1149),
.A2(n_1210),
.B(n_1135),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1103),
.A2(n_1143),
.B(n_1120),
.C(n_1179),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1103),
.B(n_1143),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1231),
.A2(n_1195),
.B(n_1136),
.Y(n_1316)
);

NAND3xp33_ASAP7_75t_L g1317 ( 
.A(n_1134),
.B(n_1155),
.C(n_1108),
.Y(n_1317)
);

INVx2_ASAP7_75t_SL g1318 ( 
.A(n_1162),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1120),
.B(n_1218),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1231),
.A2(n_1207),
.B1(n_1206),
.B2(n_1218),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1162),
.B(n_1179),
.Y(n_1321)
);

BUFx6f_ASAP7_75t_L g1322 ( 
.A(n_1168),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1218),
.B(n_1152),
.Y(n_1323)
);

AO21x1_ASAP7_75t_L g1324 ( 
.A1(n_1152),
.A2(n_1135),
.B(n_1236),
.Y(n_1324)
);

AOI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1159),
.A2(n_608),
.B1(n_969),
.B2(n_1098),
.C(n_849),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1195),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1195),
.B(n_1080),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1195),
.A2(n_1098),
.B(n_883),
.Y(n_1328)
);

O2A1O1Ixp33_ASAP7_75t_L g1329 ( 
.A1(n_1098),
.A2(n_969),
.B(n_883),
.C(n_882),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1330)
);

A2O1A1Ixp33_ASAP7_75t_L g1331 ( 
.A1(n_1098),
.A2(n_883),
.B(n_882),
.C(n_716),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1098),
.A2(n_733),
.B1(n_724),
.B2(n_1006),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1333)
);

NOR2xp33_ASAP7_75t_L g1334 ( 
.A(n_1098),
.B(n_737),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1098),
.A2(n_883),
.B(n_882),
.C(n_716),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1078),
.Y(n_1337)
);

OR2x2_ASAP7_75t_L g1338 ( 
.A(n_1099),
.B(n_978),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1098),
.A2(n_883),
.B(n_882),
.C(n_716),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1084),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1181),
.B(n_1119),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1093),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1181),
.B(n_1119),
.Y(n_1345)
);

BUFx6f_ASAP7_75t_L g1346 ( 
.A(n_1136),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1084),
.Y(n_1347)
);

CKINVDCx11_ASAP7_75t_R g1348 ( 
.A(n_1093),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1098),
.B(n_886),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1099),
.B(n_889),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1099),
.B(n_889),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1093),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1084),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1110),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1084),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1098),
.A2(n_883),
.B(n_1165),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1084),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1077),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1361)
);

INVxp67_ASAP7_75t_SL g1362 ( 
.A(n_1213),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1098),
.A2(n_733),
.B1(n_724),
.B2(n_1006),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1076),
.A2(n_1098),
.B(n_1222),
.Y(n_1365)
);

OAI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1098),
.A2(n_960),
.B1(n_1194),
.B2(n_946),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1098),
.B(n_886),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1077),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1098),
.B(n_1094),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1098),
.A2(n_883),
.B(n_1165),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1098),
.B(n_1094),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1098),
.B(n_1094),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1181),
.B(n_1119),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1374)
);

O2A1O1Ixp33_ASAP7_75t_L g1375 ( 
.A1(n_1098),
.A2(n_969),
.B(n_883),
.C(n_882),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1376)
);

CKINVDCx9p33_ASAP7_75t_R g1377 ( 
.A(n_1114),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1136),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1098),
.B(n_737),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_SL g1380 ( 
.A1(n_1098),
.A2(n_946),
.B1(n_1163),
.B2(n_1150),
.C(n_1147),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1098),
.B(n_716),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1098),
.A2(n_1239),
.A3(n_1088),
.B(n_1076),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1383)
);

NAND3xp33_ASAP7_75t_SL g1384 ( 
.A(n_1098),
.B(n_717),
.C(n_716),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1181),
.B(n_1119),
.Y(n_1387)
);

OR2x6_ASAP7_75t_L g1388 ( 
.A(n_1146),
.B(n_1027),
.Y(n_1388)
);

NOR2xp33_ASAP7_75t_SL g1389 ( 
.A(n_1098),
.B(n_883),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1391)
);

OAI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1098),
.A2(n_883),
.B(n_1165),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1098),
.B(n_716),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1181),
.B(n_1119),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1098),
.A2(n_960),
.B1(n_1194),
.B2(n_946),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1193),
.A2(n_1015),
.B(n_977),
.Y(n_1396)
);

OAI21xp5_ASAP7_75t_SL g1397 ( 
.A1(n_1098),
.A2(n_1124),
.B(n_883),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_SL g1398 ( 
.A1(n_1098),
.A2(n_883),
.B(n_882),
.C(n_946),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1076),
.A2(n_883),
.B(n_1144),
.Y(n_1399)
);

OA21x2_ASAP7_75t_L g1400 ( 
.A1(n_1193),
.A2(n_1191),
.B(n_1172),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1136),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1098),
.B(n_737),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1098),
.A2(n_883),
.B(n_1165),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1098),
.B(n_737),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_SL g1405 ( 
.A(n_1098),
.B(n_886),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1098),
.B(n_716),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1168),
.B(n_925),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1326),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1389),
.A2(n_1363),
.B1(n_1332),
.B2(n_1366),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1366),
.A2(n_1395),
.B1(n_1389),
.B2(n_1334),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1395),
.A2(n_1404),
.B1(n_1402),
.B2(n_1379),
.Y(n_1411)
);

BUFx8_ASAP7_75t_L g1412 ( 
.A(n_1355),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1260),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1270),
.B(n_1291),
.Y(n_1414)
);

INVxp33_ASAP7_75t_SL g1415 ( 
.A(n_1327),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1261),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1248),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1282),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1247),
.A2(n_1317),
.B1(n_1406),
.B2(n_1381),
.Y(n_1419)
);

CKINVDCx11_ASAP7_75t_R g1420 ( 
.A(n_1348),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1322),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1283),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1325),
.A2(n_1384),
.B1(n_1393),
.B2(n_1349),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1275),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1299),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1367),
.A2(n_1405),
.B1(n_1247),
.B2(n_1317),
.Y(n_1426)
);

BUFx2_ASAP7_75t_SL g1427 ( 
.A(n_1344),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_SL g1428 ( 
.A1(n_1281),
.A2(n_1392),
.B1(n_1358),
.B2(n_1403),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1360),
.Y(n_1429)
);

BUFx6f_ASAP7_75t_L g1430 ( 
.A(n_1305),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1369),
.A2(n_1371),
.B1(n_1372),
.B2(n_1403),
.Y(n_1431)
);

INVx6_ASAP7_75t_L g1432 ( 
.A(n_1293),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1350),
.B(n_1351),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1322),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1340),
.Y(n_1435)
);

NAND2xp33_ASAP7_75t_R g1436 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1266),
.Y(n_1437)
);

INVx6_ASAP7_75t_L g1438 ( 
.A(n_1293),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1347),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1353),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1284),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1397),
.A2(n_1274),
.B1(n_1254),
.B2(n_1279),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1397),
.A2(n_1331),
.B1(n_1339),
.B2(n_1335),
.Y(n_1443)
);

BUFx10_ASAP7_75t_L g1444 ( 
.A(n_1312),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1242),
.A2(n_1376),
.B(n_1399),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1372),
.A2(n_1370),
.B1(n_1392),
.B2(n_1358),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1368),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1354),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_1290),
.Y(n_1449)
);

AOI22x1_ASAP7_75t_L g1450 ( 
.A1(n_1272),
.A2(n_1370),
.B1(n_1257),
.B2(n_1286),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1305),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1286),
.A2(n_1328),
.B1(n_1251),
.B2(n_1281),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1328),
.A2(n_1272),
.B1(n_1265),
.B2(n_1308),
.Y(n_1453)
);

CKINVDCx11_ASAP7_75t_R g1454 ( 
.A(n_1342),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1265),
.A2(n_1258),
.B1(n_1268),
.B2(n_1365),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1356),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1338),
.B(n_1296),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1258),
.A2(n_1365),
.B1(n_1310),
.B2(n_1278),
.Y(n_1458)
);

OAI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1287),
.A2(n_1359),
.B1(n_1295),
.B2(n_1297),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1294),
.Y(n_1460)
);

CKINVDCx16_ASAP7_75t_R g1461 ( 
.A(n_1287),
.Y(n_1461)
);

BUFx12f_ASAP7_75t_L g1462 ( 
.A(n_1322),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1259),
.A2(n_1288),
.B1(n_1329),
.B2(n_1375),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1362),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1271),
.A2(n_1377),
.B(n_1320),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1342),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1315),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1345),
.Y(n_1468)
);

BUFx8_ASAP7_75t_L g1469 ( 
.A(n_1301),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1345),
.B(n_1373),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1380),
.A2(n_1241),
.B1(n_1298),
.B2(n_1297),
.Y(n_1471)
);

CKINVDCx20_ASAP7_75t_R g1472 ( 
.A(n_1253),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1302),
.A2(n_1303),
.B1(n_1394),
.B2(n_1373),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1315),
.Y(n_1474)
);

BUFx4f_ASAP7_75t_SL g1475 ( 
.A(n_1387),
.Y(n_1475)
);

BUFx2_ASAP7_75t_SL g1476 ( 
.A(n_1307),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1321),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1387),
.B(n_1394),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1346),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1346),
.Y(n_1480)
);

OAI21xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1311),
.A2(n_1319),
.B(n_1292),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1380),
.A2(n_1241),
.B1(n_1292),
.B2(n_1267),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1313),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1378),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1273),
.B(n_1318),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1300),
.A2(n_1316),
.B1(n_1269),
.B2(n_1388),
.Y(n_1486)
);

OAI21xp5_ASAP7_75t_SL g1487 ( 
.A1(n_1336),
.A2(n_1383),
.B(n_1352),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1401),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1324),
.A2(n_1398),
.B1(n_1374),
.B2(n_1361),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1364),
.A2(n_1390),
.B1(n_1391),
.B2(n_1385),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1401),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1285),
.B(n_1280),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1280),
.B(n_1263),
.Y(n_1493)
);

CKINVDCx6p67_ASAP7_75t_R g1494 ( 
.A(n_1388),
.Y(n_1494)
);

BUFx12f_ASAP7_75t_L g1495 ( 
.A(n_1388),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1407),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1273),
.A2(n_1323),
.B1(n_1319),
.B2(n_1337),
.Y(n_1497)
);

OAI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1273),
.A2(n_1252),
.B1(n_1249),
.B2(n_1264),
.Y(n_1498)
);

INVx6_ASAP7_75t_L g1499 ( 
.A(n_1407),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1314),
.Y(n_1500)
);

CKINVDCx8_ASAP7_75t_R g1501 ( 
.A(n_1264),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1280),
.Y(n_1502)
);

BUFx3_ASAP7_75t_L g1503 ( 
.A(n_1304),
.Y(n_1503)
);

CKINVDCx11_ASAP7_75t_R g1504 ( 
.A(n_1289),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1309),
.A2(n_1276),
.B1(n_1277),
.B2(n_1243),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1306),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1262),
.A2(n_1400),
.B1(n_1256),
.B2(n_1245),
.Y(n_1507)
);

CKINVDCx11_ASAP7_75t_R g1508 ( 
.A(n_1263),
.Y(n_1508)
);

BUFx4_ASAP7_75t_SL g1509 ( 
.A(n_1263),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1400),
.A2(n_1333),
.B1(n_1386),
.B2(n_1357),
.Y(n_1510)
);

INVx1_ASAP7_75t_SL g1511 ( 
.A(n_1330),
.Y(n_1511)
);

CKINVDCx11_ASAP7_75t_R g1512 ( 
.A(n_1306),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1250),
.A2(n_1382),
.B1(n_1255),
.B2(n_1396),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_SL g1514 ( 
.A1(n_1250),
.A2(n_1382),
.B1(n_1255),
.B2(n_1341),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1306),
.Y(n_1515)
);

INVx2_ASAP7_75t_SL g1516 ( 
.A(n_1255),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1250),
.A2(n_1382),
.B1(n_1343),
.B2(n_1246),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1246),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1246),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1244),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1332),
.A2(n_1098),
.B1(n_1363),
.B2(n_709),
.Y(n_1521)
);

BUFx4f_ASAP7_75t_L g1522 ( 
.A(n_1355),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1260),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1260),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1366),
.A2(n_1395),
.B1(n_1389),
.B2(n_1124),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1332),
.A2(n_1098),
.B1(n_1363),
.B2(n_709),
.Y(n_1526)
);

BUFx12f_ASAP7_75t_L g1527 ( 
.A(n_1348),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1266),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1366),
.A2(n_1124),
.B1(n_1395),
.B2(n_1379),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1362),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1305),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1366),
.A2(n_1395),
.B1(n_1389),
.B2(n_1124),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1326),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1366),
.A2(n_1124),
.B1(n_1395),
.B2(n_1379),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_L g1535 ( 
.A1(n_1366),
.A2(n_1124),
.B1(n_1395),
.B2(n_1379),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1366),
.A2(n_1124),
.B1(n_1395),
.B2(n_1379),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1355),
.Y(n_1537)
);

INVx4_ASAP7_75t_SL g1538 ( 
.A(n_1326),
.Y(n_1538)
);

INVx6_ASAP7_75t_L g1539 ( 
.A(n_1326),
.Y(n_1539)
);

BUFx2_ASAP7_75t_SL g1540 ( 
.A(n_1248),
.Y(n_1540)
);

BUFx2_ASAP7_75t_SL g1541 ( 
.A(n_1248),
.Y(n_1541)
);

INVx6_ASAP7_75t_L g1542 ( 
.A(n_1326),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1366),
.A2(n_1124),
.B1(n_1395),
.B2(n_1379),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1270),
.B(n_889),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1338),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1260),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1366),
.A2(n_1124),
.B1(n_1395),
.B2(n_1379),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1260),
.Y(n_1548)
);

BUFx12f_ASAP7_75t_L g1549 ( 
.A(n_1348),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1355),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1389),
.A2(n_1124),
.B1(n_634),
.B2(n_1332),
.Y(n_1551)
);

CKINVDCx11_ASAP7_75t_R g1552 ( 
.A(n_1355),
.Y(n_1552)
);

INVx6_ASAP7_75t_L g1553 ( 
.A(n_1326),
.Y(n_1553)
);

CKINVDCx6p67_ASAP7_75t_R g1554 ( 
.A(n_1355),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1502),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1493),
.Y(n_1556)
);

NOR2x1_ASAP7_75t_R g1557 ( 
.A(n_1420),
.B(n_1537),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1467),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1474),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1449),
.Y(n_1560)
);

BUFx2_ASAP7_75t_L g1561 ( 
.A(n_1530),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1448),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1414),
.B(n_1457),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1445),
.A2(n_1507),
.B(n_1510),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1413),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1506),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1521),
.A2(n_1526),
.B1(n_1409),
.B2(n_1442),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1416),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1435),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1497),
.B(n_1410),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1433),
.B(n_1478),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1503),
.B(n_1483),
.Y(n_1572)
);

OA21x2_ASAP7_75t_L g1573 ( 
.A1(n_1487),
.A2(n_1490),
.B(n_1489),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1464),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1518),
.Y(n_1575)
);

AO21x1_ASAP7_75t_L g1576 ( 
.A1(n_1463),
.A2(n_1551),
.B(n_1443),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1501),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1505),
.B(n_1516),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1481),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1519),
.Y(n_1580)
);

INVx2_ASAP7_75t_SL g1581 ( 
.A(n_1496),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1492),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1509),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1509),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1439),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1410),
.B(n_1485),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1515),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1450),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1456),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1545),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1523),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1507),
.A2(n_1510),
.B(n_1489),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1524),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1546),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1411),
.B(n_1525),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1548),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1418),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1411),
.B(n_1525),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1529),
.A2(n_1535),
.B(n_1543),
.C(n_1536),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1511),
.Y(n_1600)
);

BUFx12f_ASAP7_75t_L g1601 ( 
.A(n_1552),
.Y(n_1601)
);

OAI21x1_ASAP7_75t_L g1602 ( 
.A1(n_1490),
.A2(n_1486),
.B(n_1482),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1460),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1532),
.B(n_1428),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1512),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1482),
.A2(n_1446),
.B(n_1423),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1513),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1513),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1514),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1514),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1422),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1425),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1498),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1498),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1532),
.A2(n_1534),
.B1(n_1547),
.B2(n_1529),
.Y(n_1615)
);

INVx3_ASAP7_75t_L g1616 ( 
.A(n_1500),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1500),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1424),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1428),
.B(n_1455),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1517),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1495),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1517),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1455),
.B(n_1446),
.Y(n_1623)
);

INVx3_ASAP7_75t_L g1624 ( 
.A(n_1500),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1452),
.B(n_1453),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1453),
.A2(n_1452),
.B(n_1535),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1496),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1544),
.B(n_1431),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_SL g1629 ( 
.A1(n_1461),
.A2(n_1441),
.B1(n_1472),
.B2(n_1534),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1508),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1459),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1470),
.B(n_1415),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1477),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1459),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1536),
.A2(n_1547),
.B(n_1543),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1419),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1423),
.A2(n_1426),
.B(n_1471),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1426),
.B(n_1458),
.Y(n_1638)
);

NOR2xp33_ASAP7_75t_L g1639 ( 
.A(n_1440),
.B(n_1466),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1520),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1431),
.B(n_1471),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_SL g1642 ( 
.A1(n_1473),
.A2(n_1444),
.B1(n_1475),
.B2(n_1436),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1419),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1436),
.A2(n_1465),
.B1(n_1458),
.B2(n_1504),
.Y(n_1644)
);

AO21x2_ASAP7_75t_L g1645 ( 
.A1(n_1491),
.A2(n_1476),
.B(n_1494),
.Y(n_1645)
);

INVx1_ASAP7_75t_SL g1646 ( 
.A(n_1447),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1499),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1468),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1437),
.B(n_1528),
.C(n_1469),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1430),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1469),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1408),
.A2(n_1421),
.B(n_1434),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1408),
.A2(n_1421),
.B(n_1434),
.Y(n_1653)
);

INVxp67_ASAP7_75t_L g1654 ( 
.A(n_1427),
.Y(n_1654)
);

AOI21x1_ASAP7_75t_L g1655 ( 
.A1(n_1444),
.A2(n_1451),
.B(n_1531),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1429),
.A2(n_1454),
.B1(n_1475),
.B2(n_1522),
.Y(n_1656)
);

CKINVDCx11_ASAP7_75t_R g1657 ( 
.A(n_1527),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1417),
.B(n_1540),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1451),
.B(n_1432),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1484),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1479),
.A2(n_1480),
.B(n_1484),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1484),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1488),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1541),
.B(n_1550),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1432),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1438),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1538),
.B(n_1438),
.Y(n_1667)
);

AND2x4_ASAP7_75t_L g1668 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1668)
);

BUFx2_ASAP7_75t_L g1669 ( 
.A(n_1462),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1533),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1533),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1538),
.Y(n_1672)
);

A2O1A1Ixp33_ASAP7_75t_L g1673 ( 
.A1(n_1599),
.A2(n_1635),
.B(n_1595),
.C(n_1598),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1563),
.B(n_1542),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1587),
.B(n_1554),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1595),
.A2(n_1522),
.B(n_1533),
.C(n_1539),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_L g1677 ( 
.A(n_1649),
.B(n_1412),
.Y(n_1677)
);

OAI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1615),
.A2(n_1539),
.B1(n_1542),
.B2(n_1553),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1628),
.B(n_1542),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1587),
.B(n_1553),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1586),
.B(n_1549),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_SL g1683 ( 
.A1(n_1576),
.A2(n_1412),
.B(n_1644),
.Y(n_1683)
);

CKINVDCx6p67_ASAP7_75t_R g1684 ( 
.A(n_1601),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1644),
.A2(n_1567),
.B1(n_1629),
.B2(n_1642),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1571),
.B(n_1630),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1561),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1606),
.A2(n_1598),
.B(n_1602),
.Y(n_1688)
);

AO22x2_ASAP7_75t_L g1689 ( 
.A1(n_1607),
.A2(n_1608),
.B1(n_1609),
.B2(n_1610),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1630),
.B(n_1605),
.Y(n_1690)
);

AOI21xp33_ASAP7_75t_L g1691 ( 
.A1(n_1576),
.A2(n_1604),
.B(n_1625),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_L g1693 ( 
.A(n_1640),
.B(n_1643),
.C(n_1636),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1605),
.B(n_1570),
.Y(n_1694)
);

AND2x2_ASAP7_75t_SL g1695 ( 
.A(n_1579),
.B(n_1570),
.Y(n_1695)
);

AOI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1619),
.A2(n_1643),
.B1(n_1636),
.B2(n_1623),
.C(n_1588),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1619),
.B(n_1603),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1588),
.A2(n_1641),
.B(n_1637),
.Y(n_1698)
);

NOR2xp33_ASAP7_75t_L g1699 ( 
.A(n_1631),
.B(n_1634),
.Y(n_1699)
);

OA21x2_ASAP7_75t_L g1700 ( 
.A1(n_1592),
.A2(n_1564),
.B(n_1613),
.Y(n_1700)
);

AO32x2_ASAP7_75t_L g1701 ( 
.A1(n_1574),
.A2(n_1581),
.A3(n_1627),
.B1(n_1620),
.B2(n_1622),
.Y(n_1701)
);

OAI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1641),
.A2(n_1637),
.B(n_1640),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1565),
.B(n_1568),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1583),
.B(n_1584),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1638),
.A2(n_1579),
.B(n_1613),
.C(n_1614),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1569),
.B(n_1585),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1637),
.B(n_1638),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1572),
.B(n_1583),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1626),
.A2(n_1638),
.B1(n_1637),
.B2(n_1649),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1590),
.B(n_1558),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1577),
.B(n_1659),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1585),
.B(n_1589),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1589),
.B(n_1591),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1614),
.A2(n_1577),
.B(n_1624),
.C(n_1616),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1654),
.A2(n_1626),
.B1(n_1656),
.B2(n_1646),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1626),
.A2(n_1573),
.B(n_1653),
.Y(n_1716)
);

CKINVDCx20_ASAP7_75t_R g1717 ( 
.A(n_1560),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1582),
.B(n_1574),
.Y(n_1718)
);

NOR2x1_ASAP7_75t_SL g1719 ( 
.A(n_1645),
.B(n_1659),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1566),
.A2(n_1580),
.B(n_1575),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1558),
.B(n_1559),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1601),
.Y(n_1722)
);

OAI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1626),
.A2(n_1573),
.B(n_1652),
.Y(n_1723)
);

A2O1A1Ixp33_ASAP7_75t_L g1724 ( 
.A1(n_1577),
.A2(n_1616),
.B(n_1617),
.C(n_1624),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1562),
.B(n_1593),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1632),
.A2(n_1668),
.B1(n_1664),
.B2(n_1670),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1582),
.B(n_1594),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1596),
.B(n_1556),
.Y(n_1728)
);

O2A1O1Ixp33_ASAP7_75t_L g1729 ( 
.A1(n_1648),
.A2(n_1616),
.B(n_1617),
.C(n_1624),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1668),
.A2(n_1670),
.B1(n_1658),
.B2(n_1621),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1660),
.B(n_1662),
.Y(n_1731)
);

NAND4xp25_ASAP7_75t_L g1732 ( 
.A(n_1621),
.B(n_1669),
.C(n_1639),
.D(n_1559),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1666),
.B(n_1647),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1575),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1580),
.Y(n_1735)
);

BUFx12f_ASAP7_75t_L g1736 ( 
.A(n_1722),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1720),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1720),
.Y(n_1738)
);

NAND2x1_ASAP7_75t_SL g1739 ( 
.A(n_1709),
.B(n_1578),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1720),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1734),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1700),
.B(n_1578),
.Y(n_1742)
);

BUFx2_ASAP7_75t_L g1743 ( 
.A(n_1701),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1555),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_SL g1745 ( 
.A(n_1695),
.B(n_1647),
.Y(n_1745)
);

INVx2_ASAP7_75t_SL g1746 ( 
.A(n_1735),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1689),
.B(n_1697),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1716),
.B(n_1723),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1688),
.B(n_1578),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1689),
.B(n_1566),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1713),
.Y(n_1751)
);

AOI22xp5_ASAP7_75t_L g1752 ( 
.A1(n_1685),
.A2(n_1668),
.B1(n_1670),
.B2(n_1667),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1689),
.B(n_1600),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1707),
.B(n_1701),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1711),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1703),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1719),
.B(n_1572),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1701),
.B(n_1600),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1717),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1708),
.B(n_1653),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1706),
.Y(n_1761)
);

AOI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1673),
.A2(n_1669),
.B1(n_1612),
.B2(n_1597),
.C(n_1611),
.Y(n_1762)
);

BUFx2_ASAP7_75t_L g1763 ( 
.A(n_1687),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1712),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1718),
.B(n_1661),
.Y(n_1765)
);

BUFx12f_ASAP7_75t_L g1766 ( 
.A(n_1722),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1743),
.B(n_1692),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1738),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1741),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1738),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1754),
.B(n_1694),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1741),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1750),
.B(n_1725),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1736),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1754),
.B(n_1708),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1752),
.A2(n_1673),
.B1(n_1691),
.B2(n_1702),
.C(n_1696),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1754),
.B(n_1708),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1754),
.B(n_1695),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1743),
.B(n_1728),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1762),
.A2(n_1693),
.B1(n_1683),
.B2(n_1715),
.C(n_1699),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1737),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1744),
.B(n_1705),
.Y(n_1782)
);

AOI33xp33_ASAP7_75t_L g1783 ( 
.A1(n_1748),
.A2(n_1686),
.A3(n_1690),
.B1(n_1682),
.B2(n_1681),
.B3(n_1680),
.Y(n_1783)
);

INVx4_ASAP7_75t_L g1784 ( 
.A(n_1736),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1752),
.A2(n_1693),
.B1(n_1676),
.B2(n_1677),
.C(n_1679),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1747),
.B(n_1727),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1747),
.B(n_1710),
.Y(n_1787)
);

INVxp67_ASAP7_75t_L g1788 ( 
.A(n_1753),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1753),
.B(n_1740),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1752),
.A2(n_1678),
.B1(n_1762),
.B2(n_1745),
.Y(n_1790)
);

BUFx2_ASAP7_75t_L g1791 ( 
.A(n_1739),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1739),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1746),
.Y(n_1793)
);

AOI33xp33_ASAP7_75t_L g1794 ( 
.A1(n_1748),
.A2(n_1704),
.A3(n_1731),
.B1(n_1729),
.B2(n_1733),
.B3(n_1726),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_SL g1795 ( 
.A(n_1736),
.B(n_1724),
.Y(n_1795)
);

OR2x6_ASAP7_75t_L g1796 ( 
.A(n_1755),
.B(n_1711),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1740),
.Y(n_1797)
);

INVx3_ASAP7_75t_L g1798 ( 
.A(n_1760),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1744),
.B(n_1721),
.Y(n_1799)
);

OAI21xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1745),
.A2(n_1676),
.B(n_1732),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1739),
.Y(n_1801)
);

AND2x4_ASAP7_75t_L g1802 ( 
.A(n_1757),
.B(n_1704),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1742),
.B(n_1714),
.Y(n_1803)
);

INVx3_ASAP7_75t_L g1804 ( 
.A(n_1760),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1788),
.B(n_1751),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1791),
.B(n_1748),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1791),
.B(n_1742),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1792),
.B(n_1742),
.Y(n_1808)
);

AND2x4_ASAP7_75t_SL g1809 ( 
.A(n_1784),
.B(n_1755),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1788),
.B(n_1751),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1797),
.Y(n_1811)
);

OR2x6_ASAP7_75t_L g1812 ( 
.A(n_1796),
.B(n_1755),
.Y(n_1812)
);

INVxp67_ASAP7_75t_L g1813 ( 
.A(n_1782),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1779),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1787),
.B(n_1756),
.Y(n_1815)
);

OR2x2_ASAP7_75t_L g1816 ( 
.A(n_1767),
.B(n_1765),
.Y(n_1816)
);

OR2x2_ASAP7_75t_L g1817 ( 
.A(n_1767),
.B(n_1765),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1787),
.B(n_1756),
.Y(n_1818)
);

BUFx2_ASAP7_75t_L g1819 ( 
.A(n_1792),
.Y(n_1819)
);

INVx2_ASAP7_75t_SL g1820 ( 
.A(n_1793),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1787),
.B(n_1756),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1768),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1767),
.B(n_1765),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1799),
.B(n_1761),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1801),
.B(n_1803),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1769),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1799),
.B(n_1761),
.Y(n_1827)
);

INVxp67_ASAP7_75t_SL g1828 ( 
.A(n_1793),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1768),
.Y(n_1829)
);

AND2x4_ASAP7_75t_L g1830 ( 
.A(n_1804),
.B(n_1757),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1799),
.B(n_1761),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1768),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1801),
.B(n_1758),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1769),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1804),
.B(n_1757),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1782),
.B(n_1764),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1803),
.B(n_1775),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1786),
.B(n_1764),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1803),
.B(n_1758),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1775),
.B(n_1758),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1770),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1775),
.B(n_1749),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1772),
.Y(n_1843)
);

HB1xp67_ASAP7_75t_L g1844 ( 
.A(n_1779),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1814),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1814),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1837),
.B(n_1778),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1820),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1813),
.B(n_1836),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_L g1850 ( 
.A(n_1819),
.B(n_1784),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1813),
.B(n_1771),
.Y(n_1851)
);

INVxp67_ASAP7_75t_SL g1852 ( 
.A(n_1844),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1836),
.B(n_1771),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1837),
.B(n_1778),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1805),
.A2(n_1776),
.B1(n_1780),
.B2(n_1800),
.C(n_1785),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1837),
.B(n_1778),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1844),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1815),
.B(n_1789),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1826),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1815),
.B(n_1789),
.Y(n_1860)
);

OR2x2_ASAP7_75t_L g1861 ( 
.A(n_1818),
.B(n_1789),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1825),
.B(n_1771),
.Y(n_1862)
);

NAND2x1_ASAP7_75t_L g1863 ( 
.A(n_1819),
.B(n_1802),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1825),
.B(n_1777),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1820),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1820),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1805),
.B(n_1786),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1826),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1810),
.B(n_1786),
.Y(n_1869)
);

NOR2xp33_ASAP7_75t_L g1870 ( 
.A(n_1810),
.B(n_1684),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1812),
.B(n_1804),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1825),
.B(n_1777),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1818),
.B(n_1773),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1834),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1839),
.B(n_1777),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1822),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1834),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1809),
.B(n_1736),
.Y(n_1878)
);

INVx1_ASAP7_75t_SL g1879 ( 
.A(n_1809),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1821),
.B(n_1773),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1839),
.B(n_1802),
.Y(n_1881)
);

OR2x2_ASAP7_75t_L g1882 ( 
.A(n_1821),
.B(n_1824),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1839),
.B(n_1802),
.Y(n_1883)
);

BUFx6f_ASAP7_75t_L g1884 ( 
.A(n_1812),
.Y(n_1884)
);

AO221x1_ASAP7_75t_L g1885 ( 
.A1(n_1811),
.A2(n_1798),
.B1(n_1804),
.B2(n_1763),
.C(n_1663),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1842),
.B(n_1802),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1843),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1842),
.B(n_1802),
.Y(n_1888)
);

NOR2xp33_ASAP7_75t_L g1889 ( 
.A(n_1870),
.B(n_1766),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1847),
.B(n_1806),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1855),
.B(n_1783),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1851),
.B(n_1816),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1845),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1845),
.Y(n_1894)
);

NOR3xp33_ASAP7_75t_L g1895 ( 
.A(n_1855),
.B(n_1784),
.C(n_1776),
.Y(n_1895)
);

NAND2x1p5_ASAP7_75t_L g1896 ( 
.A(n_1850),
.B(n_1784),
.Y(n_1896)
);

OAI211xp5_ASAP7_75t_L g1897 ( 
.A1(n_1850),
.A2(n_1780),
.B(n_1800),
.C(n_1790),
.Y(n_1897)
);

OR2x2_ASAP7_75t_L g1898 ( 
.A(n_1851),
.B(n_1816),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1849),
.B(n_1817),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1847),
.B(n_1806),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_SL g1901 ( 
.A(n_1879),
.B(n_1557),
.Y(n_1901)
);

NOR3xp33_ASAP7_75t_L g1902 ( 
.A(n_1879),
.B(n_1784),
.C(n_1785),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1852),
.Y(n_1903)
);

OAI221xp5_ASAP7_75t_L g1904 ( 
.A1(n_1863),
.A2(n_1812),
.B1(n_1795),
.B2(n_1790),
.C(n_1774),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1849),
.B(n_1794),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1852),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1867),
.B(n_1817),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1854),
.B(n_1806),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1854),
.B(n_1842),
.Y(n_1909)
);

NOR2xp67_ASAP7_75t_R g1910 ( 
.A(n_1884),
.B(n_1766),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1878),
.A2(n_1557),
.B(n_1663),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1856),
.B(n_1833),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1856),
.B(n_1824),
.Y(n_1913)
);

NOR2x1_ASAP7_75t_L g1914 ( 
.A(n_1846),
.B(n_1774),
.Y(n_1914)
);

OR2x2_ASAP7_75t_L g1915 ( 
.A(n_1867),
.B(n_1823),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1862),
.B(n_1833),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1884),
.A2(n_1795),
.B1(n_1812),
.B2(n_1809),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1862),
.B(n_1833),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1869),
.B(n_1827),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1864),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1869),
.B(n_1827),
.Y(n_1921)
);

NAND2x1p5_ASAP7_75t_L g1922 ( 
.A(n_1863),
.B(n_1663),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1884),
.B(n_1766),
.Y(n_1923)
);

AOI211xp5_ASAP7_75t_L g1924 ( 
.A1(n_1884),
.A2(n_1774),
.B(n_1749),
.C(n_1675),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1846),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1922),
.B(n_1864),
.Y(n_1926)
);

OAI33xp33_ASAP7_75t_L g1927 ( 
.A1(n_1891),
.A2(n_1857),
.A3(n_1865),
.B1(n_1866),
.B2(n_1848),
.B3(n_1859),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1925),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1922),
.B(n_1872),
.Y(n_1929)
);

AOI21xp5_ASAP7_75t_L g1930 ( 
.A1(n_1897),
.A2(n_1857),
.B(n_1618),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1895),
.B(n_1872),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1911),
.A2(n_1885),
.B(n_1759),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1903),
.Y(n_1933)
);

AOI221xp5_ASAP7_75t_L g1934 ( 
.A1(n_1905),
.A2(n_1884),
.B1(n_1885),
.B2(n_1880),
.C(n_1848),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_L g1935 ( 
.A(n_1901),
.B(n_1766),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1912),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1893),
.B(n_1875),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1890),
.B(n_1875),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1904),
.A2(n_1884),
.B1(n_1880),
.B2(n_1866),
.C(n_1865),
.Y(n_1939)
);

OAI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1924),
.A2(n_1917),
.B1(n_1914),
.B2(n_1896),
.Y(n_1940)
);

NOR2xp67_ASAP7_75t_L g1941 ( 
.A(n_1890),
.B(n_1848),
.Y(n_1941)
);

NOR4xp25_ASAP7_75t_L g1942 ( 
.A(n_1906),
.B(n_1865),
.C(n_1866),
.D(n_1874),
.Y(n_1942)
);

OAI21xp5_ASAP7_75t_L g1943 ( 
.A1(n_1902),
.A2(n_1812),
.B(n_1873),
.Y(n_1943)
);

OAI221xp5_ASAP7_75t_L g1944 ( 
.A1(n_1923),
.A2(n_1911),
.B1(n_1896),
.B2(n_1894),
.C(n_1889),
.Y(n_1944)
);

AOI22xp5_ASAP7_75t_L g1945 ( 
.A1(n_1920),
.A2(n_1812),
.B1(n_1871),
.B2(n_1796),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1900),
.B(n_1881),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1900),
.B(n_1881),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1908),
.B(n_1883),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1899),
.B(n_1882),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1920),
.A2(n_1871),
.B1(n_1796),
.B2(n_1883),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1912),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_SL g1952 ( 
.A1(n_1935),
.A2(n_1896),
.B(n_1663),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1951),
.Y(n_1953)
);

OAI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1930),
.A2(n_1910),
.B1(n_1919),
.B2(n_1921),
.C(n_1899),
.Y(n_1954)
);

AOI322xp5_ASAP7_75t_L g1955 ( 
.A1(n_1931),
.A2(n_1908),
.A3(n_1918),
.B1(n_1916),
.B2(n_1909),
.C1(n_1913),
.C2(n_1808),
.Y(n_1955)
);

A2O1A1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1932),
.A2(n_1940),
.B(n_1939),
.C(n_1934),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1937),
.B(n_1907),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1942),
.B(n_1916),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1935),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1949),
.B(n_1907),
.Y(n_1960)
);

AOI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1927),
.A2(n_1871),
.B1(n_1915),
.B2(n_1918),
.Y(n_1961)
);

OAI21xp33_ASAP7_75t_L g1962 ( 
.A1(n_1943),
.A2(n_1915),
.B(n_1898),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1928),
.Y(n_1963)
);

XOR2x2_ASAP7_75t_L g1964 ( 
.A(n_1944),
.B(n_1651),
.Y(n_1964)
);

OAI22xp5_ASAP7_75t_L g1965 ( 
.A1(n_1941),
.A2(n_1936),
.B1(n_1949),
.B2(n_1933),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1936),
.Y(n_1966)
);

AOI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1926),
.A2(n_1909),
.B1(n_1871),
.B2(n_1808),
.Y(n_1967)
);

NOR2xp67_ASAP7_75t_L g1968 ( 
.A(n_1926),
.B(n_1892),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1946),
.B(n_1886),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1938),
.B(n_1892),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1946),
.Y(n_1971)
);

OAI222xp33_ASAP7_75t_L g1972 ( 
.A1(n_1950),
.A2(n_1898),
.B1(n_1860),
.B2(n_1861),
.C1(n_1858),
.C2(n_1882),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1956),
.A2(n_1929),
.B(n_1945),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1966),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1971),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1959),
.B(n_1657),
.Y(n_1976)
);

OAI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1958),
.A2(n_1929),
.B(n_1947),
.Y(n_1977)
);

OAI22xp33_ASAP7_75t_SL g1978 ( 
.A1(n_1958),
.A2(n_1858),
.B1(n_1860),
.B2(n_1861),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1960),
.Y(n_1979)
);

AOI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1968),
.A2(n_1954),
.B1(n_1962),
.B2(n_1964),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1953),
.B(n_1938),
.Y(n_1981)
);

OA21x2_ASAP7_75t_L g1982 ( 
.A1(n_1963),
.A2(n_1876),
.B(n_1868),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_SL g1983 ( 
.A1(n_1954),
.A2(n_1948),
.B1(n_1947),
.B2(n_1759),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1970),
.Y(n_1984)
);

NOR3xp33_ASAP7_75t_SL g1985 ( 
.A(n_1973),
.B(n_1965),
.C(n_1972),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1980),
.A2(n_1961),
.B1(n_1967),
.B2(n_1957),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1976),
.B(n_1952),
.Y(n_1987)
);

NOR2xp33_ASAP7_75t_L g1988 ( 
.A(n_1979),
.B(n_1965),
.Y(n_1988)
);

NOR3xp33_ASAP7_75t_L g1989 ( 
.A(n_1983),
.B(n_1969),
.C(n_1621),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1984),
.B(n_1955),
.Y(n_1990)
);

AOI211xp5_ASAP7_75t_L g1991 ( 
.A1(n_1978),
.A2(n_1663),
.B(n_1948),
.C(n_1668),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1982),
.Y(n_1992)
);

NAND3xp33_ASAP7_75t_L g1993 ( 
.A(n_1977),
.B(n_1876),
.C(n_1868),
.Y(n_1993)
);

AOI221xp5_ASAP7_75t_L g1994 ( 
.A1(n_1975),
.A2(n_1876),
.B1(n_1887),
.B2(n_1877),
.C(n_1874),
.Y(n_1994)
);

NAND3xp33_ASAP7_75t_SL g1995 ( 
.A(n_1981),
.B(n_1717),
.C(n_1873),
.Y(n_1995)
);

AOI222xp33_ASAP7_75t_L g1996 ( 
.A1(n_1986),
.A2(n_1974),
.B1(n_1828),
.B2(n_1982),
.C1(n_1807),
.C2(n_1808),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_R g1997 ( 
.A(n_1988),
.B(n_1671),
.Y(n_1997)
);

AOI222xp33_ASAP7_75t_L g1998 ( 
.A1(n_1995),
.A2(n_1828),
.B1(n_1807),
.B2(n_1887),
.C1(n_1877),
.C2(n_1859),
.Y(n_1998)
);

AOI222xp33_ASAP7_75t_L g1999 ( 
.A1(n_1990),
.A2(n_1807),
.B1(n_1853),
.B2(n_1674),
.C1(n_1749),
.C2(n_1781),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1992),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1993),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1985),
.A2(n_1853),
.B1(n_1823),
.B2(n_1830),
.Y(n_2002)
);

INVx1_ASAP7_75t_SL g2003 ( 
.A(n_1997),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_2000),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_2001),
.Y(n_2005)
);

AOI21xp33_ASAP7_75t_L g2006 ( 
.A1(n_1996),
.A2(n_1987),
.B(n_1998),
.Y(n_2006)
);

OAI211xp5_ASAP7_75t_L g2007 ( 
.A1(n_1999),
.A2(n_1989),
.B(n_1991),
.C(n_1994),
.Y(n_2007)
);

OAI211xp5_ASAP7_75t_L g2008 ( 
.A1(n_2002),
.A2(n_1672),
.B(n_1730),
.C(n_1886),
.Y(n_2008)
);

OAI321xp33_ASAP7_75t_L g2009 ( 
.A1(n_2001),
.A2(n_1672),
.A3(n_1796),
.B1(n_1888),
.B2(n_1655),
.C(n_1838),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_2004),
.Y(n_2010)
);

NAND4xp75_ASAP7_75t_L g2011 ( 
.A(n_2005),
.B(n_1888),
.C(n_1661),
.D(n_1840),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_2003),
.B(n_1830),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_2009),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_2006),
.B(n_1840),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_2007),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2014),
.Y(n_2016)
);

AND2x4_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_2008),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_2012),
.B(n_1830),
.Y(n_2018)
);

XNOR2xp5_ASAP7_75t_L g2019 ( 
.A(n_2016),
.B(n_2015),
.Y(n_2019)
);

AO22x2_ASAP7_75t_L g2020 ( 
.A1(n_2019),
.A2(n_2017),
.B1(n_2013),
.B2(n_2012),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2020),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_2020),
.A2(n_2015),
.B1(n_2017),
.B2(n_2013),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_SL g2023 ( 
.A1(n_2021),
.A2(n_2011),
.B1(n_2018),
.B2(n_1667),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_2022),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_SL g2025 ( 
.A1(n_2024),
.A2(n_1655),
.B(n_1831),
.Y(n_2025)
);

AOI22xp33_ASAP7_75t_L g2026 ( 
.A1(n_2023),
.A2(n_1667),
.B1(n_1830),
.B2(n_1835),
.Y(n_2026)
);

AO21x2_ASAP7_75t_L g2027 ( 
.A1(n_2025),
.A2(n_1832),
.B(n_1822),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2027),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2028),
.Y(n_2029)
);

OAI221xp5_ASAP7_75t_R g2030 ( 
.A1(n_2029),
.A2(n_2026),
.B1(n_1829),
.B2(n_1822),
.C(n_1841),
.Y(n_2030)
);

AOI211xp5_ASAP7_75t_L g2031 ( 
.A1(n_2030),
.A2(n_1667),
.B(n_1665),
.C(n_1650),
.Y(n_2031)
);


endmodule