module real_jpeg_6598_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_0),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_0),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_0),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_0),
.B(n_205),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_1),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_20)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_2),
.Y(n_167)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_2),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_2),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_2),
.Y(n_322)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_3),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_3),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_3),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_3),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_4),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_4),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_4),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_4),
.B(n_350),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_4),
.B(n_85),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_4),
.B(n_261),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_5),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_5),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g289 ( 
.A(n_5),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_5),
.B(n_315),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_5),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_6),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_6),
.B(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_6),
.B(n_109),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_6),
.B(n_71),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_6),
.B(n_189),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_6),
.B(n_371),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_6),
.B(n_214),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_7),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_7),
.B(n_111),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_7),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_7),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_7),
.B(n_186),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_7),
.B(n_355),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_7),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_7),
.B(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_8),
.Y(n_118)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_10),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_10),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_10),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_10),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_10),
.B(n_186),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_10),
.B(n_71),
.Y(n_410)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_11),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_11),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_11),
.Y(n_295)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_13),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_14),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_14),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_14),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_14),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_14),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_14),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_14),
.B(n_418),
.Y(n_417)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_16),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_16),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_16),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_16),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_16),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_16),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_16),
.B(n_259),
.Y(n_258)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_18),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_18),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_18),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_18),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_18),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_19),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_19),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_19),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_19),
.B(n_71),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_19),
.B(n_139),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_19),
.B(n_385),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_19),
.B(n_398),
.Y(n_397)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_125),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_123),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_104),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_28),
.B(n_104),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_87),
.C(n_88),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_29),
.A2(n_30),
.B1(n_523),
.B2(n_524),
.Y(n_522)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_60),
.C(n_75),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_31),
.A2(n_32),
.B1(n_504),
.B2(n_506),
.Y(n_503)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_44),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_38),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_38),
.C(n_44),
.Y(n_87)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_37),
.Y(n_144)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_37),
.Y(n_268)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_42),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_42),
.Y(n_263)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_43),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_43),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_50),
.C(n_57),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_45),
.B(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_49),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_50),
.A2(n_51),
.B1(n_57),
.B2(n_58),
.Y(n_494)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_55),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_55),
.Y(n_212)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_56),
.Y(n_278)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_60),
.A2(n_75),
.B1(n_76),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_60),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_69),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g499 ( 
.A(n_61),
.B(n_500),
.Y(n_499)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_63),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_64),
.A2(n_65),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_64),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_500)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_65),
.B(n_200),
.C(n_204),
.Y(n_501)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_67),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_68),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_83),
.C(n_86),
.Y(n_93)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx5_ASAP7_75t_L g351 ( 
.A(n_72),
.Y(n_351)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_73),
.Y(n_217)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_74),
.Y(n_382)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_81),
.B1(n_82),
.B2(n_86),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_84),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_97),
.C(n_100),
.Y(n_106)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_85),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_87),
.B(n_88),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_93),
.C(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_100),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_96),
.A2(n_97),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_99),
.Y(n_202)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_122),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_120),
.B2(n_121),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_119),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g400 ( 
.A(n_118),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_521),
.B(n_526),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_487),
.B(n_518),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_299),
.B(n_486),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_244),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_129),
.B(n_244),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g529 ( 
.A(n_129),
.Y(n_529)
);

FAx1_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_198),
.CI(n_227),
.CON(n_129),
.SN(n_129)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_130),
.B(n_198),
.C(n_227),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_169),
.C(n_180),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_131),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_145),
.C(n_156),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_132),
.B(n_472),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_133),
.B(n_138),
.C(n_141),
.Y(n_179)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_135),
.Y(n_224)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_145),
.A2(n_146),
.B1(n_156),
.B2(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_154),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_147),
.B(n_154),
.Y(n_462)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_149),
.B(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_150),
.B(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_156),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_157),
.B(n_159),
.C(n_165),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_164),
.B1(n_165),
.B2(n_168),
.Y(n_158)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_164),
.B(n_204),
.C(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_164),
.A2(n_165),
.B1(n_204),
.B2(n_208),
.Y(n_240)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_169),
.B(n_180),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_174),
.B1(n_177),
.B2(n_178),
.Y(n_170)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_171),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_174),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_174),
.B(n_177),
.C(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_178),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_178),
.B(n_232),
.C(n_237),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_192),
.C(n_194),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_181),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_188),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_182),
.B(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_185),
.B(n_188),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_187),
.Y(n_416)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_191),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_192),
.B(n_194),
.Y(n_281)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_209),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_199),
.B(n_210),
.C(n_218),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_204),
.Y(n_208)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_207),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_218),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_216),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_216),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_213),
.B(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_214),
.Y(n_366)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_220),
.B(n_223),
.C(n_225),
.Y(n_502)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_229),
.B(n_231),
.C(n_238),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_233),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_242),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.C(n_251),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_246),
.B(n_249),
.Y(n_482)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_251),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_279),
.C(n_282),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_253),
.B(n_475),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.C(n_264),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_254),
.A2(n_255),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_257),
.A2(n_258),
.B(n_260),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_257),
.B(n_264),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.C(n_274),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_430)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_273),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_274),
.B(n_430),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_275),
.B(n_366),
.Y(n_365)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_278),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g475 ( 
.A1(n_279),
.A2(n_280),
.B1(n_282),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_282),
.Y(n_476)
);

MAJx2_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_294),
.C(n_296),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_284),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.C(n_292),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_285),
.B(n_442),
.Y(n_441)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_289),
.A2(n_292),
.B1(n_293),
.B2(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_289),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_294),
.B(n_296),
.Y(n_464)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_480),
.B(n_485),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_467),
.B(n_479),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_449),
.B(n_466),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_423),
.B(n_448),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_391),
.B(n_422),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_358),
.B(n_390),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_341),
.B(n_357),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_324),
.B(n_340),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_320),
.B(n_323),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_316),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_314),
.Y(n_325)
);

INVx4_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_325),
.B(n_326),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_328),
.B1(n_332),
.B2(n_333),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_335),
.C(n_338),
.Y(n_356)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_330),
.Y(n_347)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_334),
.A2(n_335),
.B1(n_338),
.B2(n_339),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_356),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_356),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_347),
.C(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_346),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_348),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_352),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_376),
.C(n_377),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_354),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_359),
.B(n_361),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_374),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_375),
.C(n_378),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_363),
.B(n_365),
.C(n_367),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_369),
.B1(n_370),
.B2(n_373),
.Y(n_367)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_368),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_369),
.B(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_383),
.Y(n_378)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_387),
.C(n_388),
.Y(n_420)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_384),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_383)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_384),
.Y(n_388)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_387),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_392),
.B(n_421),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_421),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_403),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_402),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_394),
.B(n_402),
.C(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_401),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_401),
.B(n_437),
.C(n_438),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_411),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_413),
.C(n_419),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_410),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_406),
.B(n_409),
.C(n_410),
.Y(n_434)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_413),
.B1(n_419),
.B2(n_420),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_417),
.Y(n_433)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_446),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_446),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_435),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_427),
.C(n_435),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_458),
.C(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_433),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_434),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_439),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_440),
.C(n_445),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_444),
.B2(n_445),
.Y(n_439)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_440),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_441),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_465),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_465),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_456),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_455),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_452),
.B(n_455),
.C(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_453),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_461),
.C(n_463),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_468),
.B(n_477),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_468),
.B(n_477),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_470),
.Y(n_468)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_469),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_474),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_474),
.C(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_483),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_481),
.B(n_483),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_515),
.Y(n_487)
);

OAI21xp33_ASAP7_75t_L g518 ( 
.A1(n_488),
.A2(n_519),
.B(n_520),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_508),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_489),
.B(n_508),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_490),
.A2(n_491),
.B1(n_497),
.B2(n_507),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_490),
.B(n_498),
.C(n_503),
.Y(n_525)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.C(n_495),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_510),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_493),
.A2(n_495),
.B1(n_496),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_497),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_503),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_501),
.C(n_502),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_513),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_501),
.B(n_502),
.Y(n_513)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_504),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_512),
.C(n_514),
.Y(n_508)
);

FAx1_ASAP7_75t_L g516 ( 
.A(n_509),
.B(n_512),
.CI(n_514),
.CON(n_516),
.SN(n_516)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_516),
.B(n_517),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_517),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_516),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_522),
.B(n_525),
.Y(n_526)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_523),
.Y(n_524)
);


endmodule