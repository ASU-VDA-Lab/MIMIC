module fake_jpeg_11919_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_38),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_29),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

HAxp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_0),
.CON(n_60),
.SN(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_0),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_53),
.B1(n_52),
.B2(n_43),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_66),
.A2(n_75),
.B1(n_78),
.B2(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_77),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_53),
.B1(n_54),
.B2(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_50),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_42),
.B1(n_44),
.B2(n_41),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_93),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_81),
.Y(n_109)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_84),
.B(n_95),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_2),
.B(n_3),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_89),
.Y(n_104)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_94),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

NAND4xp25_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_22),
.C(n_35),
.D(n_33),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_3),
.Y(n_95)
);

NAND2x1p5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_4),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_17),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_5),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_100),
.B(n_105),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_106),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_85),
.B(n_7),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_90),
.B(n_7),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_98),
.B1(n_104),
.B2(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_16),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

AOI21x1_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_119),
.B(n_122),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_18),
.C(n_19),
.Y(n_118)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_120),
.C(n_24),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_23),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_117),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_128),
.B(n_129),
.Y(n_130)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_98),
.B1(n_102),
.B2(n_121),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_130),
.A2(n_126),
.B(n_129),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_113),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_132),
.B(n_125),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_96),
.B1(n_112),
.B2(n_103),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_27),
.B(n_30),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_135),
.A2(n_31),
.B(n_32),
.Y(n_136)
);


endmodule