module real_jpeg_11515_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_2),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_81),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_2),
.A2(n_60),
.B1(n_61),
.B2(n_81),
.Y(n_139)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_3),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_4),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_199)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_6),
.A2(n_41),
.B1(n_60),
.B2(n_61),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_47),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_63),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_9),
.A2(n_37),
.B1(n_38),
.B2(n_63),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_12),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_44),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g101 ( 
.A(n_14),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_137),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_101),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_14),
.B(n_61),
.C(n_84),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_14),
.B(n_36),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_14),
.A2(n_64),
.B(n_165),
.Y(n_181)
);

O2A1O1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_14),
.A2(n_27),
.B(n_35),
.C(n_192),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_101),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_15),
.A2(n_44),
.B1(n_45),
.B2(n_49),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_15),
.B(n_28),
.Y(n_74)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_125),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_20),
.B(n_103),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_89),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_21),
.A2(n_22),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_42),
.B2(n_56),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_24),
.B(n_56),
.C(n_57),
.Y(n_122)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_26),
.A2(n_31),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_27),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

AOI32xp33_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_45),
.A3(n_49),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_31),
.A2(n_39),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_32),
.B(n_40),
.Y(n_120)
);

NOR2x1_ASAP7_75t_R g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_34),
.A2(n_37),
.B(n_101),
.Y(n_192)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_37),
.A2(n_38),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_38),
.B(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_48),
.B(n_50),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_43),
.A2(n_48),
.B1(n_52),
.B2(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

O2A1O1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_45),
.A2(n_52),
.B(n_101),
.C(n_102),
.Y(n_100)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_55),
.Y(n_99)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_48),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_71),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_58),
.A2(n_71),
.B1(n_72),
.B2(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_64),
.B1(n_67),
.B2(n_70),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_59),
.A2(n_64),
.B1(n_70),
.B2(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_66),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_61),
.B1(n_84),
.B2(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_60),
.B(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_64),
.A2(n_70),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_64),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_65),
.A2(n_66),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_65),
.B(n_166),
.Y(n_179)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_66),
.B(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_70),
.A2(n_171),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_70),
.B(n_101),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_70),
.A2(n_139),
.B(n_179),
.Y(n_193)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_75),
.B(n_89),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_76),
.B(n_79),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_77),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_87),
.B2(n_88),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_82),
.B(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_87),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_82),
.A2(n_88),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_86),
.A2(n_92),
.B(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_86),
.B(n_101),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_93),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_97),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_90),
.B(n_94),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_95),
.A2(n_96),
.B(n_120),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_96),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_98),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_122),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_114),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_110),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_118),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_143),
.B(n_223),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_140),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_127),
.B(n_140),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_131),
.C(n_133),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_128),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_131),
.B(n_133),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.C(n_138),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_138),
.Y(n_209)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_218),
.B(n_222),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_203),
.B(n_217),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_187),
.B(n_202),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_167),
.B(n_186),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_156),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_148),
.B(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_149),
.A2(n_150),
.B1(n_154),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_152),
.A2(n_153),
.B(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_154),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_164),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_175),
.B(n_185),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_169),
.B(n_173),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_180),
.B(n_184),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_177),
.B(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_188),
.B(n_189),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_197),
.C(n_201),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_191),
.B(n_193),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_194)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_197),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_211),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_213),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_213),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);


endmodule