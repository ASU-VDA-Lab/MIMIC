module fake_ibex_1083_n_1861 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_357, n_88, n_412, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_411, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_1861);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_357;
input n_88;
input n_412;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_411;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_1861;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1566;
wire n_1464;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_532;
wire n_726;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_545;
wire n_887;
wire n_1162;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_423;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_648;
wire n_571;
wire n_1726;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1199;
wire n_1767;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1734;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_980;
wire n_1193;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_414;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_61),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_40),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_255),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_395),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_167),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_339),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_385),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

BUFx2_ASAP7_75t_L g421 ( 
.A(n_44),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_33),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_335),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_405),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_174),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_128),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_293),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_172),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_242),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_325),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_382),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_20),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_376),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_53),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_393),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_143),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_341),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_56),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_51),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_76),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_300),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_136),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_230),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_138),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_4),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_159),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_253),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_355),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_35),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_348),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_1),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_321),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_59),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_43),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_73),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_200),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_50),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_249),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_175),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_3),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_31),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_400),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_72),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_184),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_297),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_152),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_250),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_215),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_239),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_404),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_352),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_153),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_225),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_22),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_319),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_367),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_151),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_72),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_183),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_19),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_38),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_104),
.Y(n_486)
);

INVx1_ASAP7_75t_SL g487 ( 
.A(n_366),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_271),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_269),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_273),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_216),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_410),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_317),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_129),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_165),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_278),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_268),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_399),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_333),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_387),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_259),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_141),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_337),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_166),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_347),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_64),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_42),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_58),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_374),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_284),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_292),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_36),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_189),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_248),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_359),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_177),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_380),
.Y(n_517)
);

BUFx10_ASAP7_75t_L g518 ( 
.A(n_111),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_291),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_63),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_263),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_203),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_306),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_373),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_221),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_294),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_109),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_233),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_160),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_157),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_117),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_115),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_301),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_52),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_349),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_314),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_18),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_244),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_142),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_126),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_191),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_396),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_287),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_381),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_41),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_286),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_70),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_398),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_316),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_322),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_288),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_130),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_375),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_10),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_8),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_298),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_378),
.Y(n_557)
);

CKINVDCx16_ASAP7_75t_R g558 ( 
.A(n_81),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_411),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_358),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_12),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_89),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_320),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_84),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_38),
.Y(n_565)
);

CKINVDCx16_ASAP7_75t_R g566 ( 
.A(n_343),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_401),
.Y(n_567)
);

BUFx10_ASAP7_75t_L g568 ( 
.A(n_304),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_370),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_386),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_251),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_42),
.Y(n_572)
);

BUFx10_ASAP7_75t_L g573 ( 
.A(n_37),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_88),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_2),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_73),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_112),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_16),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_403),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_46),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_407),
.Y(n_581)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_351),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_368),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_149),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_309),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_173),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_83),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_296),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_85),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_39),
.Y(n_590)
);

CKINVDCx11_ASAP7_75t_R g591 ( 
.A(n_155),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_363),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_315),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_364),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_11),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_45),
.Y(n_596)
);

CKINVDCx14_ASAP7_75t_R g597 ( 
.A(n_369),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_150),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_28),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_277),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_360),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_310),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_102),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_390),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_35),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_12),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_50),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_234),
.Y(n_608)
);

INVx1_ASAP7_75t_SL g609 ( 
.A(n_21),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_32),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_389),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_85),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_46),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_388),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_342),
.Y(n_615)
);

BUFx10_ASAP7_75t_L g616 ( 
.A(n_156),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_217),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_187),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_356),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_106),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_340),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_2),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_285),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_379),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_111),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_265),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_270),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_93),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_91),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_357),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_226),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_383),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_39),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_377),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_74),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_312),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_228),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_108),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_402),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_290),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_372),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_26),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_408),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_346),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_98),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_208),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_392),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_76),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_145),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_328),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_170),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_345),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_185),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_17),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_362),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_74),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_354),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_186),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_262),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_45),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_97),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_114),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_119),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_210),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_82),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_302),
.Y(n_666)
);

INVxp67_ASAP7_75t_SL g667 ( 
.A(n_21),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_171),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_240),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_92),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_214),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_43),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_47),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_391),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_394),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_353),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_318),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_326),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_91),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_336),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_54),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_131),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_365),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_344),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_13),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_132),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_23),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_361),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_338),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_14),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_198),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_324),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_60),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_282),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_55),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_413),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_591),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_591),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_421),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_624),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_558),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_677),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_511),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_459),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_518),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_490),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_563),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_459),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_466),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_653),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_537),
.B(n_0),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_577),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_566),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_582),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_577),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_415),
.Y(n_716)
);

CKINVDCx16_ASAP7_75t_R g717 ( 
.A(n_518),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_506),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_506),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_415),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_447),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_540),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_418),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_540),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_681),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_681),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_418),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_453),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_561),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_492),
.Y(n_730)
);

NOR2xp67_ASAP7_75t_L g731 ( 
.A(n_607),
.B(n_0),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_661),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_672),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_674),
.B(n_419),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_561),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_426),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_492),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_523),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_440),
.Y(n_739)
);

CKINVDCx20_ASAP7_75t_R g740 ( 
.A(n_523),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_442),
.Y(n_741)
);

BUFx2_ASAP7_75t_L g742 ( 
.A(n_414),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_451),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_456),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_422),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_524),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_524),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_457),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_557),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_557),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_518),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_600),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_470),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_478),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_482),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_573),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_484),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_600),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_486),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_658),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_658),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_531),
.Y(n_762)
);

INVxp67_ASAP7_75t_SL g763 ( 
.A(n_532),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_554),
.Y(n_764)
);

CKINVDCx20_ASAP7_75t_R g765 ( 
.A(n_686),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_562),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_564),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_575),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_686),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_434),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_599),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_625),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_573),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_633),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_645),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_656),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_687),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_597),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_690),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_568),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_573),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_603),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_417),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_597),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_441),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_455),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_462),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_464),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_467),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_568),
.B(n_1),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_568),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_616),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_485),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_697),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_753),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_699),
.B(n_616),
.Y(n_796)
);

INVx3_ASAP7_75t_L g797 ( 
.A(n_753),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_698),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_703),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_788),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_788),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_712),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_728),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_732),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_715),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_733),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_725),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_751),
.B(n_427),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_704),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_717),
.A2(n_507),
.B1(n_512),
.B2(n_508),
.Y(n_810)
);

AND2x6_ASAP7_75t_L g811 ( 
.A(n_790),
.B(n_416),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_R g812 ( 
.A(n_784),
.B(n_520),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_736),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_739),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_726),
.Y(n_815)
);

NOR2xp67_ASAP7_75t_L g816 ( 
.A(n_756),
.B(n_705),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_741),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_743),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_744),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_716),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_720),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_723),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_748),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_742),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_727),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_754),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_755),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_757),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_759),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_762),
.Y(n_830)
);

CKINVDCx20_ASAP7_75t_R g831 ( 
.A(n_704),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_721),
.B(n_616),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_R g833 ( 
.A(n_784),
.B(n_527),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_780),
.B(n_534),
.Y(n_834)
);

NAND2xp33_ASAP7_75t_SL g835 ( 
.A(n_773),
.B(n_603),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_730),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_764),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_766),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_R g839 ( 
.A(n_709),
.B(n_545),
.Y(n_839)
);

XNOR2xp5_ASAP7_75t_L g840 ( 
.A(n_696),
.B(n_547),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_767),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_768),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_785),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_745),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_737),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_791),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_771),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_738),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_746),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_772),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_770),
.Y(n_851)
);

INVx5_ASAP7_75t_L g852 ( 
.A(n_783),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_747),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_774),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_792),
.B(n_555),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_786),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_750),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_775),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_700),
.B(n_667),
.Y(n_859)
);

OA21x2_ASAP7_75t_L g860 ( 
.A1(n_782),
.A2(n_481),
.B(n_470),
.Y(n_860)
);

CKINVDCx20_ASAP7_75t_R g861 ( 
.A(n_708),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_702),
.B(n_565),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_706),
.B(n_572),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_776),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_752),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_779),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_734),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_758),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_763),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_760),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_777),
.Y(n_871)
);

INVxp67_ASAP7_75t_L g872 ( 
.A(n_711),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_708),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_787),
.Y(n_874)
);

OA21x2_ASAP7_75t_L g875 ( 
.A1(n_731),
.A2(n_494),
.B(n_481),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_707),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_710),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_761),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_783),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_783),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_789),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_778),
.B(n_494),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_769),
.Y(n_883)
);

INVxp67_ASAP7_75t_SL g884 ( 
.A(n_773),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_740),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_740),
.Y(n_886)
);

BUFx2_ASAP7_75t_L g887 ( 
.A(n_793),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_749),
.Y(n_888)
);

CKINVDCx16_ASAP7_75t_R g889 ( 
.A(n_781),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_713),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_749),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_714),
.B(n_574),
.Y(n_892)
);

XOR2xp5_ASAP7_75t_L g893 ( 
.A(n_696),
.B(n_576),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_781),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_701),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_701),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_765),
.B(n_580),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_765),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_718),
.B(n_587),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_719),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_722),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_724),
.Y(n_902)
);

XOR2xp5_ASAP7_75t_L g903 ( 
.A(n_718),
.B(n_589),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_729),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_735),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_735),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_697),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_728),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_780),
.B(n_519),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_753),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_753),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_728),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_697),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_753),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_697),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_699),
.B(n_590),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_753),
.A2(n_592),
.B(n_519),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_753),
.A2(n_593),
.B(n_592),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_697),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_753),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_728),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_697),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_753),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_780),
.B(n_593),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_697),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_728),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_728),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_753),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_780),
.B(n_595),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_753),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_728),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_742),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_699),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_753),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_697),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_697),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_728),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_728),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_753),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_728),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_699),
.B(n_596),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_728),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_697),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_843),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_807),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_917),
.Y(n_947)
);

AND2x6_ASAP7_75t_L g948 ( 
.A(n_880),
.B(n_416),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_827),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_933),
.Y(n_950)
);

NAND3xp33_ASAP7_75t_L g951 ( 
.A(n_872),
.B(n_606),
.C(n_605),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_934),
.B(n_824),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_800),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_934),
.B(n_610),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_887),
.Y(n_955)
);

AND2x6_ASAP7_75t_L g956 ( 
.A(n_880),
.B(n_608),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_879),
.B(n_695),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_801),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_852),
.B(n_423),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_872),
.A2(n_613),
.B1(n_622),
.B2(n_612),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_869),
.A2(n_620),
.B1(n_603),
.B2(n_431),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_824),
.B(n_628),
.Y(n_962)
);

INVx4_ASAP7_75t_L g963 ( 
.A(n_852),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_867),
.B(n_424),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_846),
.B(n_487),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_807),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_867),
.B(n_425),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_803),
.Y(n_968)
);

INVx4_ASAP7_75t_SL g969 ( 
.A(n_811),
.Y(n_969)
);

CKINVDCx16_ASAP7_75t_R g970 ( 
.A(n_889),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_804),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_846),
.B(n_500),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_896),
.B(n_603),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_867),
.B(n_813),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_867),
.B(n_814),
.Y(n_975)
);

AND2x2_ASAP7_75t_SL g976 ( 
.A(n_856),
.B(n_620),
.Y(n_976)
);

HB1xp67_ASAP7_75t_L g977 ( 
.A(n_844),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_871),
.A2(n_635),
.B(n_629),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_876),
.B(n_428),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_844),
.B(n_638),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_806),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_908),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_912),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_807),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_852),
.B(n_430),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_877),
.B(n_432),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_852),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_827),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_921),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_851),
.B(n_642),
.Y(n_990)
);

BUFx3_ASAP7_75t_L g991 ( 
.A(n_794),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_851),
.B(n_648),
.Y(n_992)
);

OR2x2_ASAP7_75t_L g993 ( 
.A(n_916),
.B(n_436),
.Y(n_993)
);

INVx4_ASAP7_75t_SL g994 ( 
.A(n_811),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_927),
.Y(n_995)
);

BUFx10_ASAP7_75t_L g996 ( 
.A(n_798),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_827),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_834),
.B(n_433),
.Y(n_998)
);

BUFx8_ASAP7_75t_SL g999 ( 
.A(n_809),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_808),
.B(n_578),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_928),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_855),
.B(n_435),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_859),
.A2(n_620),
.B1(n_429),
.B2(n_450),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_856),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_907),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_859),
.B(n_437),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_932),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_807),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_874),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_940),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_818),
.B(n_438),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_930),
.B(n_443),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_892),
.B(n_444),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_938),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_939),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_819),
.B(n_445),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_827),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_941),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_838),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_943),
.Y(n_1020)
);

INVx4_ASAP7_75t_SL g1021 ( 
.A(n_811),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_838),
.Y(n_1022)
);

NAND3x1_ASAP7_75t_L g1023 ( 
.A(n_902),
.B(n_458),
.C(n_439),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_838),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_838),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_900),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_847),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_847),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_847),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_837),
.B(n_446),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_816),
.B(n_609),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_841),
.B(n_448),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_842),
.B(n_452),
.Y(n_1033)
);

INVx6_ASAP7_75t_L g1034 ( 
.A(n_847),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_850),
.B(n_454),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_L g1036 ( 
.A(n_811),
.B(n_694),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_901),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_854),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_854),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_854),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_795),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_854),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_858),
.B(n_460),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_795),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_802),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_832),
.B(n_468),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_805),
.Y(n_1047)
);

INVxp67_ASAP7_75t_SL g1048 ( 
.A(n_874),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_881),
.B(n_654),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_815),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_796),
.B(n_469),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_864),
.B(n_471),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_882),
.B(n_472),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_918),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_797),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_940),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_797),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_911),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_882),
.B(n_473),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_942),
.B(n_660),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_799),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_911),
.Y(n_1062)
);

AO21x2_ASAP7_75t_L g1063 ( 
.A1(n_866),
.A2(n_465),
.B(n_461),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_940),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_914),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_862),
.B(n_662),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_881),
.B(n_663),
.Y(n_1067)
);

OAI22xp33_ASAP7_75t_SL g1068 ( 
.A1(n_884),
.A2(n_670),
.B1(n_673),
.B2(n_665),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_863),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_914),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_835),
.A2(n_693),
.B1(n_685),
.B2(n_679),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_920),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_SL g1073 ( 
.A(n_884),
.B(n_475),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_920),
.Y(n_1074)
);

AND2x6_ASAP7_75t_L g1075 ( 
.A(n_890),
.B(n_608),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_940),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_810),
.B(n_620),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_929),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_860),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_929),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_913),
.B(n_476),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_910),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_899),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_923),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_924),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_918),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_931),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_817),
.B(n_480),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_823),
.B(n_488),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_935),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_826),
.B(n_489),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_828),
.B(n_491),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_829),
.B(n_493),
.Y(n_1093)
);

BUFx10_ASAP7_75t_L g1094 ( 
.A(n_915),
.Y(n_1094)
);

INVx4_ASAP7_75t_L g1095 ( 
.A(n_811),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_830),
.B(n_498),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_909),
.B(n_499),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_875),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_875),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_909),
.B(n_623),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_875),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_918),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_925),
.B(n_501),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_812),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_925),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_812),
.Y(n_1106)
);

NAND2xp33_ASAP7_75t_SL g1107 ( 
.A(n_839),
.B(n_833),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_897),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_860),
.Y(n_1109)
);

OAI221xp5_ASAP7_75t_L g1110 ( 
.A1(n_835),
.A2(n_479),
.B1(n_483),
.B2(n_477),
.C(n_474),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_839),
.B(n_623),
.Y(n_1111)
);

INVx3_ASAP7_75t_L g1112 ( 
.A(n_860),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_896),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_833),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_894),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_895),
.B(n_502),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_896),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_896),
.A2(n_496),
.B1(n_497),
.B2(n_495),
.Y(n_1118)
);

NAND2xp33_ASAP7_75t_L g1119 ( 
.A(n_944),
.B(n_692),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_919),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_922),
.B(n_509),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_926),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_936),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_820),
.B(n_513),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_906),
.B(n_904),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_821),
.Y(n_1126)
);

AO22x2_ASAP7_75t_L g1127 ( 
.A1(n_903),
.A2(n_504),
.B1(n_505),
.B2(n_503),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_937),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_822),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_898),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_898),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_825),
.B(n_515),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_836),
.B(n_640),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_898),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_893),
.B(n_3),
.Y(n_1135)
);

INVx4_ASAP7_75t_SL g1136 ( 
.A(n_898),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_845),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_848),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_849),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_853),
.A2(n_526),
.B1(n_530),
.B2(n_514),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_857),
.B(n_516),
.Y(n_1141)
);

BUFx8_ASAP7_75t_SL g1142 ( 
.A(n_831),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_865),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_905),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_868),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_870),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_878),
.Y(n_1147)
);

NAND3x1_ASAP7_75t_L g1148 ( 
.A(n_840),
.B(n_548),
.C(n_542),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_883),
.B(n_640),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_861),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_904),
.Y(n_1151)
);

NAND2xp33_ASAP7_75t_L g1152 ( 
.A(n_885),
.B(n_517),
.Y(n_1152)
);

AND2x6_ASAP7_75t_L g1153 ( 
.A(n_886),
.B(n_643),
.Y(n_1153)
);

AND2x6_ASAP7_75t_L g1154 ( 
.A(n_891),
.B(n_643),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_888),
.B(n_550),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_873),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_872),
.B(n_521),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_803),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_803),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_917),
.Y(n_1160)
);

INVxp33_ASAP7_75t_L g1161 ( 
.A(n_934),
.Y(n_1161)
);

OR2x2_ASAP7_75t_L g1162 ( 
.A(n_934),
.B(n_4),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_952),
.B(n_5),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_974),
.B(n_522),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_975),
.B(n_525),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1161),
.B(n_528),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1083),
.A2(n_570),
.B(n_584),
.C(n_551),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_968),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_971),
.B(n_981),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_982),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_983),
.B(n_529),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_989),
.B(n_533),
.Y(n_1172)
);

AND2x6_ASAP7_75t_SL g1173 ( 
.A(n_999),
.B(n_585),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_977),
.B(n_535),
.Y(n_1174)
);

AOI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1105),
.A2(n_604),
.B1(n_611),
.B2(n_602),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_947),
.A2(n_636),
.B(n_631),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_950),
.B(n_1069),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_995),
.B(n_536),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_993),
.B(n_538),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1001),
.B(n_539),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1007),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1009),
.B(n_5),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1014),
.B(n_541),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_945),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1015),
.B(n_543),
.Y(n_1185)
);

INVxp33_ASAP7_75t_L g1186 ( 
.A(n_1004),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1041),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_955),
.B(n_6),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1018),
.A2(n_644),
.B1(n_646),
.B2(n_641),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_980),
.B(n_6),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1049),
.B(n_544),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_990),
.B(n_7),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1020),
.B(n_546),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1073),
.B(n_549),
.Y(n_1194)
);

A2O1A1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1158),
.A2(n_650),
.B(n_651),
.C(n_649),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_992),
.B(n_7),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_SL g1197 ( 
.A(n_1095),
.B(n_691),
.Y(n_1197)
);

AO22x1_ASAP7_75t_L g1198 ( 
.A1(n_1061),
.A2(n_553),
.B1(n_556),
.B2(n_552),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1159),
.B(n_559),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1045),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1041),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1098),
.A2(n_659),
.B(n_666),
.C(n_655),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_991),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1095),
.B(n_976),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_947),
.A2(n_682),
.B(n_671),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1157),
.B(n_560),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1077),
.A2(n_569),
.B1(n_571),
.B2(n_567),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_L g1208 ( 
.A(n_948),
.B(n_579),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1144),
.Y(n_1209)
);

INVx5_ASAP7_75t_L g1210 ( 
.A(n_973),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1160),
.A2(n_583),
.B(n_581),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_962),
.B(n_586),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1047),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1003),
.B(n_588),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_963),
.B(n_598),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1063),
.A2(n_689),
.B1(n_614),
.B2(n_615),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_963),
.B(n_601),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_965),
.B(n_617),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1054),
.A2(n_619),
.B(n_618),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1048),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1050),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1055),
.Y(n_1222)
);

NAND2x1p5_ASAP7_75t_L g1223 ( 
.A(n_1005),
.B(n_420),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_972),
.B(n_621),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1100),
.B(n_626),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1100),
.B(n_627),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_996),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1144),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_SL g1229 ( 
.A(n_1126),
.B(n_630),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_987),
.Y(n_1230)
);

NOR2xp33_ASAP7_75t_L g1231 ( 
.A(n_1060),
.B(n_632),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1057),
.Y(n_1232)
);

AOI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_688),
.B1(n_637),
.B2(n_639),
.Y(n_1233)
);

O2A1O1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1068),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_987),
.B(n_634),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1066),
.B(n_647),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1101),
.A2(n_664),
.B1(n_668),
.B2(n_657),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1044),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1101),
.A2(n_675),
.B1(n_676),
.B2(n_669),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1160),
.A2(n_680),
.B(n_678),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1044),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1111),
.B(n_683),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1046),
.B(n_684),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1053),
.B(n_9),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1115),
.A2(n_449),
.B1(n_463),
.B2(n_420),
.Y(n_1245)
);

INVx3_ASAP7_75t_L g1246 ( 
.A(n_973),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1054),
.A2(n_449),
.B1(n_463),
.B2(n_420),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1067),
.B(n_420),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_996),
.Y(n_1249)
);

BUFx5_ASAP7_75t_L g1250 ( 
.A(n_1086),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1058),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_969),
.B(n_11),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1085),
.Y(n_1253)
);

NAND2x1p5_ASAP7_75t_L g1254 ( 
.A(n_1104),
.B(n_449),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1059),
.B(n_13),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1090),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_954),
.B(n_14),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1144),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1051),
.B(n_15),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_966),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1162),
.B(n_15),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_957),
.B(n_16),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1062),
.Y(n_1263)
);

INVxp67_ASAP7_75t_L g1264 ( 
.A(n_1142),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_957),
.B(n_17),
.Y(n_1265)
);

INVx3_ASAP7_75t_L g1266 ( 
.A(n_1131),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1079),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_960),
.B(n_18),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1065),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1000),
.B(n_19),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1081),
.B(n_449),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_SL g1272 ( 
.A(n_1128),
.B(n_463),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_966),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1082),
.A2(n_1084),
.B1(n_1087),
.B2(n_1109),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1036),
.A2(n_510),
.B1(n_594),
.B2(n_463),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_970),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1000),
.B(n_20),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1086),
.A2(n_594),
.B1(n_652),
.B2(n_510),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1094),
.B(n_22),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1070),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1103),
.B(n_23),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_SL g1282 ( 
.A(n_1026),
.B(n_24),
.C(n_25),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1072),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1099),
.A2(n_594),
.B1(n_652),
.B2(n_510),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1074),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_998),
.B(n_24),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1002),
.B(n_25),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1094),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1012),
.B(n_26),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_979),
.B(n_27),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1112),
.A2(n_594),
.B(n_510),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_986),
.B(n_27),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1078),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1013),
.B(n_28),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1151),
.B(n_29),
.Y(n_1295)
);

NOR2xp33_ASAP7_75t_R g1296 ( 
.A(n_1107),
.B(n_29),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1080),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1112),
.A2(n_652),
.B(n_134),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1099),
.A2(n_652),
.B1(n_32),
.B2(n_30),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1106),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1127),
.A2(n_33),
.B1(n_30),
.B2(n_31),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_964),
.B(n_34),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1127),
.B(n_34),
.Y(n_1303)
);

NOR3xp33_ASAP7_75t_L g1304 ( 
.A(n_1156),
.B(n_36),
.C(n_37),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_967),
.B(n_40),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1130),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1102),
.A2(n_1016),
.B(n_1011),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1030),
.B(n_41),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_966),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1033),
.B(n_44),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1035),
.B(n_47),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1079),
.A2(n_51),
.B1(n_48),
.B2(n_49),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1110),
.A2(n_1134),
.B1(n_1079),
.B2(n_978),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1135),
.A2(n_52),
.B1(n_48),
.B2(n_49),
.Y(n_1314)
);

AND2x4_ASAP7_75t_SL g1315 ( 
.A(n_1156),
.B(n_53),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1052),
.B(n_54),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1102),
.A2(n_135),
.B(n_133),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_969),
.B(n_55),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_984),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_984),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_984),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1117),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_948),
.B(n_956),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1131),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1113),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1136),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_948),
.B(n_56),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1114),
.B(n_57),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1136),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_951),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_948),
.B(n_60),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_SL g1332 ( 
.A1(n_1116),
.A2(n_139),
.B(n_140),
.C(n_137),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1149),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_SL g1334 ( 
.A(n_1037),
.B(n_61),
.C(n_62),
.Y(n_1334)
);

INVxp67_ASAP7_75t_L g1335 ( 
.A(n_1133),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_956),
.B(n_62),
.Y(n_1336)
);

XOR2xp5_ASAP7_75t_L g1337 ( 
.A(n_1150),
.B(n_953),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_994),
.B(n_1021),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1008),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1008),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1006),
.B(n_63),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_949),
.A2(n_146),
.B(n_144),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_956),
.B(n_64),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1088),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_956),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_961),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1149),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1023),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1097),
.A2(n_71),
.B1(n_68),
.B2(n_69),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1155),
.B(n_71),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1031),
.B(n_75),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_949),
.A2(n_148),
.B(n_147),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1089),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1031),
.B(n_75),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_SL g1355 ( 
.A1(n_1155),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_SL g1356 ( 
.A(n_994),
.B(n_77),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1168),
.B(n_1118),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_SL g1358 ( 
.A(n_1210),
.B(n_1146),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1250),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1210),
.B(n_1147),
.Y(n_1360)
);

BUFx8_ASAP7_75t_L g1361 ( 
.A(n_1249),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1250),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1227),
.B(n_1021),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1184),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1170),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1181),
.B(n_1125),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1169),
.B(n_1140),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1250),
.Y(n_1368)
);

NOR2x1p5_ASAP7_75t_L g1369 ( 
.A(n_1203),
.B(n_958),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1344),
.B(n_1120),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1176),
.A2(n_1071),
.B(n_1092),
.C(n_1091),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1210),
.B(n_1129),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1229),
.B(n_1137),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1230),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1250),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1250),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1276),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1186),
.B(n_1138),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1335),
.B(n_1139),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1220),
.Y(n_1380)
);

BUFx3_ASAP7_75t_L g1381 ( 
.A(n_1288),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1253),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1353),
.B(n_1153),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_L g1384 ( 
.A(n_1264),
.B(n_1122),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1337),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1256),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1267),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1163),
.B(n_1153),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1200),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1213),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1221),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1333),
.B(n_1347),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1222),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1274),
.B(n_1153),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_SL g1395 ( 
.A(n_1314),
.B(n_1123),
.C(n_1121),
.Y(n_1395)
);

AOI21xp33_ASAP7_75t_L g1396 ( 
.A1(n_1244),
.A2(n_1028),
.B(n_1025),
.Y(n_1396)
);

INVxp67_ASAP7_75t_SL g1397 ( 
.A(n_1267),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1315),
.Y(n_1398)
);

OR2x6_ASAP7_75t_L g1399 ( 
.A(n_1252),
.B(n_1143),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_SL g1400 ( 
.A(n_1252),
.B(n_1153),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1230),
.Y(n_1401)
);

BUFx4f_ASAP7_75t_L g1402 ( 
.A(n_1303),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1232),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1188),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1182),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1251),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1177),
.A2(n_1145),
.B1(n_1148),
.B2(n_1152),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1262),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1179),
.B(n_1350),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1263),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1269),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1280),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1267),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1283),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1300),
.B(n_1124),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1285),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1293),
.Y(n_1417)
);

INVx3_ASAP7_75t_L g1418 ( 
.A(n_1246),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1297),
.Y(n_1419)
);

NAND3xp33_ASAP7_75t_SL g1420 ( 
.A(n_1301),
.B(n_1141),
.C(n_1132),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1322),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1306),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1187),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1201),
.Y(n_1424)
);

NOR3xp33_ASAP7_75t_SL g1425 ( 
.A(n_1282),
.B(n_1043),
.C(n_1032),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1274),
.B(n_1154),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1265),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_SL g1429 ( 
.A(n_1272),
.B(n_1154),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1246),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1196),
.A2(n_1154),
.B1(n_1075),
.B2(n_1119),
.Y(n_1431)
);

INVx4_ASAP7_75t_L g1432 ( 
.A(n_1223),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_1231),
.B(n_1212),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1270),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1238),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1277),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1268),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1257),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1174),
.A2(n_1154),
.B1(n_1075),
.B2(n_1093),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1236),
.B(n_1096),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1166),
.B(n_959),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_SL g1442 ( 
.A(n_1296),
.B(n_985),
.Y(n_1442)
);

AOI221xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1202),
.A2(n_1038),
.B1(n_1029),
.B2(n_1039),
.C(n_1042),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1351),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1354),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1279),
.B(n_1261),
.Y(n_1446)
);

INVx2_ASAP7_75t_SL g1447 ( 
.A(n_1209),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1175),
.B(n_1075),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1241),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1175),
.B(n_1075),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1327),
.Y(n_1451)
);

INVx1_ASAP7_75t_SL g1452 ( 
.A(n_1331),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1326),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1295),
.A2(n_946),
.B1(n_1034),
.B2(n_997),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1266),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1301),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1254),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1233),
.B(n_1198),
.Y(n_1458)
);

AND2x6_ASAP7_75t_SL g1459 ( 
.A(n_1173),
.B(n_78),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_R g1460 ( 
.A(n_1271),
.B(n_1208),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_R g1461 ( 
.A(n_1334),
.B(n_946),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1266),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1228),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1325),
.Y(n_1464)
);

O2A1O1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1195),
.A2(n_1017),
.B(n_1019),
.C(n_988),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1307),
.B(n_1022),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1324),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1189),
.B(n_1024),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1349),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1233),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1258),
.B(n_1329),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1336),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_1355),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1237),
.B(n_1008),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1239),
.B(n_1010),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1308),
.Y(n_1476)
);

AOI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1291),
.A2(n_1040),
.B(n_1027),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1260),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1189),
.B(n_1056),
.Y(n_1479)
);

NOR2xp33_ASAP7_75t_L g1480 ( 
.A(n_1167),
.B(n_1034),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1345),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1328),
.Y(n_1482)
);

BUFx12f_ASAP7_75t_SL g1483 ( 
.A(n_1348),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1205),
.B(n_1076),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1310),
.Y(n_1485)
);

AND2x4_ASAP7_75t_L g1486 ( 
.A(n_1215),
.B(n_1010),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_SL g1487 ( 
.A(n_1207),
.B(n_1010),
.Y(n_1487)
);

CKINVDCx8_ASAP7_75t_R g1488 ( 
.A(n_1341),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1311),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1273),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1309),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1345),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1343),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_L g1494 ( 
.A(n_1225),
.B(n_1064),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1216),
.B(n_1064),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1216),
.B(n_1064),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1380),
.B(n_1348),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1466),
.A2(n_1298),
.B(n_1317),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1390),
.Y(n_1499)
);

INVx3_ASAP7_75t_SL g1500 ( 
.A(n_1377),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1466),
.A2(n_1255),
.B(n_1281),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1477),
.A2(n_1342),
.B(n_1284),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1481),
.A2(n_1299),
.B1(n_1284),
.B2(n_1346),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1484),
.A2(n_1287),
.B(n_1286),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1359),
.A2(n_1320),
.B(n_1319),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1469),
.A2(n_1299),
.B(n_1313),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1362),
.A2(n_1339),
.B(n_1321),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1365),
.Y(n_1508)
);

INVxp67_ASAP7_75t_SL g1509 ( 
.A(n_1400),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1484),
.A2(n_1289),
.B(n_1294),
.Y(n_1510)
);

AOI221x1_ASAP7_75t_L g1511 ( 
.A1(n_1420),
.A2(n_1304),
.B1(n_1312),
.B2(n_1278),
.C(n_1247),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1361),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1402),
.B(n_1204),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1371),
.A2(n_1259),
.B(n_1332),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1437),
.A2(n_1316),
.B(n_1275),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1456),
.B(n_1290),
.Y(n_1516)
);

AOI221xp5_ASAP7_75t_SL g1517 ( 
.A1(n_1433),
.A2(n_1234),
.B1(n_1292),
.B2(n_1248),
.C(n_1302),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1393),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1367),
.B(n_1226),
.Y(n_1519)
);

AOI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1394),
.A2(n_1219),
.B(n_1305),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1361),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1367),
.B(n_1171),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1368),
.A2(n_1340),
.B(n_1352),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1443),
.A2(n_1245),
.B(n_1275),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1375),
.A2(n_1323),
.B(n_1338),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1366),
.B(n_1370),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1432),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1366),
.B(n_1370),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_SL g1529 ( 
.A1(n_1394),
.A2(n_1346),
.B(n_1245),
.Y(n_1529)
);

A2O1A1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1476),
.A2(n_1240),
.B(n_1211),
.C(n_1330),
.Y(n_1530)
);

NOR2xp67_ASAP7_75t_L g1531 ( 
.A(n_1432),
.B(n_1191),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1389),
.B(n_1172),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1399),
.B(n_1318),
.Y(n_1533)
);

OAI21xp5_ASAP7_75t_L g1534 ( 
.A1(n_1427),
.A2(n_1219),
.B(n_1356),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1492),
.A2(n_1194),
.B1(n_1180),
.B2(n_1183),
.Y(n_1535)
);

O2A1O1Ixp5_ASAP7_75t_SL g1536 ( 
.A1(n_1453),
.A2(n_1217),
.B(n_1235),
.C(n_1242),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1402),
.B(n_1178),
.Y(n_1537)
);

BUFx3_ASAP7_75t_L g1538 ( 
.A(n_1364),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1409),
.B(n_1185),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1427),
.A2(n_1165),
.B(n_1164),
.Y(n_1540)
);

AO21x2_ASAP7_75t_L g1541 ( 
.A1(n_1426),
.A2(n_1199),
.B(n_1193),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1399),
.A2(n_1224),
.B1(n_1218),
.B2(n_1243),
.Y(n_1542)
);

AOI21xp5_ASAP7_75t_L g1543 ( 
.A1(n_1485),
.A2(n_1206),
.B(n_1197),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1425),
.B(n_1214),
.C(n_79),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_R g1545 ( 
.A(n_1385),
.B(n_80),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1400),
.B(n_80),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1391),
.B(n_81),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1489),
.A2(n_1475),
.B(n_1474),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1383),
.A2(n_1396),
.B(n_1426),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1399),
.Y(n_1550)
);

A2O1A1Ixp33_ASAP7_75t_L g1551 ( 
.A1(n_1438),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1429),
.B(n_86),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1376),
.A2(n_158),
.B(n_154),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1428),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_1554)
);

AOI21xp5_ASAP7_75t_L g1555 ( 
.A1(n_1383),
.A2(n_162),
.B(n_161),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1404),
.B(n_87),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1473),
.B(n_89),
.Y(n_1557)
);

OAI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1495),
.A2(n_90),
.B(n_92),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1495),
.A2(n_90),
.B(n_93),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1397),
.A2(n_164),
.B(n_163),
.Y(n_1560)
);

O2A1O1Ixp5_ASAP7_75t_L g1561 ( 
.A1(n_1487),
.A2(n_272),
.B(n_412),
.C(n_409),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1417),
.B(n_94),
.Y(n_1562)
);

NAND2x1_ASAP7_75t_L g1563 ( 
.A(n_1387),
.B(n_168),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1470),
.B(n_94),
.Y(n_1564)
);

A2O1A1Ixp33_ASAP7_75t_L g1565 ( 
.A1(n_1480),
.A2(n_95),
.B(n_96),
.C(n_97),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1496),
.A2(n_176),
.B(n_169),
.Y(n_1566)
);

AO21x2_ASAP7_75t_L g1567 ( 
.A1(n_1496),
.A2(n_179),
.B(n_178),
.Y(n_1567)
);

OAI22x1_ASAP7_75t_L g1568 ( 
.A1(n_1369),
.A2(n_1458),
.B1(n_1407),
.B2(n_1483),
.Y(n_1568)
);

A2O1A1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1434),
.A2(n_95),
.B(n_96),
.C(n_98),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1465),
.A2(n_181),
.B(n_180),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1429),
.B(n_99),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1403),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1406),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1381),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1395),
.B(n_99),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1453),
.A2(n_1490),
.B(n_1478),
.Y(n_1576)
);

OAI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1479),
.A2(n_100),
.B(n_101),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1410),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_SL g1579 ( 
.A(n_1457),
.B(n_100),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1576),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1498),
.A2(n_1388),
.B(n_1448),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1508),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1509),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1502),
.A2(n_1388),
.B(n_1448),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1549),
.A2(n_1450),
.B(n_1479),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1526),
.B(n_1379),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1566),
.A2(n_1450),
.B(n_1401),
.Y(n_1587)
);

BUFx2_ASAP7_75t_SL g1588 ( 
.A(n_1512),
.Y(n_1588)
);

OA21x2_ASAP7_75t_L g1589 ( 
.A1(n_1514),
.A2(n_1443),
.B(n_1396),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1523),
.A2(n_1401),
.B(n_1374),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1528),
.B(n_1419),
.Y(n_1591)
);

OAI21x1_ASAP7_75t_L g1592 ( 
.A1(n_1570),
.A2(n_1507),
.B(n_1505),
.Y(n_1592)
);

OAI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1568),
.A2(n_1398),
.B1(n_1482),
.B2(n_1405),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_SL g1594 ( 
.A1(n_1529),
.A2(n_1431),
.B(n_1439),
.Y(n_1594)
);

AOI221xp5_ASAP7_75t_L g1595 ( 
.A1(n_1542),
.A2(n_1408),
.B1(n_1539),
.B2(n_1519),
.C(n_1535),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1501),
.A2(n_1510),
.B(n_1504),
.Y(n_1596)
);

OA21x2_ASAP7_75t_L g1597 ( 
.A1(n_1506),
.A2(n_1468),
.B(n_1444),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1553),
.A2(n_1374),
.B(n_1455),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1499),
.Y(n_1599)
);

OAI21x1_ASAP7_75t_L g1600 ( 
.A1(n_1525),
.A2(n_1462),
.B(n_1468),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1503),
.A2(n_1446),
.B1(n_1488),
.B2(n_1493),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1560),
.A2(n_1421),
.B(n_1418),
.Y(n_1603)
);

OR2x6_ASAP7_75t_L g1604 ( 
.A(n_1533),
.B(n_1387),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1550),
.Y(n_1605)
);

OAI21x1_ASAP7_75t_L g1606 ( 
.A1(n_1520),
.A2(n_1418),
.B(n_1494),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1497),
.A2(n_1503),
.B1(n_1542),
.B2(n_1535),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1578),
.Y(n_1608)
);

BUFx6f_ASAP7_75t_L g1609 ( 
.A(n_1563),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1538),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1506),
.A2(n_1445),
.B(n_1436),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1522),
.B(n_1378),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1558),
.A2(n_1357),
.B(n_1461),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1548),
.A2(n_1467),
.B(n_1422),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1561),
.A2(n_1372),
.B(n_1360),
.Y(n_1615)
);

OAI21x1_ASAP7_75t_L g1616 ( 
.A1(n_1555),
.A2(n_1358),
.B(n_1454),
.Y(n_1616)
);

NAND2x1p5_ASAP7_75t_L g1617 ( 
.A(n_1527),
.B(n_1387),
.Y(n_1617)
);

NAND2x1p5_ASAP7_75t_L g1618 ( 
.A(n_1527),
.B(n_1413),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1518),
.Y(n_1619)
);

OA21x2_ASAP7_75t_L g1620 ( 
.A1(n_1534),
.A2(n_1452),
.B(n_1451),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1530),
.A2(n_1415),
.B(n_1441),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1607),
.B(n_1573),
.Y(n_1622)
);

BUFx8_ASAP7_75t_SL g1623 ( 
.A(n_1605),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1591),
.B(n_1556),
.Y(n_1624)
);

OAI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1595),
.A2(n_1557),
.B1(n_1544),
.B2(n_1564),
.C(n_1575),
.Y(n_1625)
);

OR2x6_ASAP7_75t_L g1626 ( 
.A(n_1604),
.B(n_1533),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1596),
.A2(n_1559),
.B(n_1558),
.Y(n_1627)
);

NAND2xp33_ASAP7_75t_R g1628 ( 
.A(n_1583),
.B(n_1524),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1602),
.A2(n_1516),
.B1(n_1522),
.B2(n_1533),
.Y(n_1629)
);

INVx8_ASAP7_75t_L g1630 ( 
.A(n_1604),
.Y(n_1630)
);

OAI22xp33_ASAP7_75t_L g1631 ( 
.A1(n_1586),
.A2(n_1577),
.B1(n_1559),
.B2(n_1516),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1599),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1621),
.A2(n_1577),
.B1(n_1540),
.B2(n_1579),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1591),
.B(n_1574),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1588),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1582),
.Y(n_1636)
);

OAI22xp5_ASAP7_75t_L g1637 ( 
.A1(n_1593),
.A2(n_1565),
.B1(n_1551),
.B2(n_1554),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1601),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1610),
.B(n_1608),
.Y(n_1639)
);

AOI222xp33_ASAP7_75t_L g1640 ( 
.A1(n_1612),
.A2(n_1545),
.B1(n_1521),
.B2(n_1532),
.C1(n_1537),
.C2(n_1513),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1594),
.A2(n_1524),
.B(n_1515),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1583),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1605),
.B(n_1532),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1604),
.A2(n_1569),
.B1(n_1562),
.B2(n_1547),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1599),
.Y(n_1645)
);

AOI221xp5_ASAP7_75t_L g1646 ( 
.A1(n_1594),
.A2(n_1562),
.B1(n_1547),
.B2(n_1392),
.C(n_1540),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1613),
.A2(n_1541),
.B1(n_1515),
.B2(n_1546),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1604),
.B(n_1531),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1613),
.A2(n_1541),
.B1(n_1534),
.B2(n_1552),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1619),
.Y(n_1650)
);

AND2x4_ASAP7_75t_SL g1651 ( 
.A(n_1619),
.B(n_1363),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1614),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1611),
.B(n_1471),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1634),
.B(n_1624),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1629),
.A2(n_1611),
.B1(n_1613),
.B2(n_1597),
.Y(n_1655)
);

OAI211xp5_ASAP7_75t_L g1656 ( 
.A1(n_1640),
.A2(n_1373),
.B(n_1384),
.C(n_1442),
.Y(n_1656)
);

CKINVDCx14_ASAP7_75t_R g1657 ( 
.A(n_1635),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1629),
.A2(n_1611),
.B1(n_1597),
.B2(n_1571),
.Y(n_1658)
);

OAI211xp5_ASAP7_75t_L g1659 ( 
.A1(n_1633),
.A2(n_1517),
.B(n_1463),
.C(n_1447),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1625),
.A2(n_1597),
.B1(n_1588),
.B2(n_1452),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1626),
.A2(n_1500),
.B1(n_1459),
.B2(n_1617),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1639),
.B(n_1617),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1643),
.B(n_1620),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1636),
.Y(n_1664)
);

OAI22xp33_ASAP7_75t_SL g1665 ( 
.A1(n_1626),
.A2(n_1617),
.B1(n_1618),
.B2(n_1430),
.Y(n_1665)
);

AOI221xp5_ASAP7_75t_L g1666 ( 
.A1(n_1643),
.A2(n_1543),
.B1(n_1471),
.B2(n_1411),
.C(n_1416),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1638),
.Y(n_1667)
);

INVx4_ASAP7_75t_SL g1668 ( 
.A(n_1626),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1630),
.B(n_1642),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1631),
.A2(n_1567),
.B(n_1603),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1633),
.A2(n_1451),
.B1(n_1472),
.B2(n_1620),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1631),
.A2(n_1567),
.B(n_1603),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1645),
.Y(n_1674)
);

OAI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1630),
.A2(n_1618),
.B1(n_1511),
.B2(n_1472),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1646),
.A2(n_1620),
.B1(n_1584),
.B2(n_1589),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1630),
.A2(n_1357),
.B1(n_1609),
.B2(n_1580),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1637),
.A2(n_1414),
.B1(n_1412),
.B2(n_1440),
.C(n_1464),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

OAI221xp5_ASAP7_75t_L g1680 ( 
.A1(n_1647),
.A2(n_1449),
.B1(n_1435),
.B2(n_1423),
.C(n_1424),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1674),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1668),
.B(n_1653),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1664),
.B(n_1667),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1669),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1654),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1663),
.B(n_1653),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1679),
.Y(n_1687)
);

OAI31xp33_ASAP7_75t_L g1688 ( 
.A1(n_1656),
.A2(n_1651),
.A3(n_1644),
.B(n_1648),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1668),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1662),
.B(n_1622),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1669),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1678),
.A2(n_1627),
.B1(n_1623),
.B2(n_1648),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1668),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1669),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1655),
.B(n_1652),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1676),
.B(n_1632),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1677),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1657),
.Y(n_1699)
);

OAI221xp5_ASAP7_75t_SL g1700 ( 
.A1(n_1678),
.A2(n_1660),
.B1(n_1659),
.B2(n_1658),
.C(n_1666),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1680),
.Y(n_1701)
);

OAI211xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1671),
.A2(n_1647),
.B(n_1649),
.C(n_1641),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1670),
.B(n_1627),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1685),
.B(n_1690),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1701),
.A2(n_1661),
.B1(n_1675),
.B2(n_1680),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1692),
.B(n_1585),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1683),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1699),
.Y(n_1708)
);

INVx2_ASAP7_75t_SL g1709 ( 
.A(n_1699),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1686),
.B(n_1649),
.Y(n_1710)
);

NAND4xp25_ASAP7_75t_L g1711 ( 
.A(n_1693),
.B(n_1672),
.C(n_1628),
.D(n_1363),
.Y(n_1711)
);

OAI31xp33_ASAP7_75t_L g1712 ( 
.A1(n_1700),
.A2(n_1665),
.A3(n_1651),
.B(n_1486),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1701),
.A2(n_1589),
.B1(n_1585),
.B2(n_1614),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1692),
.B(n_1580),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1702),
.A2(n_1589),
.B1(n_1606),
.B2(n_1616),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1681),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1688),
.A2(n_1606),
.B1(n_1616),
.B2(n_1615),
.Y(n_1717)
);

OAI33xp33_ASAP7_75t_L g1718 ( 
.A1(n_1698),
.A2(n_101),
.A3(n_102),
.B1(n_103),
.B2(n_104),
.B3(n_105),
.Y(n_1718)
);

NOR4xp25_ASAP7_75t_SL g1719 ( 
.A(n_1707),
.B(n_1684),
.C(n_1689),
.D(n_1695),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1716),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1710),
.B(n_1684),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1706),
.B(n_1689),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1704),
.B(n_1686),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1705),
.B(n_1681),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1708),
.B(n_1695),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1714),
.B(n_1692),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1709),
.Y(n_1727)
);

NAND2x1p5_ASAP7_75t_L g1728 ( 
.A(n_1718),
.B(n_1691),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1712),
.Y(n_1730)
);

BUFx2_ASAP7_75t_L g1731 ( 
.A(n_1705),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1713),
.B(n_1696),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1713),
.B(n_1687),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1715),
.B(n_1687),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1721),
.B(n_1694),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_SL g1736 ( 
.A1(n_1731),
.A2(n_1691),
.B1(n_1694),
.B2(n_1703),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1722),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1694),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1728),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1730),
.B(n_1717),
.C(n_1715),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1730),
.A2(n_1729),
.B1(n_1724),
.B2(n_1732),
.C(n_1721),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1739),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1735),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_1738),
.Y(n_1744)
);

AND2x2_ASAP7_75t_SL g1745 ( 
.A(n_1741),
.B(n_1730),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1745),
.A2(n_1730),
.B1(n_1740),
.B2(n_1736),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1743),
.B(n_1732),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1747),
.B(n_1742),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1746),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1747),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1747),
.B(n_1740),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_L g1752 ( 
.A(n_1749),
.B(n_1744),
.Y(n_1752)
);

NOR3xp33_ASAP7_75t_SL g1753 ( 
.A(n_1750),
.B(n_1745),
.C(n_1734),
.Y(n_1753)
);

XOR2xp5_ASAP7_75t_L g1754 ( 
.A(n_1751),
.B(n_1728),
.Y(n_1754)
);

OAI211xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1748),
.A2(n_1717),
.B(n_1727),
.C(n_1737),
.Y(n_1755)
);

CKINVDCx20_ASAP7_75t_L g1756 ( 
.A(n_1748),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1748),
.Y(n_1757)
);

HB1xp67_ASAP7_75t_L g1758 ( 
.A(n_1748),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1754),
.A2(n_1727),
.B1(n_1719),
.B2(n_1725),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1752),
.B(n_1725),
.C(n_1733),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1756),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1758),
.Y(n_1762)
);

NOR4xp25_ASAP7_75t_L g1763 ( 
.A(n_1757),
.B(n_1723),
.C(n_1720),
.D(n_1386),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1755),
.A2(n_1725),
.B(n_1723),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1753),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1758),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1752),
.A2(n_1691),
.B1(n_1698),
.B2(n_1703),
.C(n_1726),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1758),
.B(n_1722),
.Y(n_1768)
);

AOI211xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1758),
.A2(n_1722),
.B(n_1682),
.C(n_106),
.Y(n_1769)
);

OAI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1691),
.B1(n_1628),
.B2(n_1682),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1761),
.A2(n_1691),
.B1(n_1682),
.B2(n_1697),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1765),
.B(n_1687),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1762),
.Y(n_1773)
);

AOI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1760),
.A2(n_1691),
.B1(n_1682),
.B2(n_1696),
.Y(n_1774)
);

OAI211xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1766),
.A2(n_1767),
.B(n_1759),
.C(n_1768),
.Y(n_1775)
);

AOI311xp33_ASAP7_75t_L g1776 ( 
.A1(n_1764),
.A2(n_103),
.A3(n_105),
.B(n_107),
.C(n_108),
.Y(n_1776)
);

NAND4xp75_ASAP7_75t_L g1777 ( 
.A(n_1763),
.B(n_107),
.C(n_109),
.D(n_110),
.Y(n_1777)
);

NAND4xp75_ASAP7_75t_L g1778 ( 
.A(n_1763),
.B(n_110),
.C(n_112),
.D(n_113),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_R g1779 ( 
.A(n_1761),
.B(n_113),
.Y(n_1779)
);

AOI222xp33_ASAP7_75t_L g1780 ( 
.A1(n_1762),
.A2(n_1697),
.B1(n_1486),
.B2(n_1382),
.C1(n_1609),
.C2(n_1615),
.Y(n_1780)
);

AOI211x1_ASAP7_75t_SL g1781 ( 
.A1(n_1761),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_1781)
);

AOI321xp33_ASAP7_75t_L g1782 ( 
.A1(n_1761),
.A2(n_1697),
.A3(n_117),
.B1(n_118),
.B2(n_119),
.C(n_120),
.Y(n_1782)
);

NAND3xp33_ASAP7_75t_SL g1783 ( 
.A(n_1761),
.B(n_1460),
.C(n_1536),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1769),
.A2(n_1609),
.B1(n_118),
.B2(n_120),
.C(n_121),
.Y(n_1784)
);

AOI21xp33_ASAP7_75t_L g1785 ( 
.A1(n_1773),
.A2(n_116),
.B(n_121),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1784),
.A2(n_122),
.B(n_123),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1781),
.A2(n_1697),
.B1(n_1609),
.B2(n_124),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1779),
.Y(n_1788)
);

XOR2xp5_ASAP7_75t_L g1789 ( 
.A(n_1777),
.B(n_122),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1770),
.B(n_123),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_SL g1791 ( 
.A1(n_1775),
.A2(n_124),
.B(n_125),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_R g1792 ( 
.A(n_1783),
.B(n_125),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_SL g1793 ( 
.A(n_1776),
.B(n_1609),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1772),
.A2(n_126),
.B(n_127),
.Y(n_1794)
);

OAI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1782),
.A2(n_127),
.B(n_128),
.C(n_1491),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1778),
.B(n_1491),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1774),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1771),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1780),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1773),
.Y(n_1800)
);

BUFx8_ASAP7_75t_SL g1801 ( 
.A(n_1788),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1798),
.A2(n_1491),
.B1(n_1413),
.B2(n_1581),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1790),
.B(n_182),
.Y(n_1803)
);

OAI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1797),
.A2(n_1491),
.B1(n_1413),
.B2(n_1581),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1791),
.A2(n_1584),
.B1(n_1587),
.B2(n_1590),
.Y(n_1805)
);

OAI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1787),
.A2(n_188),
.B1(n_190),
.B2(n_192),
.C(n_193),
.Y(n_1806)
);

OAI21xp33_ASAP7_75t_L g1807 ( 
.A1(n_1795),
.A2(n_1590),
.B(n_1587),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1786),
.B(n_194),
.Y(n_1808)
);

AOI311xp33_ASAP7_75t_L g1809 ( 
.A1(n_1800),
.A2(n_195),
.A3(n_196),
.B(n_197),
.C(n_199),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1789),
.B(n_201),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1794),
.B(n_202),
.Y(n_1811)
);

NAND4xp75_ASAP7_75t_L g1812 ( 
.A(n_1793),
.B(n_204),
.C(n_205),
.D(n_206),
.Y(n_1812)
);

OAI211xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1785),
.A2(n_207),
.B(n_209),
.C(n_211),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1796),
.Y(n_1814)
);

OAI211xp5_ASAP7_75t_L g1815 ( 
.A1(n_1792),
.A2(n_212),
.B(n_213),
.C(n_218),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1799),
.Y(n_1816)
);

NOR3xp33_ASAP7_75t_L g1817 ( 
.A(n_1785),
.B(n_219),
.C(n_220),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1801),
.Y(n_1818)
);

NOR3xp33_ASAP7_75t_L g1819 ( 
.A(n_1815),
.B(n_222),
.C(n_223),
.Y(n_1819)
);

NAND3xp33_ASAP7_75t_SL g1820 ( 
.A(n_1816),
.B(n_224),
.C(n_227),
.Y(n_1820)
);

NAND5xp2_ASAP7_75t_L g1821 ( 
.A(n_1809),
.B(n_229),
.C(n_231),
.D(n_232),
.E(n_235),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1806),
.B(n_236),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_SL g1823 ( 
.A(n_1812),
.B(n_237),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1810),
.A2(n_238),
.B1(n_241),
.B2(n_243),
.Y(n_1824)
);

OAI222xp33_ASAP7_75t_L g1825 ( 
.A1(n_1814),
.A2(n_1803),
.B1(n_1811),
.B2(n_1808),
.C1(n_1802),
.C2(n_1804),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1817),
.A2(n_1807),
.B1(n_1813),
.B2(n_1805),
.Y(n_1826)
);

NAND4xp25_ASAP7_75t_SL g1827 ( 
.A(n_1806),
.B(n_245),
.C(n_246),
.D(n_247),
.Y(n_1827)
);

CKINVDCx20_ASAP7_75t_R g1828 ( 
.A(n_1801),
.Y(n_1828)
);

OAI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1806),
.A2(n_252),
.B1(n_254),
.B2(n_256),
.C(n_257),
.Y(n_1829)
);

NOR2x1_ASAP7_75t_L g1830 ( 
.A(n_1828),
.B(n_258),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1818),
.Y(n_1831)
);

CKINVDCx5p33_ASAP7_75t_R g1832 ( 
.A(n_1820),
.Y(n_1832)
);

BUFx4f_ASAP7_75t_SL g1833 ( 
.A(n_1825),
.Y(n_1833)
);

CKINVDCx12_ASAP7_75t_R g1834 ( 
.A(n_1824),
.Y(n_1834)
);

OAI21xp33_ASAP7_75t_L g1835 ( 
.A1(n_1821),
.A2(n_1823),
.B(n_1826),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1822),
.Y(n_1836)
);

INVxp67_ASAP7_75t_L g1837 ( 
.A(n_1829),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1819),
.B(n_260),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1831),
.Y(n_1839)
);

INVx2_ASAP7_75t_SL g1840 ( 
.A(n_1830),
.Y(n_1840)
);

NAND4xp25_ASAP7_75t_L g1841 ( 
.A(n_1835),
.B(n_1827),
.C(n_264),
.D(n_266),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1834),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1833),
.Y(n_1843)
);

OAI22xp33_ASAP7_75t_SL g1844 ( 
.A1(n_1838),
.A2(n_261),
.B1(n_267),
.B2(n_274),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1832),
.Y(n_1845)
);

AOI32xp33_ASAP7_75t_L g1846 ( 
.A1(n_1839),
.A2(n_1836),
.A3(n_1837),
.B1(n_1598),
.B2(n_1600),
.Y(n_1846)
);

AOI21xp33_ASAP7_75t_L g1847 ( 
.A1(n_1843),
.A2(n_275),
.B(n_276),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1841),
.A2(n_279),
.B(n_280),
.Y(n_1848)
);

AOI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1842),
.A2(n_1845),
.B(n_1840),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1849),
.Y(n_1850)
);

OR3x1_ASAP7_75t_L g1851 ( 
.A(n_1847),
.B(n_1844),
.C(n_283),
.Y(n_1851)
);

NOR2x1p5_ASAP7_75t_L g1852 ( 
.A(n_1848),
.B(n_281),
.Y(n_1852)
);

OA21x2_ASAP7_75t_L g1853 ( 
.A1(n_1850),
.A2(n_1846),
.B(n_1598),
.Y(n_1853)
);

NOR2x1_ASAP7_75t_L g1854 ( 
.A(n_1851),
.B(n_289),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1854),
.Y(n_1855)
);

AOI222xp33_ASAP7_75t_L g1856 ( 
.A1(n_1853),
.A2(n_1852),
.B1(n_1600),
.B2(n_1592),
.C1(n_305),
.C2(n_307),
.Y(n_1856)
);

AOI21xp33_ASAP7_75t_SL g1857 ( 
.A1(n_1853),
.A2(n_295),
.B(n_299),
.Y(n_1857)
);

OAI221xp5_ASAP7_75t_R g1858 ( 
.A1(n_1855),
.A2(n_303),
.B1(n_308),
.B2(n_311),
.C(n_313),
.Y(n_1858)
);

AOI22xp33_ASAP7_75t_L g1859 ( 
.A1(n_1856),
.A2(n_1592),
.B1(n_323),
.B2(n_327),
.Y(n_1859)
);

OAI221xp5_ASAP7_75t_R g1860 ( 
.A1(n_1859),
.A2(n_1857),
.B1(n_329),
.B2(n_330),
.C(n_331),
.Y(n_1860)
);

AOI211xp5_ASAP7_75t_L g1861 ( 
.A1(n_1860),
.A2(n_1858),
.B(n_332),
.C(n_334),
.Y(n_1861)
);


endmodule