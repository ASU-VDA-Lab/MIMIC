module fake_netlist_1_7043_n_21 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_21);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_21;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
INVx8_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
OAI22xp33_ASAP7_75t_L g11 ( .A1(n_5), .A2(n_1), .B1(n_7), .B2(n_4), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_6), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_3), .B(n_0), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_2), .B(n_0), .Y(n_14) );
AO21x2_ASAP7_75t_L g15 ( .A1(n_12), .A2(n_8), .B(n_14), .Y(n_15) );
INVx2_ASAP7_75t_SL g16 ( .A(n_15), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
NAND3xp33_ASAP7_75t_L g18 ( .A(n_17), .B(n_13), .C(n_11), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_10), .Y(n_21) );
endmodule