module real_jpeg_21806_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_164;
wire n_48;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_1),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_1),
.A2(n_3),
.B1(n_38),
.B2(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_1),
.A2(n_5),
.B1(n_24),
.B2(n_38),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_2),
.A2(n_57),
.B(n_60),
.C(n_63),
.Y(n_59)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_62),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_3),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_3),
.A2(n_7),
.B1(n_40),
.B2(n_57),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_3),
.A2(n_40),
.B(n_62),
.C(n_107),
.Y(n_106)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_4),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_5),
.B(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_5),
.A2(n_8),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_5),
.A2(n_9),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_10),
.B1(n_24),
.B2(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_5),
.A2(n_7),
.B1(n_24),
.B2(n_40),
.Y(n_84)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_5),
.A2(n_7),
.B(n_10),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_33),
.B1(n_35),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_7),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_52)
);

AOI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_7),
.A2(n_45),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_66),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_7),
.A2(n_35),
.B(n_49),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_8),
.A2(n_25),
.B1(n_33),
.B2(n_35),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_10),
.Y(n_34)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_115),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_113),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_95),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_15),
.B(n_95),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_79),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_68),
.B2(n_69),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_41),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_20),
.A2(n_30),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_21),
.B(n_22),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_23),
.A2(n_26),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_24),
.B(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_27),
.A2(n_83),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_28),
.B(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_30),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_30),
.A2(n_100),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_30),
.B(n_108),
.C(n_165),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_30),
.A2(n_100),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_30),
.B(n_183),
.C(n_188),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_31),
.B(n_39),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_31),
.B(n_36),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_36),
.Y(n_31)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_35),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_34),
.A2(n_35),
.B(n_40),
.C(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_36),
.A2(n_71),
.B(n_72),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_36),
.B(n_40),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_39),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_40),
.B(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_40),
.B(n_48),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_40),
.A2(n_45),
.B(n_50),
.C(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_55),
.B2(n_67),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_42),
.A2(n_43),
.B1(n_122),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_42),
.A2(n_43),
.B1(n_85),
.B2(n_86),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_43),
.B(n_93),
.C(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_43),
.B(n_86),
.C(n_171),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_47),
.B(n_51),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_44),
.Y(n_112)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_48),
.B(n_49),
.C(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_47),
.B(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_48),
.A2(n_52),
.B1(n_53),
.B2(n_112),
.Y(n_111)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_55),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_104),
.C(n_110),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_67),
.B1(n_110),
.B2(n_111),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_58),
.B1(n_64),
.B2(n_66),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_66),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_65),
.Y(n_94)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_78),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_70),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_77),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_89),
.C(n_93),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_85),
.B1(n_86),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_81),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_85),
.A2(n_86),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_86),
.B(n_149),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_93),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_98),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.C(n_102),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_96),
.B(n_99),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_102),
.A2(n_103),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

NOR2x1_ASAP7_75t_R g156 ( 
.A(n_108),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_108),
.B(n_157),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_108),
.A2(n_133),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_109),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_110),
.A2(n_111),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_135),
.C(n_137),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

O2A1O1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_140),
.B(n_196),
.C(n_201),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_117),
.B(n_127),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_119),
.B(n_121),
.C(n_125),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_122),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_124),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_134),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_128),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_129),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_134),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_147),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_195),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_190),
.B(n_194),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_180),
.B(n_189),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_168),
.B(n_179),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_160),
.B(n_167),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_151),
.B(n_159),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_156),
.B(n_158),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_162),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_163),
.Y(n_166)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_170),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_177),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_172),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_177),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_182),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_197),
.B(n_198),
.Y(n_201)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);


endmodule