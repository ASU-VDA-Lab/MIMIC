module real_aes_9316_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_905;
wire n_673;
wire n_386;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_102;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_602;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_546;
wire n_151;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
wire n_862;
NAND2xp5_ASAP7_75t_L g632 ( .A(n_0), .B(n_232), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_1), .A2(n_81), .B1(n_631), .B2(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_2), .B(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_3), .B(n_165), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g636 ( .A(n_4), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_5), .A2(n_37), .B1(n_156), .B2(n_562), .Y(n_647) );
INVx1_ASAP7_75t_L g107 ( .A(n_6), .Y(n_107) );
NOR2xp67_ASAP7_75t_L g124 ( .A(n_6), .B(n_83), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_7), .B(n_162), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_8), .B(n_144), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_9), .A2(n_61), .B1(n_156), .B2(n_221), .Y(n_563) );
NAND3xp33_ASAP7_75t_L g595 ( .A(n_10), .B(n_156), .C(n_199), .Y(n_595) );
NAND2x1p5_ASAP7_75t_L g188 ( .A(n_11), .B(n_144), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_12), .B(n_198), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_13), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_14), .B(n_591), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_15), .B(n_153), .Y(n_618) );
AND2x2_ASAP7_75t_L g220 ( .A(n_16), .B(n_221), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_17), .B(n_157), .C(n_162), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_18), .Y(n_913) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_19), .A2(n_27), .B1(n_162), .B2(n_562), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_20), .B(n_591), .Y(n_605) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_21), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_22), .B(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_23), .B(n_231), .Y(n_256) );
NAND2xp33_ASAP7_75t_L g181 ( .A(n_24), .B(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g906 ( .A(n_25), .Y(n_906) );
NAND2xp33_ASAP7_75t_L g243 ( .A(n_26), .B(n_182), .Y(n_243) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_28), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_29), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_30), .B(n_582), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_31), .A2(n_51), .B1(n_182), .B2(n_221), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_32), .B(n_157), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_33), .B(n_164), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_34), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g123 ( .A(n_34), .Y(n_123) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_35), .A2(n_64), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_36), .A2(n_184), .B(n_226), .C(n_228), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_38), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_39), .B(n_156), .Y(n_155) );
NAND2xp33_ASAP7_75t_L g202 ( .A(n_40), .B(n_196), .Y(n_202) );
AND2x6_ASAP7_75t_L g170 ( .A(n_41), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g565 ( .A(n_42), .B(n_173), .Y(n_565) );
NAND2x1p5_ASAP7_75t_L g596 ( .A(n_43), .B(n_173), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_44), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_45), .B(n_227), .Y(n_242) );
NAND2xp33_ASAP7_75t_L g255 ( .A(n_46), .B(n_196), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_47), .B(n_153), .Y(n_607) );
INVx1_ASAP7_75t_L g171 ( .A(n_48), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_49), .Y(n_290) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_50), .A2(n_546), .B1(n_547), .B2(n_900), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_50), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g901 ( .A1(n_50), .A2(n_132), .B1(n_133), .B2(n_546), .Y(n_901) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_52), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_53), .B(n_173), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_54), .B(n_162), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_55), .Y(n_150) );
AND2x2_ASAP7_75t_L g110 ( .A(n_56), .B(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_57), .B(n_162), .Y(n_580) );
AND2x2_ASAP7_75t_L g230 ( .A(n_58), .B(n_231), .Y(n_230) );
NAND2x1_ASAP7_75t_L g612 ( .A(n_59), .B(n_173), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_60), .B(n_199), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_62), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_63), .B(n_573), .Y(n_572) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_65), .Y(n_186) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_66), .Y(n_577) );
OAI22xp33_ASAP7_75t_L g131 ( .A1(n_67), .A2(n_132), .B1(n_133), .B2(n_532), .Y(n_131) );
INVx1_ASAP7_75t_L g532 ( .A(n_67), .Y(n_532) );
NAND2xp33_ASAP7_75t_L g263 ( .A(n_68), .B(n_153), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_69), .B(n_199), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_70), .A2(n_74), .B1(n_162), .B2(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_71), .B(n_180), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g640 ( .A(n_72), .Y(n_640) );
BUFx10_ASAP7_75t_L g536 ( .A(n_73), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_75), .B(n_152), .Y(n_239) );
INVx1_ASAP7_75t_SL g677 ( .A(n_76), .Y(n_677) );
NAND2xp33_ASAP7_75t_L g269 ( .A(n_77), .B(n_162), .Y(n_269) );
CKINVDCx5p33_ASAP7_75t_R g650 ( .A(n_78), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_79), .B(n_182), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_80), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_82), .Y(n_229) );
INVx1_ASAP7_75t_L g106 ( .A(n_83), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_84), .Y(n_115) );
INVx2_ASAP7_75t_L g147 ( .A(n_85), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_86), .B(n_199), .Y(n_594) );
INVx1_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
OR2x2_ASAP7_75t_L g120 ( .A(n_87), .B(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g544 ( .A(n_87), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_87), .B(n_122), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_88), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_89), .B(n_196), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_90), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_91), .B(n_173), .Y(n_204) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_92), .Y(n_250) );
INVx1_ASAP7_75t_L g111 ( .A(n_93), .Y(n_111) );
INVx1_ASAP7_75t_L g219 ( .A(n_94), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_95), .Y(n_284) );
AND2x2_ASAP7_75t_L g291 ( .A(n_96), .B(n_144), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_97), .B(n_218), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_98), .B(n_231), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_113), .B(n_912), .Y(n_99) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx4_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx5_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
BUFx3_ASAP7_75t_L g915 ( .A(n_104), .Y(n_915) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
NOR2xp33_ASAP7_75t_SL g105 ( .A(n_106), .B(n_107), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g109 ( .A(n_110), .B(n_112), .Y(n_109) );
OR2x6_ASAP7_75t_L g113 ( .A(n_114), .B(n_125), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_114), .A2(n_127), .B(n_131), .Y(n_126) );
NOR2x1_ASAP7_75t_R g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx4_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx4_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_120), .Y(n_130) );
AND2x2_ASAP7_75t_L g543 ( .A(n_121), .B(n_544), .Y(n_543) );
AND2x4_ASAP7_75t_L g903 ( .A(n_121), .B(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_533), .B(n_537), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx12f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR3x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_385), .C(n_468), .Y(n_135) );
NAND4xp75_ASAP7_75t_L g136 ( .A(n_137), .B(n_320), .C(n_351), .D(n_366), .Y(n_136) );
NOR2x1_ASAP7_75t_L g137 ( .A(n_138), .B(n_257), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_205), .Y(n_138) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_139), .A2(n_342), .B(n_349), .Y(n_341) );
INVx2_ASAP7_75t_L g388 ( .A(n_139), .Y(n_388) );
AND2x2_ASAP7_75t_L g448 ( .A(n_139), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_175), .Y(n_139) );
AND2x4_ASAP7_75t_L g364 ( .A(n_140), .B(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g443 ( .A(n_140), .B(n_311), .Y(n_443) );
INVx2_ASAP7_75t_L g473 ( .A(n_140), .Y(n_473) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g344 ( .A(n_142), .Y(n_344) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_142), .Y(n_395) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_148), .B(n_172), .Y(n_142) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_143), .A2(n_177), .B(n_188), .Y(n_176) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_143), .A2(n_248), .B(n_256), .Y(n_247) );
OA21x2_ASAP7_75t_L g297 ( .A1(n_143), .A2(n_177), .B(n_188), .Y(n_297) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_143), .A2(n_148), .B(n_172), .Y(n_313) );
BUFx4f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
INVx4_ASAP7_75t_L g213 ( .A(n_144), .Y(n_213) );
OA21x2_ASAP7_75t_L g260 ( .A1(n_144), .A2(n_261), .B(n_270), .Y(n_260) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_144), .A2(n_261), .B(n_270), .Y(n_300) );
OA21x2_ASAP7_75t_L g348 ( .A1(n_144), .A2(n_261), .B(n_270), .Y(n_348) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_144), .Y(n_721) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_145), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g232 ( .A(n_146), .Y(n_232) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_158), .B(n_168), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_155), .C(n_157), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
INVx2_ASAP7_75t_L g265 ( .A(n_153), .Y(n_265) );
INVx1_ASAP7_75t_L g609 ( .A(n_153), .Y(n_609) );
INVx2_ASAP7_75t_L g631 ( .A(n_153), .Y(n_631) );
INVx2_ASAP7_75t_L g638 ( .A(n_153), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_153), .B(n_640), .Y(n_639) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_154), .Y(n_156) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
INVx2_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
INVx1_ASAP7_75t_L g223 ( .A(n_154), .Y(n_223) );
INVx5_ASAP7_75t_L g268 ( .A(n_156), .Y(n_268) );
BUFx12f_ASAP7_75t_L g167 ( .A(n_157), .Y(n_167) );
INVx5_ASAP7_75t_L g184 ( .A(n_157), .Y(n_184) );
INVx5_ASAP7_75t_L g199 ( .A(n_157), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_157), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
OAI321xp33_ASAP7_75t_L g628 ( .A1(n_157), .A2(n_162), .A3(n_629), .B1(n_630), .B2(n_631), .C(n_632), .Y(n_628) );
O2A1O1Ixp33_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_160), .B(n_163), .C(n_166), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_L g185 ( .A1(n_160), .A2(n_166), .B(n_186), .C(n_187), .Y(n_185) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g180 ( .A(n_162), .Y(n_180) );
INVx2_ASAP7_75t_SL g227 ( .A(n_162), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_162), .B(n_282), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_L g576 ( .A1(n_162), .A2(n_199), .B(n_577), .C(n_578), .Y(n_576) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g182 ( .A(n_165), .Y(n_182) );
INVx2_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
O2A1O1Ixp5_ASAP7_75t_L g249 ( .A1(n_166), .A2(n_250), .B(n_251), .C(n_252), .Y(n_249) );
OA22x2_ASAP7_75t_L g560 ( .A1(n_166), .A2(n_183), .B1(n_561), .B2(n_563), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_166), .A2(n_183), .B1(n_673), .B2(n_674), .Y(n_672) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_167), .A2(n_201), .B(n_202), .Y(n_200) );
BUFx2_ASAP7_75t_L g224 ( .A(n_167), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_167), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_167), .A2(n_580), .B(n_581), .Y(n_579) );
AOI21x1_ASAP7_75t_L g606 ( .A1(n_167), .A2(n_607), .B(n_608), .Y(n_606) );
OAI21x1_ASAP7_75t_L g177 ( .A1(n_168), .A2(n_178), .B(n_185), .Y(n_177) );
OAI21x1_ASAP7_75t_L g236 ( .A1(n_168), .A2(n_237), .B(n_241), .Y(n_236) );
OAI21xp5_ASAP7_75t_L g248 ( .A1(n_168), .A2(n_249), .B(n_253), .Y(n_248) );
OAI21x1_ASAP7_75t_L g261 ( .A1(n_168), .A2(n_262), .B(n_266), .Y(n_261) );
AND2x2_ASAP7_75t_L g645 ( .A(n_168), .B(n_192), .Y(n_645) );
AO31x2_ASAP7_75t_L g671 ( .A1(n_168), .A2(n_213), .A3(n_672), .B(n_676), .Y(n_671) );
INVx8_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp67_ASAP7_75t_L g211 ( .A(n_169), .B(n_212), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_169), .A2(n_280), .B(n_286), .Y(n_279) );
INVx1_ASAP7_75t_L g559 ( .A(n_169), .Y(n_559) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_169), .A2(n_632), .B(n_642), .Y(n_641) );
INVx8_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
BUFx2_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
INVx1_ASAP7_75t_L g584 ( .A(n_170), .Y(n_584) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_170), .A2(n_588), .B(n_593), .Y(n_587) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_170), .A2(n_617), .B(n_620), .Y(n_616) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g370 ( .A(n_175), .Y(n_370) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_175), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_189), .Y(n_175) );
INVx2_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_181), .B(n_183), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_182), .B(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_183), .A2(n_254), .B(n_255), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_183), .A2(n_263), .B(n_264), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_183), .A2(n_240), .B1(n_647), .B2(n_648), .Y(n_646) );
CKINVDCx6p67_ASAP7_75t_R g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_SL g285 ( .A(n_184), .Y(n_285) );
AOI21x1_ASAP7_75t_L g603 ( .A1(n_184), .A2(n_604), .B(n_605), .Y(n_603) );
AOI21x1_ASAP7_75t_L g617 ( .A1(n_184), .A2(n_618), .B(n_619), .Y(n_617) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_184), .A2(n_634), .B(n_639), .Y(n_633) );
INVx2_ASAP7_75t_L g275 ( .A(n_189), .Y(n_275) );
OR2x2_ASAP7_75t_L g336 ( .A(n_189), .B(n_313), .Y(n_336) );
AND2x2_ASAP7_75t_L g365 ( .A(n_189), .B(n_274), .Y(n_365) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_193), .B(n_204), .Y(n_190) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_191), .A2(n_236), .B(n_245), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_191), .A2(n_193), .B(n_204), .Y(n_302) );
OAI21x1_ASAP7_75t_L g586 ( .A1(n_191), .A2(n_587), .B(n_596), .Y(n_586) );
OAI21x1_ASAP7_75t_L g658 ( .A1(n_191), .A2(n_587), .B(n_596), .Y(n_658) );
INVx2_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
OAI21x1_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_200), .B(n_203), .Y(n_193) );
AOI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_197), .B(n_199), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_196), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g251 ( .A(n_198), .Y(n_251) );
INVx1_ASAP7_75t_L g244 ( .A(n_199), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_199), .A2(n_267), .B(n_269), .Y(n_266) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_203), .A2(n_603), .B(n_606), .Y(n_602) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_233), .Y(n_206) );
OR2x2_ASAP7_75t_L g436 ( .A(n_207), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g467 ( .A(n_207), .Y(n_467) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g276 ( .A(n_208), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g500 ( .A(n_208), .B(n_353), .Y(n_500) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_209), .B(n_318), .Y(n_340) );
INVx1_ASAP7_75t_L g446 ( .A(n_209), .Y(n_446) );
INVxp67_ASAP7_75t_SL g515 ( .A(n_209), .Y(n_515) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g307 ( .A(n_210), .Y(n_307) );
AOI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_230), .Y(n_210) );
OAI21x1_ASAP7_75t_L g601 ( .A1(n_212), .A2(n_602), .B(n_612), .Y(n_601) );
OAI21x1_ASAP7_75t_L g615 ( .A1(n_212), .A2(n_616), .B(n_624), .Y(n_615) );
OAI21x1_ASAP7_75t_L g655 ( .A1(n_212), .A2(n_602), .B(n_612), .Y(n_655) );
OAI21x1_ASAP7_75t_L g668 ( .A1(n_212), .A2(n_616), .B(n_624), .Y(n_668) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AO21x2_ASAP7_75t_L g278 ( .A1(n_213), .A2(n_279), .B(n_291), .Y(n_278) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_213), .A2(n_279), .B(n_291), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_225), .Y(n_214) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B(n_224), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_219), .Y(n_216) );
NOR2xp33_ASAP7_75t_SL g289 ( .A(n_217), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g562 ( .A(n_218), .Y(n_562) );
INVx2_ASAP7_75t_L g582 ( .A(n_218), .Y(n_582) );
INVx2_ASAP7_75t_L g591 ( .A(n_218), .Y(n_591) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g675 ( .A(n_223), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g593 ( .A1(n_226), .A2(n_594), .B(n_595), .Y(n_593) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx2_ASAP7_75t_L g558 ( .A(n_231), .Y(n_558) );
BUFx5_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g574 ( .A(n_232), .Y(n_574) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_232), .Y(n_642) );
INVx1_ASAP7_75t_SL g308 ( .A(n_233), .Y(n_308) );
INVx1_ASAP7_75t_L g431 ( .A(n_233), .Y(n_431) );
OR2x2_ASAP7_75t_L g519 ( .A(n_233), .B(n_335), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_233), .B(n_403), .Y(n_528) );
OR2x2_ASAP7_75t_L g233 ( .A(n_234), .B(n_246), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g277 ( .A(n_235), .B(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g324 ( .A(n_235), .B(n_246), .Y(n_324) );
INVx1_ASAP7_75t_L g339 ( .A(n_235), .Y(n_339) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_235), .Y(n_375) );
AND2x2_ASAP7_75t_L g411 ( .A(n_235), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g439 ( .A(n_235), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_240), .Y(n_237) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_240), .A2(n_287), .B(n_289), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_244), .Y(n_241) );
BUFx3_ASAP7_75t_L g392 ( .A(n_246), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_246), .B(n_306), .Y(n_497) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g318 ( .A(n_247), .Y(n_318) );
OAI21xp5_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_276), .B(n_292), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_271), .Y(n_259) );
INVx2_ASAP7_75t_L g331 ( .A(n_260), .Y(n_331) );
INVx2_ASAP7_75t_L g363 ( .A(n_260), .Y(n_363) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_260), .Y(n_449) );
AND2x2_ASAP7_75t_L g501 ( .A(n_260), .B(n_301), .Y(n_501) );
NOR2xp67_ASAP7_75t_L g283 ( .A(n_268), .B(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_271), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g394 ( .A(n_272), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x2_ASAP7_75t_L g312 ( .A(n_273), .B(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g381 ( .A(n_273), .B(n_348), .Y(n_381) );
AND2x2_ASAP7_75t_L g427 ( .A(n_273), .B(n_348), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_273), .Y(n_434) );
OR2x2_ASAP7_75t_L g499 ( .A(n_273), .B(n_299), .Y(n_499) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g311 ( .A(n_275), .Y(n_311) );
AND2x2_ASAP7_75t_L g332 ( .A(n_275), .B(n_297), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g387 ( .A1(n_276), .A2(n_383), .B1(n_388), .B2(n_389), .Y(n_387) );
INVx2_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
OR2x2_ASAP7_75t_L g383 ( .A(n_277), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g325 ( .A(n_278), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g350 ( .A(n_278), .B(n_307), .Y(n_350) );
OAI21xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B(n_285), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_303), .B1(n_309), .B2(n_314), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_294), .A2(n_337), .B1(n_407), .B2(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
AND2x2_ASAP7_75t_L g484 ( .A(n_295), .B(n_328), .Y(n_484) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_296), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_296), .B(n_344), .Y(n_494) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g335 ( .A(n_299), .Y(n_335) );
INVx2_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_SL g358 ( .A(n_300), .Y(n_358) );
BUFx2_ASAP7_75t_L g425 ( .A(n_300), .Y(n_425) );
INVx1_ASAP7_75t_L g493 ( .A(n_300), .Y(n_493) );
BUFx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g329 ( .A(n_302), .B(n_313), .Y(n_329) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_308), .Y(n_303) );
AND2x2_ASAP7_75t_L g405 ( .A(n_304), .B(n_392), .Y(n_405) );
AND2x4_ASAP7_75t_L g476 ( .A(n_304), .B(n_324), .Y(n_476) );
INVx1_ASAP7_75t_L g491 ( .A(n_304), .Y(n_491) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_305), .Y(n_510) );
INVx2_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_306), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g403 ( .A(n_306), .Y(n_403) );
INVx1_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
INVx1_ASAP7_75t_L g412 ( .A(n_307), .Y(n_412) );
INVx1_ASAP7_75t_L g407 ( .A(n_309), .Y(n_407) );
AND2x4_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x4_ASAP7_75t_SL g417 ( .A(n_311), .B(n_344), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_313), .Y(n_420) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g428 ( .A(n_316), .B(n_384), .Y(n_428) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
INVxp67_ASAP7_75t_L g466 ( .A(n_317), .Y(n_466) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g374 ( .A(n_318), .B(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_318), .B(n_319), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_318), .B(n_403), .Y(n_409) );
AND2x2_ASAP7_75t_L g438 ( .A(n_318), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_318), .B(n_446), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_327), .B(n_333), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g480 ( .A(n_323), .Y(n_480) );
NAND2xp67_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g349 ( .A(n_324), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g397 ( .A(n_324), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_324), .B(n_350), .Y(n_460) );
AND2x4_ASAP7_75t_L g372 ( .A(n_325), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g399 ( .A(n_325), .Y(n_399) );
INVx1_ASAP7_75t_L g384 ( .A(n_326), .Y(n_384) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
AND2x2_ASAP7_75t_L g379 ( .A(n_328), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g389 ( .A(n_328), .Y(n_389) );
BUFx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g360 ( .A(n_329), .Y(n_360) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OAI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_337), .B(n_341), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_334), .A2(n_463), .B1(n_465), .B2(n_466), .Y(n_462) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g459 ( .A(n_335), .Y(n_459) );
OR2x2_ASAP7_75t_L g337 ( .A(n_338), .B(n_340), .Y(n_337) );
INVx1_ASAP7_75t_L g353 ( .A(n_338), .Y(n_353) );
OR2x2_ASAP7_75t_L g444 ( .A(n_338), .B(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
AND2x2_ASAP7_75t_L g475 ( .A(n_343), .B(n_427), .Y(n_475) );
INVx1_ASAP7_75t_L g517 ( .A(n_343), .Y(n_517) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx2_ASAP7_75t_L g371 ( .A(n_344), .Y(n_371) );
AND2x2_ASAP7_75t_L g472 ( .A(n_345), .B(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVxp67_ASAP7_75t_SL g507 ( .A(n_346), .Y(n_507) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_348), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g430 ( .A(n_350), .B(n_431), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_350), .B(n_456), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_350), .B(n_483), .Y(n_482) );
NAND2x1_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_361), .Y(n_354) );
INVxp33_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_359), .Y(n_356) );
AND2x2_ASAP7_75t_L g525 ( .A(n_357), .B(n_443), .Y(n_525) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2x1_ASAP7_75t_SL g498 ( .A(n_360), .B(n_499), .Y(n_498) );
INVxp67_ASAP7_75t_L g486 ( .A(n_361), .Y(n_486) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
AND2x2_ASAP7_75t_L g391 ( .A(n_363), .B(n_392), .Y(n_391) );
AO22x1_ASAP7_75t_L g376 ( .A1(n_364), .A2(n_377), .B1(n_379), .B2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g423 ( .A(n_365), .B(n_424), .Y(n_423) );
AND2x2_ASAP7_75t_L g516 ( .A(n_365), .B(n_517), .Y(n_516) );
O2A1O1Ixp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_371), .B(n_372), .C(n_376), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_368), .A2(n_448), .B1(n_450), .B2(n_452), .C(n_457), .Y(n_447) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g464 ( .A(n_369), .B(n_441), .Y(n_464) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_371), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g401 ( .A(n_374), .Y(n_401) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g531 ( .A(n_381), .Y(n_531) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g523 ( .A(n_384), .Y(n_523) );
NAND4xp75_ASAP7_75t_L g385 ( .A(n_386), .B(n_413), .C(n_447), .D(n_461), .Y(n_385) );
AOI221x1_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B1(n_393), .B2(n_396), .C(n_406), .Y(n_386) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g483 ( .A(n_392), .Y(n_483) );
INVx2_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_397), .A2(n_398), .B(n_400), .C(n_404), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_397), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g465 ( .A(n_401), .Y(n_465) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_429), .Y(n_413) );
OAI21xp5_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_421), .B(n_428), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_418), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g520 ( .A1(n_416), .A2(n_521), .B(n_522), .Y(n_520) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_417), .B(n_531), .Y(n_530) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g441 ( .A(n_419), .Y(n_441) );
BUFx2_ASAP7_75t_L g479 ( .A(n_420), .Y(n_479) );
NAND2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B(n_435), .Y(n_429) );
AND2x2_ASAP7_75t_L g513 ( .A(n_431), .B(n_514), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_432), .A2(n_480), .B(n_504), .C(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_440), .B1(n_442), .B2(n_444), .Y(n_435) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_438), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g456 ( .A(n_439), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_441), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_443), .B(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g487 ( .A(n_445), .Y(n_487) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_467), .Y(n_461) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND4xp75_ASAP7_75t_L g468 ( .A(n_469), .B(n_485), .C(n_502), .D(n_511), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_476), .B(n_477), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx2_ASAP7_75t_L g504 ( .A(n_473), .Y(n_504) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AO22x1_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_480), .B1(n_481), .B2(n_484), .Y(n_477) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_488), .Y(n_485) );
OAI21xp5_ASAP7_75t_SL g488 ( .A1(n_489), .A2(n_492), .B(n_495), .Y(n_488) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_490), .A2(n_525), .B1(n_526), .B2(n_529), .Y(n_524) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OR2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_498), .B1(n_500), .B2(n_501), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_504), .A2(n_506), .B(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g521 ( .A(n_509), .Y(n_521) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_524), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_516), .B1(n_518), .B2(n_520), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
INVx11_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx12f_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx6_ASAP7_75t_L g542 ( .A(n_536), .Y(n_542) );
INVx2_ASAP7_75t_SL g910 ( .A(n_536), .Y(n_910) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_545), .B1(n_901), .B2(n_902), .C(n_905), .Y(n_537) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_543), .Y(n_540) );
AND2x6_ASAP7_75t_SL g902 ( .A(n_541), .B(n_903), .Y(n_902) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g904 ( .A(n_544), .Y(n_904) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g900 ( .A(n_548), .Y(n_900) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_807), .Y(n_549) );
NOR3xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_730), .C(n_770), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_685), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_566), .B1(n_660), .B2(n_669), .C1(n_678), .C2(n_683), .Y(n_552) );
INVx2_ASAP7_75t_L g782 ( .A(n_553), .Y(n_782) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g751 ( .A(n_554), .B(n_704), .Y(n_751) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g796 ( .A(n_555), .B(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g845 ( .A(n_555), .B(n_689), .Y(n_845) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_556), .B(n_671), .Y(n_681) );
INVx1_ASAP7_75t_L g690 ( .A(n_556), .Y(n_690) );
INVx1_ASAP7_75t_L g708 ( .A(n_556), .Y(n_708) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_556), .Y(n_801) );
INVxp67_ASAP7_75t_SL g869 ( .A(n_556), .Y(n_869) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_564), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
OA21x2_ASAP7_75t_L g720 ( .A1(n_560), .A2(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVxp67_ASAP7_75t_L g722 ( .A(n_565), .Y(n_722) );
OAI21xp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_597), .B(n_651), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g767 ( .A(n_568), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_568), .B(n_748), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_568), .B(n_768), .Y(n_886) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_585), .Y(n_569) );
AND2x4_ASAP7_75t_L g689 ( .A(n_570), .B(n_670), .Y(n_689) );
AND2x2_ASAP7_75t_L g728 ( .A(n_570), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx2_ASAP7_75t_L g706 ( .A(n_571), .Y(n_706) );
AND2x2_ASAP7_75t_L g794 ( .A(n_571), .B(n_658), .Y(n_794) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_574), .B(n_650), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_574), .B(n_677), .Y(n_676) );
OAI21x1_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_579), .B(n_583), .Y(n_575) );
AND2x2_ASAP7_75t_L g669 ( .A(n_585), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g701 ( .A(n_585), .Y(n_701) );
AND2x2_ASAP7_75t_L g704 ( .A(n_585), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g719 ( .A(n_586), .B(n_720), .Y(n_719) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_590), .B(n_592), .Y(n_588) );
INVxp67_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_625), .Y(n_597) );
INVx2_ASAP7_75t_SL g778 ( .A(n_598), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_598), .B(n_695), .Y(n_795) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_613), .Y(n_598) );
AND2x2_ASAP7_75t_L g700 ( .A(n_599), .B(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_599), .B(n_613), .Y(n_734) );
INVx1_ASAP7_75t_L g774 ( .A(n_599), .Y(n_774) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_600), .Y(n_694) );
OR2x2_ASAP7_75t_L g824 ( .A(n_600), .B(n_643), .Y(n_824) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g725 ( .A(n_601), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g622 ( .A(n_609), .Y(n_622) );
INVx4_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g743 ( .A(n_613), .B(n_667), .Y(n_743) );
AND2x2_ASAP7_75t_L g872 ( .A(n_613), .B(n_776), .Y(n_872) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_SL g659 ( .A(n_614), .Y(n_659) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g780 ( .A(n_615), .Y(n_780) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g709 ( .A(n_626), .B(n_710), .Y(n_709) );
BUFx3_ASAP7_75t_L g769 ( .A(n_626), .Y(n_769) );
AND2x2_ASAP7_75t_L g817 ( .A(n_626), .B(n_711), .Y(n_817) );
AND2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_643), .Y(n_626) );
INVx1_ASAP7_75t_L g656 ( .A(n_627), .Y(n_656) );
INVx2_ASAP7_75t_L g667 ( .A(n_627), .Y(n_667) );
OAI21x1_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_633), .B(n_641), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g665 ( .A(n_643), .Y(n_665) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_643), .Y(n_759) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g697 ( .A(n_644), .Y(n_697) );
AOI21x1_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_646), .B(n_649), .Y(n_644) );
INVxp33_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NOR3xp33_ASAP7_75t_L g652 ( .A(n_653), .B(n_657), .C(n_659), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g815 ( .A(n_654), .B(n_684), .Y(n_815) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx2_ASAP7_75t_L g664 ( .A(n_655), .Y(n_664) );
AND2x2_ASAP7_75t_L g696 ( .A(n_656), .B(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_656), .B(n_725), .Y(n_724) );
INVx2_ASAP7_75t_L g740 ( .A(n_656), .Y(n_740) );
INVx2_ASAP7_75t_L g682 ( .A(n_657), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_657), .B(n_749), .Y(n_885) );
BUFx3_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g797 ( .A(n_658), .B(n_706), .Y(n_797) );
AND2x4_ASAP7_75t_L g830 ( .A(n_659), .B(n_831), .Y(n_830) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_659), .A2(n_821), .B1(n_882), .B2(n_886), .Y(n_881) );
AND2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_666), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
INVx2_ASAP7_75t_L g746 ( .A(n_664), .Y(n_746) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_665), .Y(n_684) );
INVx1_ASAP7_75t_L g777 ( .A(n_665), .Y(n_777) );
AND2x2_ASAP7_75t_L g683 ( .A(n_666), .B(n_684), .Y(n_683) );
INVx2_ASAP7_75t_L g713 ( .A(n_666), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_666), .B(n_774), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_666), .B(n_876), .Y(n_875) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OR2x2_ASAP7_75t_L g733 ( .A(n_667), .B(n_697), .Y(n_733) );
AND2x2_ASAP7_75t_L g804 ( .A(n_667), .B(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g711 ( .A(n_668), .Y(n_711) );
INVx1_ASAP7_75t_L g805 ( .A(n_668), .Y(n_805) );
INVx1_ASAP7_75t_L g729 ( .A(n_670), .Y(n_729) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g717 ( .A(n_671), .Y(n_717) );
INVx1_ASAP7_75t_L g749 ( .A(n_671), .Y(n_749) );
AND2x2_ASAP7_75t_L g768 ( .A(n_671), .B(n_720), .Y(n_768) );
INVxp67_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .Y(n_679) );
AND2x2_ASAP7_75t_L g832 ( .A(n_680), .B(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_680), .B(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVxp67_ASAP7_75t_L g756 ( .A(n_681), .Y(n_756) );
AND2x4_ASAP7_75t_L g783 ( .A(n_682), .B(n_689), .Y(n_783) );
OR2x2_ASAP7_75t_L g877 ( .A(n_682), .B(n_878), .Y(n_877) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_691), .B1(n_698), .B2(n_709), .C(n_712), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI21xp33_ASAP7_75t_L g698 ( .A1(n_687), .A2(n_699), .B(n_702), .Y(n_698) );
OR2x6_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g878 ( .A(n_689), .Y(n_878) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_693), .B(n_896), .Y(n_895) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g762 ( .A(n_694), .B(n_739), .Y(n_762) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x4_ASAP7_75t_L g822 ( .A(n_696), .B(n_787), .Y(n_822) );
AND2x2_ASAP7_75t_L g842 ( .A(n_696), .B(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_697), .B(n_711), .Y(n_789) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_697), .Y(n_806) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g844 ( .A(n_700), .B(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_701), .B(n_801), .Y(n_800) );
OR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_707), .Y(n_702) );
INVx2_ASAP7_75t_L g766 ( .A(n_703), .Y(n_766) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g745 ( .A(n_704), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g755 ( .A(n_704), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g718 ( .A(n_705), .Y(n_718) );
AND2x2_ASAP7_75t_L g840 ( .A(n_705), .B(n_720), .Y(n_840) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g858 ( .A(n_707), .Y(n_858) );
AND2x2_ASAP7_75t_L g899 ( .A(n_707), .B(n_849), .Y(n_899) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g727 ( .A(n_708), .B(n_728), .Y(n_727) );
NOR2x1_ASAP7_75t_L g792 ( .A(n_708), .B(n_765), .Y(n_792) );
INVx2_ASAP7_75t_SL g827 ( .A(n_709), .Y(n_827) );
AND2x2_ASAP7_75t_L g836 ( .A(n_709), .B(n_837), .Y(n_836) );
AND2x4_ASAP7_75t_L g739 ( .A(n_710), .B(n_740), .Y(n_739) );
NOR2xp67_ASAP7_75t_L g753 ( .A(n_710), .B(n_733), .Y(n_753) );
AND2x2_ASAP7_75t_L g812 ( .A(n_710), .B(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_723), .B2(n_726), .Y(n_712) );
INVx1_ASAP7_75t_L g846 ( .A(n_713), .Y(n_846) );
INVx1_ASAP7_75t_L g818 ( .A(n_714), .Y(n_818) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_719), .Y(n_715) );
NOR2xp67_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g765 ( .A(n_717), .Y(n_765) );
INVx1_ASAP7_75t_L g892 ( .A(n_718), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_719), .A2(n_732), .B1(n_735), .B2(n_736), .C(n_741), .Y(n_731) );
AND2x4_ASAP7_75t_L g735 ( .A(n_719), .B(n_728), .Y(n_735) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g776 ( .A(n_725), .B(n_777), .Y(n_776) );
BUFx2_ASAP7_75t_L g837 ( .A(n_725), .Y(n_837) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp67_ASAP7_75t_L g862 ( .A(n_728), .Y(n_862) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_731), .B(n_754), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
OR2x2_ASAP7_75t_L g773 ( .A(n_733), .B(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g860 ( .A(n_733), .B(n_734), .Y(n_860) );
OR2x2_ASAP7_75t_L g879 ( .A(n_733), .B(n_857), .Y(n_879) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OR2x2_ASAP7_75t_L g828 ( .A(n_738), .B(n_774), .Y(n_828) );
INVx4_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g779 ( .A(n_740), .B(n_780), .Y(n_779) );
OAI32xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .A3(n_747), .B1(n_750), .B2(n_752), .Y(n_741) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g823 ( .A(n_743), .B(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AND2x2_ASAP7_75t_L g855 ( .A(n_745), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g788 ( .A(n_746), .Y(n_788) );
AND2x2_ASAP7_75t_L g831 ( .A(n_746), .B(n_777), .Y(n_831) );
AND2x2_ASAP7_75t_L g851 ( .A(n_746), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g799 ( .A(n_748), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
NOR2x1_ASAP7_75t_L g849 ( .A(n_749), .B(n_850), .Y(n_849) );
INVx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVxp67_ASAP7_75t_SL g752 ( .A(n_753), .Y(n_752) );
AOI222xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_757), .B1(n_760), .B2(n_763), .C1(n_767), .C2(n_769), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_L g865 ( .A(n_765), .Y(n_865) );
INVx1_ASAP7_75t_L g820 ( .A(n_766), .Y(n_820) );
OAI211xp5_ASAP7_75t_L g798 ( .A1(n_768), .A2(n_793), .B(n_799), .C(n_802), .Y(n_798) );
INVx2_ASAP7_75t_L g893 ( .A(n_769), .Y(n_893) );
OAI21xp33_ASAP7_75t_L g770 ( .A1(n_771), .A2(n_781), .B(n_784), .Y(n_770) );
NOR4xp25_ASAP7_75t_SL g771 ( .A(n_772), .B(n_775), .C(n_778), .D(n_779), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
BUFx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND2x1_ASAP7_75t_SL g889 ( .A(n_778), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g843 ( .A(n_780), .Y(n_843) );
NAND2x1p5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
AOI221xp5_ASAP7_75t_L g841 ( .A1(n_783), .A2(n_842), .B1(n_844), .B2(n_846), .C(n_847), .Y(n_841) );
AOI322xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_790), .A3(n_793), .B1(n_795), .B2(n_796), .C1(n_798), .C2(n_803), .Y(n_784) );
INVx2_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g852 ( .A(n_789), .Y(n_852) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
O2A1O1Ixp33_ASAP7_75t_L g819 ( .A1(n_791), .A2(n_820), .B(n_821), .C(n_823), .Y(n_819) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g833 ( .A(n_793), .Y(n_833) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
NAND2x1p5_ASAP7_75t_L g867 ( .A(n_794), .B(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g850 ( .A(n_797), .Y(n_850) );
AND2x2_ASAP7_75t_L g803 ( .A(n_804), .B(n_806), .Y(n_803) );
INVx2_ASAP7_75t_L g897 ( .A(n_804), .Y(n_897) );
INVx1_ASAP7_75t_L g813 ( .A(n_806), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_853), .Y(n_807) );
NAND3xp33_ASAP7_75t_SL g808 ( .A(n_809), .B(n_825), .C(n_841), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_818), .B(n_819), .Y(n_809) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .C(n_816), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g876 ( .A(n_824), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_832), .B(n_834), .Y(n_825) );
NAND3xp33_ASAP7_75t_SL g826 ( .A(n_827), .B(n_828), .C(n_829), .Y(n_826) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx2_ASAP7_75t_L g884 ( .A(n_840), .Y(n_884) );
INVx1_ASAP7_75t_L g898 ( .A(n_842), .Y(n_898) );
INVx2_ASAP7_75t_L g857 ( .A(n_843), .Y(n_857) );
INVxp67_ASAP7_75t_L g880 ( .A(n_845), .Y(n_880) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_849), .B(n_851), .Y(n_848) );
INVx2_ASAP7_75t_L g873 ( .A(n_851), .Y(n_873) );
NAND3xp33_ASAP7_75t_SL g853 ( .A(n_854), .B(n_863), .C(n_887), .Y(n_853) );
AOI21xp5_ASAP7_75t_L g854 ( .A1(n_855), .A2(n_858), .B(n_859), .Y(n_854) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
AOI21xp33_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_861), .B(n_862), .Y(n_859) );
AOI211xp5_ASAP7_75t_SL g863 ( .A1(n_864), .A2(n_870), .B(n_874), .C(n_881), .Y(n_863) );
AND2x4_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_871), .B(n_873), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
OAI22xp33_ASAP7_75t_SL g874 ( .A1(n_875), .A2(n_877), .B1(n_879), .B2(n_880), .Y(n_874) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NOR2x1p5_ASAP7_75t_SL g883 ( .A(n_884), .B(n_885), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_888), .A2(n_893), .B1(n_894), .B2(n_899), .Y(n_887) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_895), .B(n_898), .Y(n_894) );
INVx2_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
NOR2xp33_ASAP7_75t_L g905 ( .A(n_906), .B(n_907), .Y(n_905) );
BUFx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
BUFx12f_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OR2x2_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NOR2xp33_ASAP7_75t_SL g912 ( .A(n_913), .B(n_914), .Y(n_912) );
BUFx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
endmodule