module fake_jpeg_29669_n_315 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_9),
.B(n_11),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_7),
.B(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_48),
.Y(n_87)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_27),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_61),
.Y(n_101)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_30),
.B(n_8),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_69),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_68),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_66),
.B(n_39),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_70),
.B(n_81),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_44),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_74),
.B(n_103),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_39),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_28),
.B1(n_42),
.B2(n_40),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_84),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_43),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_102),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_55),
.A2(n_28),
.B1(n_42),
.B2(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_22),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_50),
.A2(n_28),
.B1(n_42),
.B2(n_40),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_34),
.B1(n_42),
.B2(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_22),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_105),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_37),
.B1(n_18),
.B2(n_23),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_96),
.B1(n_104),
.B2(n_62),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_37),
.B1(n_41),
.B2(n_38),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_95),
.A2(n_18),
.B1(n_23),
.B2(n_27),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_43),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_41),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_37),
.B1(n_35),
.B2(n_18),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_26),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_113),
.B(n_9),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_64),
.A2(n_38),
.B1(n_21),
.B2(n_24),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_59),
.B(n_29),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_47),
.B(n_24),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_29),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_115),
.B(n_120),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_73),
.B1(n_76),
.B2(n_89),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_69),
.B1(n_33),
.B2(n_20),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_141),
.B1(n_140),
.B2(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_122),
.Y(n_158)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_35),
.B1(n_33),
.B2(n_21),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_35),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_87),
.C(n_74),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_72),
.B1(n_97),
.B2(n_108),
.Y(n_173)
);

AO21x1_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_12),
.B(n_1),
.Y(n_180)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_135),
.Y(n_162)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_100),
.Y(n_136)
);

BUFx2_ASAP7_75t_SL g178 ( 
.A(n_136),
.Y(n_178)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_81),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_144),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_90),
.A2(n_80),
.B1(n_88),
.B2(n_110),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_146),
.Y(n_176)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_113),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_145),
.B(n_147),
.Y(n_184)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_7),
.B(n_1),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_150),
.Y(n_169)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_112),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_152),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_128),
.B(n_80),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_109),
.B(n_90),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_172),
.B(n_174),
.Y(n_187)
);

O2A1O1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_92),
.B(n_84),
.C(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_166),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_171),
.B1(n_182),
.B2(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_112),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_83),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_170),
.B(n_181),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_83),
.B(n_91),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_180),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_129),
.A2(n_72),
.B(n_91),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_127),
.A2(n_97),
.B(n_0),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_175),
.A2(n_123),
.B(n_0),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_12),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_129),
.A2(n_89),
.B1(n_76),
.B2(n_73),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_89),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_126),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_178),
.Y(n_185)
);

INVx11_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_114),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_190),
.Y(n_218)
);

AO21x2_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_116),
.B(n_137),
.Y(n_189)
);

AO21x1_ASAP7_75t_L g226 ( 
.A1(n_189),
.A2(n_173),
.B(n_155),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_119),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_191),
.A2(n_170),
.B(n_177),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_184),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_194),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_176),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_201),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_118),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_172),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_199),
.A2(n_202),
.B1(n_209),
.B2(n_177),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_159),
.B(n_166),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_154),
.A2(n_149),
.B1(n_147),
.B2(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_135),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

BUFx8_ASAP7_75t_L g208 ( 
.A(n_167),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_175),
.A2(n_146),
.B1(n_130),
.B2(n_124),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_164),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_169),
.B(n_121),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_164),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_165),
.B(n_179),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_169),
.B(n_10),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_161),
.C(n_168),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_227),
.B(n_228),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_204),
.B1(n_209),
.B2(n_205),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_238),
.C(n_212),
.Y(n_240)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_226),
.A2(n_189),
.B(n_204),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_187),
.A2(n_180),
.B(n_152),
.Y(n_227)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_196),
.A2(n_152),
.B(n_159),
.C(n_182),
.D(n_158),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_229),
.A2(n_204),
.B1(n_189),
.B2(n_199),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_186),
.A2(n_168),
.A3(n_161),
.B1(n_165),
.B2(n_163),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_223),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_187),
.A2(n_179),
.B(n_163),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_237),
.A2(n_239),
.B(n_185),
.Y(n_253)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_162),
.C(n_2),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_189),
.A2(n_186),
.B(n_202),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_225),
.C(n_224),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_227),
.B(n_239),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_242),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_220),
.A2(n_189),
.B(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_243),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_244),
.B(n_253),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_198),
.C(n_193),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_246),
.C(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_193),
.C(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_248),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_213),
.C(n_207),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_208),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_252),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_229),
.A2(n_195),
.B1(n_208),
.B2(n_210),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_214),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_255),
.B(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_162),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_76),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_259),
.B(n_216),
.Y(n_260)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_260),
.Y(n_283)
);

OAI322xp33_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_235),
.A3(n_230),
.B1(n_228),
.B2(n_219),
.C1(n_231),
.C2(n_232),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_261),
.B(n_249),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_226),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_267),
.C(n_259),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_245),
.B(n_226),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_246),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_273),
.A2(n_258),
.B1(n_230),
.B2(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_276),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_281),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_258),
.B1(n_252),
.B2(n_253),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_270),
.A2(n_241),
.B1(n_242),
.B2(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_282),
.B1(n_263),
.B2(n_260),
.Y(n_286)
);

AOI31xp67_ASAP7_75t_L g278 ( 
.A1(n_271),
.A2(n_252),
.A3(n_251),
.B(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_266),
.A2(n_251),
.B(n_232),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_219),
.B1(n_225),
.B2(n_217),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_221),
.C(n_2),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_264),
.C(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_10),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_13),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_286),
.A2(n_288),
.B1(n_221),
.B2(n_5),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_277),
.A2(n_271),
.B1(n_265),
.B2(n_267),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_284),
.B(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_290),
.B(n_293),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_269),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_281),
.C(n_283),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_295),
.B(n_13),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_297),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_294),
.B(n_289),
.C(n_291),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_263),
.C(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_300),
.A2(n_287),
.B1(n_292),
.B2(n_298),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_276),
.C(n_274),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_302),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_306),
.B(n_17),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_300),
.A2(n_288),
.B1(n_5),
.B2(n_6),
.Y(n_306)
);

XOR2x2_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_5),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_307),
.C(n_303),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_309),
.A2(n_310),
.B(n_306),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_304),
.A2(n_7),
.B(n_10),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.Y(n_313)
);

AOI321xp33_ASAP7_75t_SL g314 ( 
.A1(n_313),
.A2(n_0),
.A3(n_14),
.B1(n_17),
.B2(n_305),
.C(n_278),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_14),
.Y(n_315)
);


endmodule