module fake_jpeg_16590_n_349 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_2),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_45),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_32),
.A2(n_0),
.B(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_21),
.Y(n_65)
);

OA22x2_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_44),
.A2(n_30),
.B1(n_29),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_58),
.B1(n_70),
.B2(n_78),
.Y(n_102)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_45),
.A2(n_30),
.B1(n_22),
.B2(n_24),
.Y(n_58)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_65),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_39),
.Y(n_66)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g90 ( 
.A(n_68),
.Y(n_90)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_44),
.A2(n_30),
.B1(n_29),
.B2(n_31),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_26),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_26),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_38),
.A2(n_24),
.B1(n_36),
.B2(n_19),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_79),
.Y(n_94)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_107),
.Y(n_118)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_46),
.B1(n_51),
.B2(n_45),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_88),
.A2(n_99),
.B1(n_103),
.B2(n_54),
.Y(n_138)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_101),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_45),
.B1(n_24),
.B2(n_18),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_53),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_58),
.A2(n_42),
.B1(n_46),
.B2(n_52),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_41),
.B1(n_40),
.B2(n_20),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_111),
.B1(n_66),
.B2(n_54),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_18),
.B1(n_23),
.B2(n_19),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_20),
.B1(n_36),
.B2(n_37),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_75),
.Y(n_108)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_49),
.C(n_47),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_39),
.C(n_47),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_40),
.B1(n_41),
.B2(n_19),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_128),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_18),
.B1(n_23),
.B2(n_25),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_133),
.B1(n_140),
.B2(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_77),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_77),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_80),
.B1(n_69),
.B2(n_63),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_124),
.A2(n_82),
.B1(n_94),
.B2(n_108),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_93),
.B(n_25),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_127),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_63),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_99),
.B(n_49),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_88),
.A2(n_28),
.B(n_23),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_138),
.Y(n_150)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_25),
.B(n_35),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_142),
.C(n_49),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_137),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_83),
.B(n_26),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_136),
.B(n_83),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_88),
.A2(n_68),
.B1(n_62),
.B2(n_40),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_49),
.C(n_47),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_144),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_126),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_164),
.B1(n_141),
.B2(n_119),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_90),
.B(n_112),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_155),
.B(n_137),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_97),
.A3(n_82),
.B1(n_36),
.B2(n_20),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_162),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_165),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_121),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_142),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_138),
.A2(n_109),
.B1(n_86),
.B2(n_92),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_94),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_86),
.B1(n_105),
.B2(n_98),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_166),
.A2(n_115),
.B1(n_119),
.B2(n_141),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_100),
.Y(n_167)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_84),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_168),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_170),
.B1(n_188),
.B2(n_189),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_124),
.B1(n_134),
.B2(n_114),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_125),
.B(n_118),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_179),
.B(n_159),
.Y(n_196)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_176),
.A2(n_148),
.B1(n_84),
.B2(n_120),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_158),
.B(n_152),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_186),
.Y(n_200)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_182),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_184),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_146),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_162),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_157),
.A2(n_125),
.B1(n_117),
.B2(n_113),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_129),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_27),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx3_ASAP7_75t_SL g194 ( 
.A(n_182),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_218),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_145),
.B(n_159),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_197),
.A2(n_198),
.B(n_199),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_152),
.B(n_167),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_163),
.B(n_152),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_209),
.C(n_216),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_204),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_176),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_205),
.B(n_211),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_184),
.B(n_180),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_207),
.B(n_212),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_SL g207 ( 
.A(n_172),
.B(n_153),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_149),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g210 ( 
.A1(n_172),
.A2(n_149),
.B(n_164),
.C(n_151),
.D(n_166),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_188),
.C(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_144),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_165),
.B1(n_129),
.B2(n_96),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_175),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_213),
.B(n_171),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_27),
.C(n_120),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_217),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_123),
.B(n_126),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_170),
.B(n_27),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_123),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_169),
.B1(n_178),
.B2(n_191),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_220),
.A2(n_221),
.B1(n_224),
.B2(n_214),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_210),
.A2(n_193),
.B1(n_207),
.B2(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_215),
.A2(n_177),
.B1(n_175),
.B2(n_171),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_200),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_234),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_201),
.B(n_177),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_235),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_160),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_237),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_117),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_120),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_241),
.Y(n_248)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_1),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_230),
.B1(n_236),
.B2(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_219),
.A2(n_242),
.B1(n_232),
.B2(n_225),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_228),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_196),
.C(n_199),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_238),
.B(n_239),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_202),
.C(n_216),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_258),
.C(n_259),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_253),
.B(n_260),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_123),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_261),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_130),
.C(n_71),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_130),
.C(n_161),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_226),
.B(n_238),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_130),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_161),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_33),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_74),
.C(n_27),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_28),
.C(n_33),
.Y(n_279)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_220),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_268),
.C(n_277),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_231),
.C(n_224),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_253),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_249),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_223),
.Y(n_276)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_11),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_28),
.C(n_33),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_257),
.B(n_261),
.C(n_255),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_28),
.C(n_33),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_249),
.C(n_245),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_10),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_264),
.C(n_270),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_283),
.B(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_286),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_296),
.C(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_293),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_35),
.B1(n_41),
.B2(n_9),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_254),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_272),
.B(n_247),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_294),
.B(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_246),
.C(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_282),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_265),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_300),
.Y(n_302)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_275),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_303),
.C(n_306),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_275),
.C(n_270),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_289),
.A2(n_256),
.B(n_284),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_305),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_279),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_10),
.B(n_15),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_285),
.B(n_33),
.C(n_37),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_311),
.C(n_312),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_12),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_33),
.C(n_37),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_12),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_298),
.B(n_292),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_316),
.B(n_320),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_295),
.B1(n_35),
.B2(n_8),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_13),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_310),
.B(n_15),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_321),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_308),
.A2(n_301),
.B1(n_312),
.B2(n_307),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_33),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_14),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_325),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_2),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_14),
.B(n_13),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_3),
.C(n_4),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_328),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_325),
.B(n_2),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_334),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_3),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_323),
.A2(n_3),
.B(n_4),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_316),
.B(n_5),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_338),
.B(n_330),
.C(n_327),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_341),
.Y(n_344)
);

O2A1O1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_332),
.A2(n_321),
.B(n_324),
.C(n_6),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_4),
.C(n_5),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_329),
.Y(n_342)
);

OAI311xp33_ASAP7_75t_L g345 ( 
.A1(n_342),
.A2(n_343),
.A3(n_340),
.B1(n_6),
.C1(n_7),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_344),
.B(n_6),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_346),
.B(n_5),
.C(n_7),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_5),
.B(n_7),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g349 ( 
.A(n_348),
.Y(n_349)
);


endmodule