module fake_jpeg_1144_n_131 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_131);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_12),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_35),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_42),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_61),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_37),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_70),
.Y(n_82)
);

OAI32xp33_ASAP7_75t_L g67 ( 
.A1(n_57),
.A2(n_32),
.A3(n_39),
.B1(n_33),
.B2(n_36),
.Y(n_67)
);

AO22x1_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_43),
.B1(n_36),
.B2(n_53),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_76),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_0),
.Y(n_81)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_89),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_69),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_88),
.B1(n_70),
.B2(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_3),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_92),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_19),
.C(n_28),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_98),
.C(n_21),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_79),
.B(n_5),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_6),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_80),
.C(n_87),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_103),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_17),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_97),
.B1(n_102),
.B2(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_112),
.B1(n_115),
.B2(n_94),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_15),
.C(n_24),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_16),
.B(n_27),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_119),
.A2(n_120),
.B1(n_113),
.B2(n_110),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_106),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_121),
.B(n_116),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_118),
.C(n_114),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_124),
.B(n_125),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_111),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_127),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_128),
.A2(n_122),
.B(n_105),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_129),
.A2(n_109),
.B(n_14),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_13),
.Y(n_131)
);


endmodule