module fake_jpeg_23192_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_7),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_39),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_18),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_27),
.B1(n_31),
.B2(n_18),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_46),
.B1(n_48),
.B2(n_38),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_31),
.B1(n_18),
.B2(n_28),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_43),
.B1(n_46),
.B2(n_48),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_39),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_58),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_76),
.B(n_78),
.Y(n_96)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_62),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_45),
.B1(n_48),
.B2(n_46),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_65),
.B1(n_75),
.B2(n_77),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_71),
.B1(n_41),
.B2(n_47),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_52),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_73),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_64),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_52),
.A2(n_42),
.B1(n_30),
.B2(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_66),
.B(n_67),
.Y(n_95)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_74),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_30),
.B1(n_19),
.B2(n_34),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_0),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_72),
.A2(n_34),
.B1(n_23),
.B2(n_29),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_33),
.C(n_25),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_37),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_41),
.B(n_37),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_87),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_59),
.A2(n_21),
.B(n_17),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_63),
.B(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_91),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_17),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_100),
.Y(n_111)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_20),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_20),
.B1(n_33),
.B2(n_49),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_74),
.B1(n_68),
.B2(n_57),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_49),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_70),
.Y(n_123)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_70),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_96),
.A2(n_56),
.B(n_60),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_96),
.B(n_81),
.Y(n_129)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_106),
.A2(n_110),
.B(n_125),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_102),
.B(n_72),
.C(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_120),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_61),
.B(n_75),
.C(n_33),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_67),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_112),
.B(n_119),
.C(n_93),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_82),
.B1(n_81),
.B2(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_90),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_118),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_55),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_83),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_126),
.Y(n_133)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_124),
.A2(n_104),
.B1(n_93),
.B2(n_91),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_49),
.B(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_1),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_97),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_88),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_142),
.B(n_110),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_134),
.B1(n_138),
.B2(n_152),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_87),
.B1(n_103),
.B2(n_82),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_137),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_82),
.B1(n_95),
.B2(n_85),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_140),
.B(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_105),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_147),
.Y(n_154)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_146),
.A2(n_118),
.B(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_85),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_115),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_125),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_110),
.A2(n_93),
.B1(n_89),
.B2(n_5),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_155),
.A2(n_156),
.B(n_159),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_142),
.A2(n_127),
.B(n_117),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_109),
.Y(n_157)
);

AOI21x1_ASAP7_75t_L g179 ( 
.A1(n_157),
.A2(n_156),
.B(n_160),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_110),
.B1(n_111),
.B2(n_106),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_173),
.B1(n_3),
.B2(n_4),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_139),
.B1(n_110),
.B2(n_152),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_138),
.B1(n_134),
.B2(n_139),
.Y(n_174)
);

AOI21xp33_ASAP7_75t_L g168 ( 
.A1(n_147),
.A2(n_130),
.B(n_148),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_172),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_154),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_133),
.B(n_126),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_132),
.A2(n_128),
.B1(n_4),
.B2(n_5),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_143),
.C(n_150),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_160),
.C(n_154),
.Y(n_189)
);

AO22x1_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_140),
.B1(n_145),
.B2(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_164),
.A2(n_136),
.B1(n_135),
.B2(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_185),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_163),
.B(n_6),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_162),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_158),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_197),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_165),
.C(n_171),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_192),
.A2(n_195),
.B(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_166),
.Y(n_194)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_165),
.C(n_181),
.Y(n_195)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_178),
.A2(n_179),
.B(n_157),
.C(n_181),
.D(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_182),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_200),
.A2(n_183),
.B1(n_185),
.B2(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_210),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_188),
.A2(n_157),
.B1(n_159),
.B2(n_158),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_173),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_206),
.B(n_193),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g208 ( 
.A(n_195),
.B(n_169),
.CI(n_180),
.CON(n_208),
.SN(n_208)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_208),
.B(n_197),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_169),
.B1(n_161),
.B2(n_10),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_198),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_207),
.C(n_203),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_189),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_215),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_213),
.B(n_161),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_205),
.C(n_209),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_219),
.A2(n_222),
.B1(n_210),
.B2(n_208),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_211),
.B(n_217),
.C(n_208),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_224),
.A3(n_226),
.B1(n_196),
.B2(n_9),
.C1(n_11),
.C2(n_12),
.Y(n_228)
);

AOI21x1_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_211),
.B(n_206),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_225),
.A2(n_8),
.B(n_11),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_8),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_14),
.B(n_12),
.Y(n_232)
);

NOR3xp33_ASAP7_75t_SL g233 ( 
.A(n_232),
.B(n_230),
.C(n_12),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_13),
.Y(n_234)
);


endmodule