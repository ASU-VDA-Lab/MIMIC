module fake_ariane_1549_n_62 (n_8, n_7, n_22, n_1, n_6, n_13, n_20, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_62);

input n_8;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;

output n_62;

wire n_56;
wire n_60;
wire n_24;
wire n_43;
wire n_49;
wire n_27;
wire n_48;
wire n_29;
wire n_41;
wire n_50;
wire n_38;
wire n_55;
wire n_47;
wire n_32;
wire n_28;
wire n_37;
wire n_58;
wire n_51;
wire n_45;
wire n_34;
wire n_26;
wire n_46;
wire n_52;
wire n_36;
wire n_33;
wire n_44;
wire n_30;
wire n_40;
wire n_39;
wire n_59;
wire n_31;
wire n_42;
wire n_57;
wire n_53;
wire n_61;
wire n_35;
wire n_54;
wire n_25;

INVx5_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_6),
.B(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_R g39 ( 
.A(n_37),
.B(n_32),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_3),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_22),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_34),
.B1(n_27),
.B2(n_33),
.Y(n_46)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_27),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_35),
.B(n_25),
.C(n_24),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_36),
.Y(n_49)
);

OR2x6_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_43),
.Y(n_51)
);

NAND4xp25_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_41),
.C(n_39),
.D(n_45),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_48),
.Y(n_53)
);

AOI211x1_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_45),
.B(n_24),
.C(n_36),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_24),
.Y(n_56)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_24),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_R g58 ( 
.A(n_56),
.B(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

AO22x2_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_4),
.B1(n_7),
.B2(n_9),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_58),
.A3(n_12),
.B1(n_14),
.B2(n_16),
.C1(n_21),
.C2(n_10),
.Y(n_62)
);


endmodule