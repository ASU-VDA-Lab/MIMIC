module fake_ariane_260_n_186 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_186);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_186;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_30;
wire n_82;
wire n_178;
wire n_42;
wire n_31;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_101;
wire n_94;
wire n_134;
wire n_185;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_28),
.Y(n_31)
);

INVxp67_ASAP7_75t_SL g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_0),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

AND2x4_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_34),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_71),
.B(n_31),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_46),
.B1(n_50),
.B2(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_50),
.B1(n_5),
.B2(n_6),
.Y(n_78)
);

NOR2xp67_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_43),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_60),
.Y(n_81)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_7),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_85)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_19),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_66),
.B(n_61),
.C(n_58),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

OR2x6_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_62),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_73),
.A2(n_54),
.B1(n_56),
.B2(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_R g95 ( 
.A(n_88),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_66),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_87),
.B(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_68),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_99),
.A2(n_80),
.B(n_89),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_63),
.B(n_57),
.Y(n_103)
);

HB1xp67_ASAP7_75t_SL g104 ( 
.A(n_96),
.Y(n_104)
);

O2A1O1Ixp5_ASAP7_75t_L g105 ( 
.A1(n_100),
.A2(n_68),
.B(n_59),
.C(n_52),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_78),
.B1(n_74),
.B2(n_86),
.Y(n_106)
);

AND2x4_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_63),
.Y(n_107)
);

OA21x2_ASAP7_75t_L g108 ( 
.A1(n_101),
.A2(n_57),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_83),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_98),
.Y(n_111)
);

OR2x6_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_92),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_90),
.B(n_93),
.C(n_52),
.Y(n_113)
);

NOR2x1_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_92),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_76),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_107),
.Y(n_120)
);

OA21x2_ASAP7_75t_L g121 ( 
.A1(n_113),
.A2(n_102),
.B(n_105),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_115),
.Y(n_123)
);

AND4x1_ASAP7_75t_L g124 ( 
.A(n_120),
.B(n_90),
.C(n_82),
.D(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_83),
.C(n_67),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

OAI21x1_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_102),
.B(n_103),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_82),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_59),
.B(n_52),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_134),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_125),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

NOR2xp67_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_127),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_142),
.B(n_126),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_126),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_112),
.Y(n_159)
);

NOR2x1p5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_158),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_141),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_145),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_153),
.B(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_59),
.C(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_155),
.Y(n_170)
);

AND2x4_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_153),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_152),
.Y(n_172)
);

AOI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_161),
.A2(n_159),
.B(n_85),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_164),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_86),
.B1(n_112),
.B2(n_156),
.Y(n_175)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_167),
.A2(n_74),
.B1(n_156),
.B2(n_157),
.C(n_124),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_170),
.A2(n_165),
.B1(n_166),
.B2(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

OAI221xp5_ASAP7_75t_L g180 ( 
.A1(n_175),
.A2(n_112),
.B1(n_132),
.B2(n_97),
.C(n_94),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_177),
.A2(n_176),
.B1(n_174),
.B2(n_171),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_180),
.A2(n_173),
.B1(n_108),
.B2(n_103),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_178),
.A2(n_108),
.B1(n_94),
.B2(n_97),
.Y(n_183)
);

NAND4xp25_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_179),
.C(n_95),
.D(n_25),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_181),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_185),
.A2(n_182),
.B1(n_108),
.B2(n_103),
.Y(n_186)
);


endmodule