module fake_jpeg_27847_n_173 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_12),
.Y(n_42)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_27),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_16),
.B1(n_23),
.B2(n_18),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_28),
.B1(n_17),
.B2(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_44),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_19),
.B(n_23),
.C(n_18),
.Y(n_44)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_29),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_30),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_47),
.B(n_57),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_16),
.B1(n_19),
.B2(n_28),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_50),
.B1(n_31),
.B2(n_32),
.Y(n_84)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_55),
.Y(n_66)
);

OR2x4_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_29),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_25),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_26),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_63),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_60),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_27),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_32),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_25),
.C(n_27),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_50),
.B1(n_45),
.B2(n_53),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_65),
.A2(n_75),
.B1(n_84),
.B2(n_33),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_78),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_32),
.C(n_25),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_60),
.C(n_24),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_76),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g77 ( 
.A1(n_49),
.A2(n_31),
.B(n_27),
.C(n_25),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_33),
.B(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_12),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_15),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_15),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_62),
.A2(n_31),
.B1(n_17),
.B2(n_33),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_51),
.B1(n_17),
.B2(n_56),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_96),
.C(n_77),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_102),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_97),
.B1(n_79),
.B2(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_94),
.B(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_33),
.C(n_56),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_24),
.B1(n_21),
.B2(n_13),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_106),
.B1(n_13),
.B2(n_2),
.Y(n_122)
);

CKINVDCx12_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_22),
.B(n_21),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_107),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_65),
.A2(n_59),
.B1(n_21),
.B2(n_24),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_0),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_81),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_116),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_74),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_77),
.B1(n_67),
.B2(n_72),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_121),
.B1(n_122),
.B2(n_90),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_77),
.B1(n_80),
.B2(n_83),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_120),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_92),
.Y(n_119)
);

AO221x1_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_89),
.B1(n_103),
.B2(n_104),
.C(n_106),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_13),
.B1(n_2),
.B2(n_3),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_130),
.B(n_118),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_105),
.B(n_102),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_121),
.B(n_108),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_98),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_133),
.B(n_135),
.C(n_109),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_98),
.C(n_96),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_143),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_114),
.C(n_109),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_142),
.C(n_144),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_117),
.C(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_115),
.C(n_11),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_141),
.A2(n_134),
.B(n_129),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_148),
.B(n_146),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_133),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_5),
.Y(n_159)
);

FAx1_ASAP7_75t_SL g151 ( 
.A(n_140),
.B(n_128),
.CI(n_129),
.CON(n_151),
.SN(n_151)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_151),
.B(n_11),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_153),
.B(n_5),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_155),
.A2(n_158),
.B1(n_160),
.B2(n_150),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_10),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_149),
.B(n_1),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_147),
.A2(n_1),
.B(n_4),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_152),
.C(n_147),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_161),
.B(n_160),
.C(n_6),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_164),
.B(n_165),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_159),
.A2(n_151),
.B1(n_150),
.B2(n_152),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_167),
.A2(n_168),
.B(n_163),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_5),
.C(n_6),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_166),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_162),
.C(n_170),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_7),
.Y(n_173)
);


endmodule