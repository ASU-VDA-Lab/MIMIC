module fake_jpeg_24332_n_288 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_288);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_1),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_13),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_23),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_56),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_36),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_63),
.B1(n_65),
.B2(n_78),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_36),
.B1(n_19),
.B2(n_23),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_58),
.B1(n_19),
.B2(n_17),
.Y(n_109)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_57),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_33),
.Y(n_55)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_30),
.B1(n_36),
.B2(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_35),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_59),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_60),
.B(n_66),
.Y(n_87)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_61),
.B(n_69),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_29),
.B1(n_35),
.B2(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_34),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_68),
.B(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_74),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_34),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_32),
.B(n_27),
.Y(n_75)
);

OR2x2_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_76),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_2),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_26),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_16),
.C(n_15),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_32),
.B1(n_17),
.B2(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_81),
.Y(n_103)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_20),
.B1(n_25),
.B2(n_18),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_20),
.B(n_25),
.C(n_18),
.Y(n_101)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_97),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_104),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_76),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_67),
.C(n_79),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_22),
.B1(n_31),
.B2(n_21),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_102),
.B1(n_110),
.B2(n_82),
.Y(n_137)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_72),
.B1(n_64),
.B2(n_62),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_22),
.B1(n_31),
.B2(n_19),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_22),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_108),
.Y(n_123)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_112),
.B1(n_69),
.B2(n_5),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g110 ( 
.A1(n_70),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_70),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_74),
.Y(n_128)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_119),
.Y(n_131)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_121),
.B(n_128),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_126),
.C(n_93),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_86),
.C(n_85),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_94),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_127),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_137),
.B1(n_93),
.B2(n_102),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_132),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_88),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_135),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_15),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_136),
.B(n_139),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_82),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_109),
.Y(n_160)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_91),
.B(n_3),
.Y(n_142)
);

NAND2x1_ASAP7_75t_SL g162 ( 
.A(n_142),
.B(n_149),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_5),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_143),
.Y(n_172)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_97),
.B1(n_89),
.B2(n_110),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_72),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_151),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_5),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_100),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_161),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_158),
.B1(n_165),
.B2(n_135),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_148),
.B(n_136),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_157),
.A2(n_159),
.B(n_168),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_102),
.B1(n_96),
.B2(n_92),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_118),
.B(n_103),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_160),
.B(n_147),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_100),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_144),
.A2(n_106),
.B(n_107),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_64),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_6),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_6),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_128),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_181),
.Y(n_200)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_142),
.B(n_6),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_182),
.A2(n_151),
.B(n_131),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_185),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_187),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_180),
.B(n_140),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_188),
.B(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_149),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_190),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_192),
.B(n_196),
.Y(n_213)
);

OA21x2_ASAP7_75t_L g193 ( 
.A1(n_164),
.A2(n_130),
.B(n_127),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_154),
.B(n_169),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_178),
.B(n_163),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_197),
.B(n_202),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_201),
.B1(n_206),
.B2(n_162),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_168),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_160),
.B(n_133),
.Y(n_205)
);

OAI321xp33_ASAP7_75t_L g209 ( 
.A1(n_205),
.A2(n_162),
.A3(n_182),
.B1(n_172),
.B2(n_158),
.C(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

OA21x2_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_164),
.B(n_157),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_214),
.Y(n_241)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_161),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_215),
.C(n_204),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_152),
.C(n_181),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_219),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_175),
.B1(n_173),
.B2(n_121),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_132),
.B1(n_153),
.B2(n_154),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_222),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_206),
.A2(n_169),
.B1(n_145),
.B2(n_155),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_218),
.B(n_191),
.CI(n_184),
.CON(n_228),
.SN(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_203),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_201),
.C(n_186),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_204),
.C(n_184),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_196),
.C(n_194),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_225),
.C(n_187),
.Y(n_256)
);

NOR2x1_ASAP7_75t_R g237 ( 
.A(n_223),
.B(n_193),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_223),
.B(n_218),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_200),
.Y(n_238)
);

NOR2xp67_ASAP7_75t_SL g243 ( 
.A(n_231),
.B(n_219),
.Y(n_243)
);

NOR2xp67_ASAP7_75t_SL g266 ( 
.A(n_243),
.B(n_228),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_213),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_230),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_221),
.B1(n_208),
.B2(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_254),
.B1(n_255),
.B2(n_237),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_195),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_250),
.B(n_252),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_234),
.B(n_207),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_224),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_233),
.A2(n_208),
.B1(n_207),
.B2(n_214),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_242),
.A2(n_239),
.B1(n_240),
.B2(n_235),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_232),
.C(n_188),
.Y(n_264)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_257),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_249),
.B1(n_246),
.B2(n_255),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_261),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_205),
.B(n_197),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_271)
);

NAND4xp25_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_192),
.C(n_183),
.D(n_226),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_265),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_245),
.B(n_200),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_248),
.C(n_244),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_248),
.C(n_244),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_261),
.B1(n_256),
.B2(n_264),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g269 ( 
.A(n_258),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_275),
.B(n_277),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_267),
.C(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_210),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_272),
.B1(n_271),
.B2(n_262),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_279),
.B(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_281),
.B(n_282),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_273),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_SL g286 ( 
.A(n_284),
.B(n_285),
.C(n_228),
.Y(n_286)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_247),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g287 ( 
.A(n_286),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_283),
.Y(n_288)
);


endmodule