module fake_jpeg_662_n_11 (n_3, n_2, n_1, n_0, n_4, n_11);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_11;

wire n_10;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

XNOR2xp5_ASAP7_75t_L g5 ( 
.A(n_1),
.B(n_0),
.Y(n_5)
);

XOR2xp5_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_1),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_3),
.B(n_2),
.Y(n_7)
);

MAJx2_ASAP7_75t_L g8 ( 
.A(n_6),
.B(n_0),
.C(n_2),
.Y(n_8)
);

OAI22xp5_ASAP7_75t_L g10 ( 
.A1(n_8),
.A2(n_9),
.B1(n_7),
.B2(n_6),
.Y(n_10)
);

A2O1A1Ixp33_ASAP7_75t_SL g9 ( 
.A1(n_6),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_9)
);

FAx1_ASAP7_75t_SL g11 ( 
.A(n_10),
.B(n_8),
.CI(n_9),
.CON(n_11),
.SN(n_11)
);


endmodule