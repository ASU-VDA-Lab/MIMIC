module fake_netlist_1_5768_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
XNOR2xp5_ASAP7_75t_L g14 ( .A(n_0), .B(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_12), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
INVx6_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_14), .B1(n_13), .B2(n_15), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_18), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_14), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
OAI21xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_10), .B(n_17), .Y(n_26) );
NOR4xp25_ASAP7_75t_L g27 ( .A(n_25), .B(n_13), .C(n_12), .D(n_11), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_25), .A2(n_19), .B1(n_11), .B2(n_10), .Y(n_28) );
NAND4xp75_ASAP7_75t_L g29 ( .A(n_26), .B(n_0), .C(n_1), .D(n_2), .Y(n_29) );
XOR2xp5_ASAP7_75t_L g30 ( .A(n_28), .B(n_2), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_27), .B(n_3), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g33 ( .A(n_30), .B(n_27), .Y(n_33) );
AOI22xp5_ASAP7_75t_SL g34 ( .A1(n_33), .A2(n_29), .B1(n_4), .B2(n_5), .Y(n_34) );
OA331x2_ASAP7_75t_L g35 ( .A1(n_34), .A2(n_3), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_32), .C1(n_9), .Y(n_35) );
endmodule