module fake_jpeg_29314_n_403 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_403);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_403;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_11),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_67),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_61),
.Y(n_113)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_62),
.Y(n_120)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_63),
.Y(n_122)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_27),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_21),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_74),
.Y(n_107)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_49),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_36),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_81),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_46),
.B(n_11),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_40),
.B1(n_49),
.B2(n_47),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_102),
.B1(n_61),
.B2(n_78),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_84),
.B1(n_83),
.B2(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_48),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_124),
.Y(n_153)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_119),
.Y(n_160)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_125),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_107),
.A2(n_88),
.A3(n_103),
.B1(n_99),
.B2(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_129),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_113),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_128),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_88),
.B(n_54),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_152),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_43),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_134),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_30),
.B(n_39),
.C(n_31),
.Y(n_134)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_136),
.A2(n_121),
.B1(n_118),
.B2(n_47),
.Y(n_174)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_86),
.A2(n_39),
.B(n_26),
.C(n_30),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_159),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_98),
.A2(n_77),
.B1(n_59),
.B2(n_79),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_146),
.A2(n_149),
.B1(n_128),
.B2(n_70),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_92),
.A2(n_61),
.B1(n_66),
.B2(n_73),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_97),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_94),
.A2(n_34),
.B1(n_22),
.B2(n_47),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_151),
.A2(n_158),
.B1(n_47),
.B2(n_25),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_70),
.B(n_32),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_159),
.C(n_131),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_96),
.A2(n_33),
.B1(n_41),
.B2(n_22),
.Y(n_155)
);

NOR2x1_ASAP7_75t_R g171 ( 
.A(n_155),
.B(n_87),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_119),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_87),
.C(n_34),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_22),
.B1(n_34),
.B2(n_25),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_32),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_153),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_129),
.B1(n_160),
.B2(n_115),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_58),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_173),
.A2(n_174),
.B1(n_180),
.B2(n_146),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_175),
.A2(n_138),
.B1(n_140),
.B2(n_154),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_141),
.A2(n_121),
.B1(n_126),
.B2(n_97),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_184),
.A2(n_156),
.B(n_157),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_127),
.A2(n_109),
.B1(n_117),
.B2(n_122),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_128),
.B1(n_122),
.B2(n_137),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_106),
.C(n_111),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_155),
.C(n_133),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_192),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_197),
.B(n_208),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_184),
.B(n_161),
.C(n_157),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_202),
.B1(n_208),
.B2(n_197),
.Y(n_222)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_171),
.A2(n_150),
.B1(n_145),
.B2(n_117),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_164),
.B1(n_183),
.B2(n_174),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_181),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_144),
.B1(n_147),
.B2(n_142),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_186),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_206),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_163),
.B(n_134),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_164),
.B(n_154),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_208),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_149),
.B(n_143),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_209),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_206),
.A2(n_188),
.B(n_179),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_205),
.B(n_165),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_215),
.B(n_218),
.Y(n_251)
);

BUFx24_ASAP7_75t_L g217 ( 
.A(n_194),
.Y(n_217)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_198),
.A2(n_167),
.B1(n_176),
.B2(n_181),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_168),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_130),
.C(n_178),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_199),
.B1(n_202),
.B2(n_201),
.Y(n_243)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_132),
.B1(n_169),
.B2(n_185),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_202),
.B1(n_193),
.B2(n_203),
.Y(n_238)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_162),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_168),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_229),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_170),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_189),
.B(n_170),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_203),
.B1(n_190),
.B2(n_182),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_234),
.A2(n_41),
.B(n_57),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_191),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_227),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_236),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_243),
.B1(n_255),
.B2(n_225),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_224),
.A2(n_209),
.B(n_192),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_239),
.A2(n_226),
.B(n_229),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_196),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_242),
.C(n_246),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_195),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_215),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_191),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_210),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_200),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_247),
.B(n_250),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_162),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_219),
.B(n_178),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_252),
.B(n_48),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.C(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_166),
.C(n_130),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_185),
.B1(n_182),
.B2(n_148),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_256),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_237),
.A2(n_222),
.B1(n_230),
.B2(n_212),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_258),
.A2(n_272),
.B1(n_273),
.B2(n_283),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_232),
.A2(n_251),
.B(n_237),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_263),
.B(n_274),
.C(n_275),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_232),
.A2(n_214),
.B(n_223),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_258),
.B(n_276),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_216),
.C(n_213),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_266),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_251),
.A2(n_239),
.B(n_247),
.Y(n_266)
);

AOI22x1_ASAP7_75t_L g273 ( 
.A1(n_238),
.A2(n_216),
.B1(n_217),
.B2(n_135),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_217),
.C(n_120),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_217),
.C(n_91),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_255),
.B1(n_110),
.B2(n_249),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_257),
.A2(n_60),
.B(n_43),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_278),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_236),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_26),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_233),
.A2(n_50),
.B(n_69),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_281),
.B(n_46),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_241),
.B(n_50),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_243),
.A2(n_68),
.B1(n_56),
.B2(n_72),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_284),
.A2(n_287),
.B1(n_294),
.B2(n_302),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_287),
.B(n_286),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_264),
.A2(n_280),
.B1(n_279),
.B2(n_273),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_250),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_296),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_280),
.B(n_233),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_290),
.B(n_307),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_253),
.C(n_254),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_293),
.C(n_275),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_259),
.B(n_246),
.C(n_256),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_273),
.A2(n_245),
.B1(n_244),
.B2(n_248),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_295),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_248),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_259),
.B(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_260),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_272),
.A2(n_25),
.B1(n_75),
.B2(n_45),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_301),
.A2(n_292),
.B1(n_299),
.B2(n_300),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_14),
.B1(n_20),
.B2(n_19),
.Y(n_302)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_305),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_278),
.B(n_14),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_311),
.B1(n_313),
.B2(n_319),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_318),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_310),
.B(n_303),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_267),
.B1(n_270),
.B2(n_269),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_312),
.A2(n_9),
.B(n_18),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_261),
.B1(n_266),
.B2(n_283),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_291),
.C(n_289),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_324),
.C(n_325),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_262),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_38),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_281),
.C(n_277),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_282),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_31),
.C(n_58),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_326),
.B(n_327),
.C(n_284),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_300),
.B(n_65),
.C(n_36),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_298),
.B(n_12),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_328),
.B(n_14),
.Y(n_337)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_310),
.Y(n_333)
);

INVx11_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_322),
.B(n_302),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_334),
.B(n_335),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_336),
.B(n_340),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_339),
.Y(n_355)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_294),
.B1(n_301),
.B2(n_2),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_329),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_314),
.B(n_10),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_308),
.A2(n_10),
.B1(n_20),
.B2(n_19),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_9),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_36),
.C(n_38),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_343),
.B(n_309),
.C(n_318),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_344),
.A2(n_18),
.B(n_16),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_9),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_18),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_335),
.A2(n_317),
.B(n_324),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_38),
.B(n_13),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_348),
.B(n_354),
.Y(n_369)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_349),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_338),
.A2(n_326),
.B1(n_327),
.B2(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_350),
.B(n_351),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_320),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_331),
.B(n_320),
.C(n_325),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_330),
.C(n_336),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_358),
.B(n_332),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_SL g362 ( 
.A(n_351),
.B(n_333),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_362),
.B(n_365),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_368),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_330),
.C(n_343),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_371),
.Y(n_377)
);

NOR2xp67_ASAP7_75t_SL g365 ( 
.A(n_359),
.B(n_344),
.Y(n_365)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_366),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_356),
.A2(n_16),
.B(n_15),
.Y(n_367)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_346),
.A2(n_38),
.B1(n_16),
.B2(n_15),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_357),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_347),
.C(n_349),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_363),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_375),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_360),
.B(n_359),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_378),
.A2(n_381),
.B(n_382),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_361),
.A2(n_353),
.B(n_350),
.Y(n_379)
);

OAI21x1_ASAP7_75t_SL g390 ( 
.A1(n_379),
.A2(n_36),
.B(n_5),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_369),
.A2(n_349),
.B(n_355),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_354),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_377),
.A2(n_364),
.B(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_384),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_376),
.A2(n_13),
.B(n_1),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_385),
.B(n_389),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_372),
.A2(n_13),
.B1(n_1),
.B2(n_2),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_388),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_36),
.C(n_1),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_378),
.A2(n_0),
.B(n_2),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_390),
.A2(n_375),
.B(n_373),
.Y(n_391)
);

AO21x2_ASAP7_75t_L g397 ( 
.A1(n_391),
.A2(n_395),
.B(n_36),
.Y(n_397)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_383),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_392),
.A2(n_386),
.B(n_5),
.Y(n_396)
);

AO21x1_ASAP7_75t_L g399 ( 
.A1(n_396),
.A2(n_397),
.B(n_398),
.Y(n_399)
);

OAI311xp33_ASAP7_75t_L g398 ( 
.A1(n_394),
.A2(n_0),
.A3(n_6),
.B1(n_7),
.C1(n_8),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_396),
.A2(n_393),
.B(n_6),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_0),
.C(n_6),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_401),
.B(n_399),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_7),
.C(n_8),
.Y(n_403)
);


endmodule