module fake_netlist_1_11055_n_907 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_204, n_221, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_237, n_181, n_101, n_62, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_242, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_191, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_224, n_96, n_225, n_39, n_907);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_204;
input n_221;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_237;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_242;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_224;
input n_96;
input n_225;
input n_39;
output n_907;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_903;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_857;
wire n_786;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_466;
wire n_302;
wire n_900;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_446;
wire n_420;
wire n_285;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_880;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_898;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_409;
wire n_363;
wire n_315;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_267;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_819;
wire n_290;
wire n_405;
wire n_772;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g244 ( .A(n_85), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_238), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_107), .Y(n_246) );
NOR2xp67_ASAP7_75t_L g247 ( .A(n_214), .B(n_126), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_242), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_27), .Y(n_249) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_172), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_38), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_231), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_157), .Y(n_253) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_65), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_147), .Y(n_255) );
CKINVDCx5p33_ASAP7_75t_R g256 ( .A(n_110), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_202), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_74), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_55), .Y(n_259) );
CKINVDCx14_ASAP7_75t_R g260 ( .A(n_166), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_182), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_75), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_200), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_62), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_125), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_103), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_139), .Y(n_267) );
CKINVDCx5p33_ASAP7_75t_R g268 ( .A(n_81), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_9), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_191), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_152), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_120), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_115), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_212), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_57), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_9), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g277 ( .A(n_1), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_197), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_150), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_91), .Y(n_280) );
CKINVDCx20_ASAP7_75t_R g281 ( .A(n_39), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_30), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_95), .Y(n_283) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_168), .Y(n_284) );
CKINVDCx5p33_ASAP7_75t_R g285 ( .A(n_138), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_241), .B(n_101), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_34), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_117), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_144), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_43), .Y(n_290) );
CKINVDCx16_ASAP7_75t_R g291 ( .A(n_72), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_173), .Y(n_292) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_52), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_105), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_89), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_155), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_1), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_183), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_169), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_25), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_132), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_206), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_171), .Y(n_303) );
CKINVDCx5p33_ASAP7_75t_R g304 ( .A(n_102), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_78), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_31), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_22), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_161), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_127), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_36), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_228), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_195), .Y(n_313) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_154), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_179), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_109), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_104), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_187), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_2), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_188), .B(n_220), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_45), .B(n_106), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_6), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_177), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_239), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_203), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_60), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_237), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_128), .Y(n_328) );
BUFx8_ASAP7_75t_SL g329 ( .A(n_46), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_88), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_67), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_186), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_87), .Y(n_333) );
BUFx10_ASAP7_75t_L g334 ( .A(n_233), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_13), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_234), .Y(n_336) );
CKINVDCx5p33_ASAP7_75t_R g337 ( .A(n_73), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_59), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_71), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_164), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_63), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_170), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_44), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_194), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_178), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_97), .Y(n_346) );
BUFx8_ASAP7_75t_SL g347 ( .A(n_70), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_180), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_209), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_11), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_111), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_32), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_199), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_113), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_19), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g356 ( .A(n_222), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_137), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_47), .Y(n_358) );
BUFx8_ASAP7_75t_SL g359 ( .A(n_198), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_15), .Y(n_360) );
CKINVDCx14_ASAP7_75t_R g361 ( .A(n_42), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_25), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_174), .Y(n_363) );
CKINVDCx5p33_ASAP7_75t_R g364 ( .A(n_131), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_18), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g366 ( .A(n_226), .Y(n_366) );
NOR2xp67_ASAP7_75t_L g367 ( .A(n_13), .B(n_230), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_335), .B(n_0), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_257), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_246), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_244), .A2(n_28), .B(n_26), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_255), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_249), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_350), .Y(n_374) );
BUFx3_ASAP7_75t_L g375 ( .A(n_289), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_269), .B(n_0), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_272), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_360), .B(n_3), .Y(n_378) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_270), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_258), .A2(n_33), .B(n_29), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_305), .Y(n_381) );
INVx3_ASAP7_75t_L g382 ( .A(n_276), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_270), .Y(n_383) );
AND2x6_ASAP7_75t_L g384 ( .A(n_324), .B(n_35), .Y(n_384) );
BUFx6f_ASAP7_75t_L g385 ( .A(n_270), .Y(n_385) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_259), .A2(n_40), .B(n_37), .Y(n_386) );
BUFx12f_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
INVxp67_ASAP7_75t_L g388 ( .A(n_297), .Y(n_388) );
OAI22x1_ASAP7_75t_R g389 ( .A1(n_245), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_389) );
BUFx6f_ASAP7_75t_L g390 ( .A(n_270), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_261), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_355), .B(n_4), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_262), .Y(n_393) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_282), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_282), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_276), .Y(n_396) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_282), .Y(n_397) );
INVx3_ASAP7_75t_L g398 ( .A(n_392), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_379), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_370), .B(n_253), .Y(n_400) );
INVx3_ASAP7_75t_L g401 ( .A(n_392), .Y(n_401) );
NOR2x1p5_ASAP7_75t_L g402 ( .A(n_387), .B(n_277), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
NAND2xp5_ASAP7_75t_SL g404 ( .A(n_388), .B(n_264), .Y(n_404) );
NAND2xp33_ASAP7_75t_L g405 ( .A(n_384), .B(n_282), .Y(n_405) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_369), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_379), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_368), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_368), .Y(n_409) );
INVx3_ASAP7_75t_L g410 ( .A(n_392), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
INVx3_ASAP7_75t_L g412 ( .A(n_378), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_379), .Y(n_413) );
NAND2xp33_ASAP7_75t_L g414 ( .A(n_384), .B(n_250), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_397), .Y(n_415) );
OA22x2_ASAP7_75t_L g416 ( .A1(n_378), .A2(n_308), .B1(n_319), .B2(n_300), .Y(n_416) );
INVx8_ASAP7_75t_L g417 ( .A(n_384), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_378), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_370), .B(n_291), .Y(n_419) );
AO21x2_ASAP7_75t_L g420 ( .A1(n_371), .A2(n_267), .B(n_265), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_373), .B(n_366), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_376), .B(n_365), .C(n_322), .Y(n_422) );
AND3x2_ASAP7_75t_L g423 ( .A(n_389), .B(n_311), .C(n_273), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_397), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_372), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_400), .B(n_373), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_425), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_412), .A2(n_391), .B1(n_393), .B2(n_384), .Y(n_428) );
NAND2xp5_ASAP7_75t_SL g429 ( .A(n_417), .B(n_371), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g430 ( .A1(n_403), .A2(n_374), .B1(n_393), .B2(n_391), .C(n_377), .Y(n_430) );
INVx8_ASAP7_75t_L g431 ( .A(n_417), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g433 ( .A(n_422), .B(n_372), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_406), .B(n_375), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_406), .B(n_384), .Y(n_435) );
INVx2_ASAP7_75t_SL g436 ( .A(n_412), .Y(n_436) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_408), .A2(n_381), .B(n_377), .C(n_361), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_409), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_418), .B(n_384), .Y(n_439) );
OAI22xp33_ASAP7_75t_L g440 ( .A1(n_416), .A2(n_248), .B1(n_281), .B2(n_254), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_416), .A2(n_284), .B1(n_312), .B2(n_293), .Y(n_441) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_417), .B(n_271), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_419), .B(n_381), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_398), .A2(n_260), .B1(n_361), .B2(n_276), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_398), .B(n_251), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_398), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_421), .B(n_404), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_401), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_401), .B(n_252), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_401), .Y(n_450) );
INVx2_ASAP7_75t_SL g451 ( .A(n_410), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_410), .B(n_256), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_414), .A2(n_362), .B1(n_276), .B2(n_274), .Y(n_453) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_405), .A2(n_275), .B(n_287), .C(n_278), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_420), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_414), .A2(n_367), .B1(n_292), .B2(n_296), .C(n_341), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_405), .B(n_263), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
AND2x4_ASAP7_75t_L g459 ( .A(n_402), .B(n_314), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_438), .A2(n_363), .B1(n_351), .B2(n_362), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_426), .A2(n_362), .B1(n_303), .B2(n_306), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_441), .B(n_420), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_426), .B(n_266), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_431), .B(n_268), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_L g465 ( .A1(n_432), .A2(n_307), .B(n_310), .C(n_288), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_439), .A2(n_386), .B(n_380), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_446), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_447), .B(n_423), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_450), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_440), .A2(n_316), .B(n_317), .C(n_315), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_429), .A2(n_386), .B(n_380), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_448), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_440), .A2(n_326), .B(n_327), .C(n_318), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_455), .A2(n_338), .B(n_332), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_435), .A2(n_340), .B(n_339), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_458), .A2(n_343), .B(n_342), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_428), .A2(n_346), .B(n_344), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_447), .B(n_334), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_431), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_442), .A2(n_349), .B(n_348), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_459), .B(n_301), .C(n_299), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_443), .B(n_427), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_442), .A2(n_358), .B(n_354), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_434), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_443), .B(n_279), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_444), .B(n_280), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
AND3x2_ASAP7_75t_L g488 ( .A(n_459), .B(n_347), .C(n_329), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_433), .B(n_283), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_451), .B(n_285), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_445), .A2(n_407), .B(n_399), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_456), .A2(n_345), .B(n_396), .C(n_382), .Y(n_492) );
NAND2xp33_ASAP7_75t_L g493 ( .A(n_431), .B(n_290), .Y(n_493) );
NOR2xp33_ASAP7_75t_SL g494 ( .A(n_454), .B(n_359), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_437), .A2(n_247), .B(n_286), .C(n_320), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_467), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_474), .A2(n_476), .B(n_475), .Y(n_497) );
INVx5_ASAP7_75t_L g498 ( .A(n_479), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_460), .B(n_449), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_474), .A2(n_453), .B(n_452), .Y(n_500) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_471), .A2(n_457), .B(n_430), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_468), .B(n_294), .Y(n_502) );
OAI21x1_ASAP7_75t_SL g503 ( .A1(n_477), .A2(n_5), .B(n_7), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_471), .A2(n_321), .B(n_320), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_479), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_466), .A2(n_413), .B(n_411), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_478), .B(n_362), .Y(n_507) );
OR2x6_ASAP7_75t_L g508 ( .A(n_470), .B(n_473), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_482), .A2(n_424), .B(n_415), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_472), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_492), .A2(n_382), .B(n_396), .C(n_385), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_491), .A2(n_424), .B(n_415), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_495), .A2(n_413), .B(n_298), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_484), .B(n_295), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_481), .B(n_7), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_462), .B(n_465), .Y(n_516) );
AOI21x1_ASAP7_75t_L g517 ( .A1(n_477), .A2(n_385), .B(n_383), .Y(n_517) );
AO22x2_ASAP7_75t_L g518 ( .A1(n_461), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_518) );
AO31x2_ASAP7_75t_L g519 ( .A1(n_480), .A2(n_397), .A3(n_395), .B(n_394), .Y(n_519) );
INVx2_ASAP7_75t_SL g520 ( .A(n_488), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_485), .A2(n_304), .B(n_302), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_463), .A2(n_313), .B(n_309), .Y(n_522) );
OA22x2_ASAP7_75t_L g523 ( .A1(n_487), .A2(n_357), .B1(n_323), .B2(n_325), .Y(n_523) );
OAI21x1_ASAP7_75t_L g524 ( .A1(n_483), .A2(n_48), .B(n_41), .Y(n_524) );
INVx3_ASAP7_75t_L g525 ( .A(n_490), .Y(n_525) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_486), .A2(n_330), .B(n_328), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_493), .B(n_331), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_464), .B(n_333), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_489), .Y(n_529) );
OAI21x1_ASAP7_75t_L g530 ( .A1(n_494), .A2(n_50), .B(n_49), .Y(n_530) );
NOR2xp67_ASAP7_75t_L g531 ( .A(n_460), .B(n_8), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_469), .Y(n_532) );
INVx2_ASAP7_75t_SL g533 ( .A(n_488), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_484), .B(n_336), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_479), .B(n_10), .Y(n_535) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_517), .A2(n_385), .B(n_383), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g537 ( .A1(n_511), .A2(n_148), .B(n_243), .C(n_240), .Y(n_537) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_504), .A2(n_352), .B(n_337), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_508), .A2(n_397), .B1(n_395), .B2(n_394), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_516), .A2(n_364), .B1(n_356), .B2(n_353), .Y(n_540) );
INVx3_ASAP7_75t_L g541 ( .A(n_505), .Y(n_541) );
AO21x2_ASAP7_75t_L g542 ( .A1(n_513), .A2(n_395), .B(n_394), .Y(n_542) );
OAI21x1_ASAP7_75t_L g543 ( .A1(n_512), .A2(n_395), .B(n_394), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_515), .B(n_12), .Y(n_544) );
OAI21x1_ASAP7_75t_L g545 ( .A1(n_501), .A2(n_390), .B(n_140), .Y(n_545) );
NAND2x1p5_ASAP7_75t_L g546 ( .A(n_498), .B(n_12), .Y(n_546) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_531), .A2(n_497), .B(n_500), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_496), .Y(n_548) );
INVxp33_ASAP7_75t_L g549 ( .A(n_514), .Y(n_549) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_505), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_503), .A2(n_390), .B(n_141), .Y(n_552) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_524), .A2(n_390), .B(n_142), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_508), .B(n_14), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_510), .Y(n_555) );
OAI21x1_ASAP7_75t_L g556 ( .A1(n_509), .A2(n_136), .B(n_236), .Y(n_556) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_520), .Y(n_557) );
OAI21xp5_ASAP7_75t_L g558 ( .A1(n_510), .A2(n_15), .B(n_16), .Y(n_558) );
OAI21x1_ASAP7_75t_L g559 ( .A1(n_530), .A2(n_143), .B(n_235), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_533), .Y(n_560) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_532), .A2(n_135), .B(n_229), .Y(n_561) );
BUFx3_ASAP7_75t_L g562 ( .A(n_498), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_529), .B(n_16), .Y(n_563) );
OA21x2_ASAP7_75t_L g564 ( .A1(n_507), .A2(n_134), .B(n_227), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_505), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_534), .B(n_17), .Y(n_567) );
NAND2x1p5_ASAP7_75t_L g568 ( .A(n_525), .B(n_17), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_535), .B(n_18), .Y(n_569) );
BUFx3_ASAP7_75t_L g570 ( .A(n_523), .Y(n_570) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_499), .A2(n_145), .B(n_225), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_526), .A2(n_19), .B(n_20), .Y(n_573) );
OAI21x1_ASAP7_75t_L g574 ( .A1(n_521), .A2(n_146), .B(n_224), .Y(n_574) );
CKINVDCx11_ASAP7_75t_R g575 ( .A(n_518), .Y(n_575) );
OAI21x1_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_133), .B(n_223), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_518), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_519), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_528), .Y(n_579) );
AO21x2_ASAP7_75t_L g580 ( .A1(n_527), .A2(n_130), .B(n_221), .Y(n_580) );
OAI21x1_ASAP7_75t_L g581 ( .A1(n_522), .A2(n_129), .B(n_219), .Y(n_581) );
AO21x2_ASAP7_75t_L g582 ( .A1(n_502), .A2(n_124), .B(n_218), .Y(n_582) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_518), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_583) );
OAI21x1_ASAP7_75t_L g584 ( .A1(n_517), .A2(n_149), .B(n_217), .Y(n_584) );
BUFx2_ASAP7_75t_L g585 ( .A(n_535), .Y(n_585) );
AND2x4_ASAP7_75t_L g586 ( .A(n_525), .B(n_21), .Y(n_586) );
OAI21x1_ASAP7_75t_L g587 ( .A1(n_517), .A2(n_123), .B(n_216), .Y(n_587) );
CKINVDCx20_ASAP7_75t_R g588 ( .A(n_520), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_496), .B(n_23), .Y(n_589) );
OAI21x1_ASAP7_75t_L g590 ( .A1(n_517), .A2(n_122), .B(n_215), .Y(n_590) );
AO21x1_ASAP7_75t_L g591 ( .A1(n_504), .A2(n_23), .B(n_24), .Y(n_591) );
OAI21x1_ASAP7_75t_SL g592 ( .A1(n_503), .A2(n_24), .B(n_51), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_506), .A2(n_53), .B(n_54), .Y(n_593) );
OA21x2_ASAP7_75t_L g594 ( .A1(n_504), .A2(n_56), .B(n_58), .Y(n_594) );
OA21x2_ASAP7_75t_L g595 ( .A1(n_504), .A2(n_61), .B(n_64), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_548), .B(n_66), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_555), .Y(n_597) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_547), .A2(n_68), .B(n_69), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_551), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_572), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_589), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_577), .B(n_76), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_589), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_562), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_562), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_563), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_568), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_579), .B(n_77), .Y(n_608) );
NOR2xp67_ASAP7_75t_SL g609 ( .A(n_565), .B(n_79), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_578), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_578), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_586), .B(n_80), .Y(n_612) );
INVx3_ASAP7_75t_L g613 ( .A(n_565), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g614 ( .A1(n_583), .A2(n_213), .B1(n_83), .B2(n_84), .Y(n_614) );
OA21x2_ASAP7_75t_L g615 ( .A1(n_545), .A2(n_82), .B(n_86), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_566), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_550), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_568), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_586), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_575), .A2(n_90), .B1(n_92), .B2(n_93), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_546), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_585), .B(n_211), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_569), .Y(n_624) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_536), .A2(n_94), .B(n_96), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_558), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_558), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_550), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_554), .Y(n_629) );
OAI21x1_ASAP7_75t_L g630 ( .A1(n_543), .A2(n_553), .B(n_590), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_549), .B(n_98), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_554), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_541), .Y(n_633) );
AO21x2_ASAP7_75t_L g634 ( .A1(n_542), .A2(n_99), .B(n_100), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_557), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_576), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_570), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_544), .Y(n_638) );
OAI21xp5_ASAP7_75t_L g639 ( .A1(n_573), .A2(n_108), .B(n_112), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_591), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_541), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_567), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_594), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_575), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_573), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_539), .A2(n_210), .B1(n_116), .B2(n_118), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_592), .Y(n_647) );
BUFx12f_ASAP7_75t_L g648 ( .A(n_557), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g649 ( .A(n_588), .Y(n_649) );
BUFx12f_ASAP7_75t_L g650 ( .A(n_560), .Y(n_650) );
AO21x1_ASAP7_75t_SL g651 ( .A1(n_539), .A2(n_114), .B(n_119), .Y(n_651) );
OA21x2_ASAP7_75t_L g652 ( .A1(n_559), .A2(n_121), .B(n_151), .Y(n_652) );
OAI21x1_ASAP7_75t_L g653 ( .A1(n_584), .A2(n_153), .B(n_156), .Y(n_653) );
BUFx2_ASAP7_75t_SL g654 ( .A(n_588), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_538), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_560), .Y(n_657) );
INVx2_ASAP7_75t_SL g658 ( .A(n_538), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_574), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_582), .Y(n_661) );
INVx3_ASAP7_75t_L g662 ( .A(n_564), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_556), .Y(n_663) );
BUFx2_ASAP7_75t_L g664 ( .A(n_582), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_540), .B(n_158), .Y(n_665) );
OAI21x1_ASAP7_75t_L g666 ( .A1(n_587), .A2(n_159), .B(n_160), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_580), .Y(n_667) );
OR2x6_ASAP7_75t_L g668 ( .A(n_593), .B(n_162), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_580), .Y(n_669) );
OAI21x1_ASAP7_75t_L g670 ( .A1(n_561), .A2(n_163), .B(n_165), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_564), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g672 ( .A(n_571), .B(n_167), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_540), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_571), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_595), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_644), .B(n_542), .Y(n_676) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_600), .Y(n_677) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_600), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_599), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_629), .A2(n_595), .B1(n_594), .B2(n_593), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_597), .Y(n_681) );
AND2x4_ASAP7_75t_L g682 ( .A(n_613), .B(n_175), .Y(n_682) );
BUFx3_ASAP7_75t_L g683 ( .A(n_613), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_624), .B(n_176), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_638), .B(n_181), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_602), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_642), .B(n_632), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_604), .B(n_184), .Y(n_688) );
INVx3_ASAP7_75t_L g689 ( .A(n_616), .Y(n_689) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_610), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_641), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_605), .B(n_185), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_637), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_619), .Y(n_694) );
INVx1_ASAP7_75t_SL g695 ( .A(n_617), .Y(n_695) );
AND2x2_ASAP7_75t_L g696 ( .A(n_654), .B(n_189), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_657), .B(n_190), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_616), .Y(n_698) );
AND2x4_ASAP7_75t_L g699 ( .A(n_607), .B(n_192), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_618), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_658), .Y(n_701) );
AND2x4_ASAP7_75t_L g702 ( .A(n_621), .B(n_193), .Y(n_702) );
AND2x4_ASAP7_75t_L g703 ( .A(n_622), .B(n_196), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_601), .B(n_537), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_649), .B(n_208), .Y(n_705) );
INVxp67_ASAP7_75t_L g706 ( .A(n_633), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_596), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_628), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_603), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_635), .B(n_201), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_596), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_649), .Y(n_712) );
NOR2x1p5_ASAP7_75t_L g713 ( .A(n_648), .B(n_204), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_606), .B(n_205), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_631), .B(n_207), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_631), .B(n_673), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_623), .B(n_612), .Y(n_717) );
NOR2x1_ASAP7_75t_R g718 ( .A(n_650), .B(n_665), .Y(n_718) );
INVxp67_ASAP7_75t_SL g719 ( .A(n_610), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_608), .Y(n_720) );
BUFx2_ASAP7_75t_L g721 ( .A(n_668), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_608), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_611), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_640), .Y(n_724) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_611), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_647), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_626), .B(n_627), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_645), .B(n_655), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_655), .B(n_661), .Y(n_729) );
BUFx6f_ASAP7_75t_L g730 ( .A(n_651), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_620), .B(n_614), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_620), .B(n_614), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_639), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_639), .B(n_664), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_668), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_659), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_660), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_662), .Y(n_738) );
NAND2x1_ASAP7_75t_L g739 ( .A(n_609), .B(n_668), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_653), .Y(n_740) );
INVxp67_ASAP7_75t_L g741 ( .A(n_667), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_666), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_646), .B(n_669), .Y(n_743) );
BUFx3_ASAP7_75t_L g744 ( .A(n_625), .Y(n_744) );
AND2x2_ASAP7_75t_L g745 ( .A(n_646), .B(n_598), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_671), .B(n_634), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_670), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_656), .B(n_672), .Y(n_748) );
INVxp67_ASAP7_75t_L g749 ( .A(n_662), .Y(n_749) );
AND2x4_ASAP7_75t_SL g750 ( .A(n_636), .B(n_663), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_672), .B(n_643), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_652), .B(n_643), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_674), .Y(n_753) );
AND2x4_ASAP7_75t_SL g754 ( .A(n_675), .B(n_615), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_675), .B(n_615), .Y(n_755) );
NOR2xp67_ASAP7_75t_L g756 ( .A(n_630), .B(n_635), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_687), .B(n_709), .Y(n_757) );
NAND2x1p5_ASAP7_75t_L g758 ( .A(n_739), .B(n_735), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_679), .Y(n_759) );
AND2x4_ASAP7_75t_L g760 ( .A(n_735), .B(n_756), .Y(n_760) );
BUFx3_ASAP7_75t_L g761 ( .A(n_683), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_681), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_718), .B(n_693), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_712), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_700), .B(n_717), .Y(n_765) );
BUFx3_ASAP7_75t_L g766 ( .A(n_683), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_694), .Y(n_767) );
BUFx3_ASAP7_75t_L g768 ( .A(n_689), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_691), .B(n_677), .Y(n_769) );
INVx2_ASAP7_75t_L g770 ( .A(n_736), .Y(n_770) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_677), .Y(n_771) );
AND2x4_ASAP7_75t_L g772 ( .A(n_721), .B(n_726), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_678), .B(n_716), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_706), .B(n_695), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_676), .B(n_724), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_698), .B(n_706), .Y(n_776) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_690), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_689), .B(n_686), .Y(n_778) );
INVx3_ASAP7_75t_L g779 ( .A(n_750), .Y(n_779) );
INVx1_ASAP7_75t_SL g780 ( .A(n_705), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_737), .Y(n_781) );
HB1xp67_ASAP7_75t_L g782 ( .A(n_690), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_708), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_720), .B(n_722), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_707), .B(n_711), .Y(n_785) );
INVx3_ASAP7_75t_L g786 ( .A(n_750), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_741), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_727), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_725), .Y(n_789) );
NAND2x1p5_ASAP7_75t_L g790 ( .A(n_682), .B(n_730), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_731), .B(n_732), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_723), .Y(n_792) );
INVx3_ASAP7_75t_L g793 ( .A(n_730), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_728), .Y(n_794) );
AND2x2_ASAP7_75t_L g795 ( .A(n_688), .B(n_696), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_753), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_729), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_749), .B(n_738), .Y(n_798) );
AND2x2_ASAP7_75t_L g799 ( .A(n_697), .B(n_684), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_733), .B(n_743), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_729), .Y(n_801) );
AND2x4_ASAP7_75t_L g802 ( .A(n_749), .B(n_738), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_713), .A2(n_745), .B1(n_734), .B2(n_704), .Y(n_803) );
HB1xp67_ASAP7_75t_L g804 ( .A(n_701), .Y(n_804) );
AND2x4_ASAP7_75t_L g805 ( .A(n_719), .B(n_701), .Y(n_805) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_685), .A2(n_714), .B1(n_710), .B2(n_680), .C(n_704), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_752), .Y(n_807) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_751), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_702), .Y(n_809) );
AND2x2_ASAP7_75t_L g810 ( .A(n_692), .B(n_699), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_755), .Y(n_811) );
INVx1_ASAP7_75t_SL g812 ( .A(n_703), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_699), .B(n_703), .Y(n_813) );
AND2x2_ASAP7_75t_L g814 ( .A(n_746), .B(n_715), .Y(n_814) );
INVx2_ASAP7_75t_L g815 ( .A(n_755), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_759), .Y(n_816) );
AND2x2_ASAP7_75t_L g817 ( .A(n_807), .B(n_748), .Y(n_817) );
AND2x2_ASAP7_75t_L g818 ( .A(n_773), .B(n_742), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_767), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_791), .B(n_740), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_757), .Y(n_821) );
INVx3_ASAP7_75t_L g822 ( .A(n_758), .Y(n_822) );
INVx2_ASAP7_75t_L g823 ( .A(n_770), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_761), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_787), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_781), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_775), .B(n_754), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_775), .B(n_754), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_788), .B(n_680), .Y(n_829) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_804), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_775), .B(n_744), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_814), .B(n_747), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_771), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_771), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_797), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_800), .B(n_774), .Y(n_836) );
INVx1_ASAP7_75t_SL g837 ( .A(n_764), .Y(n_837) );
OR2x2_ASAP7_75t_L g838 ( .A(n_789), .B(n_777), .Y(n_838) );
INVx2_ASAP7_75t_L g839 ( .A(n_811), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_765), .B(n_769), .Y(n_840) );
AND2x2_ASAP7_75t_L g841 ( .A(n_794), .B(n_801), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_784), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_808), .B(n_796), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_811), .B(n_815), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_815), .B(n_805), .Y(n_845) );
AND2x2_ASAP7_75t_L g846 ( .A(n_805), .B(n_792), .Y(n_846) );
INVx2_ASAP7_75t_SL g847 ( .A(n_761), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_805), .B(n_792), .Y(n_848) );
OR2x2_ASAP7_75t_L g849 ( .A(n_836), .B(n_782), .Y(n_849) );
INVx1_ASAP7_75t_L g850 ( .A(n_816), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_842), .B(n_785), .Y(n_851) );
INVx3_ASAP7_75t_SL g852 ( .A(n_847), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_837), .B(n_763), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_SL g854 ( .A1(n_847), .A2(n_763), .B(n_780), .C(n_812), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_819), .Y(n_855) );
INVx3_ASAP7_75t_L g856 ( .A(n_824), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_841), .B(n_762), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_832), .B(n_772), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_826), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_838), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_838), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_843), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_832), .B(n_776), .Y(n_863) );
AND2x4_ASAP7_75t_L g864 ( .A(n_831), .B(n_760), .Y(n_864) );
AOI22xp33_ASAP7_75t_SL g865 ( .A1(n_822), .A2(n_813), .B1(n_758), .B2(n_810), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_830), .Y(n_866) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_833), .B(n_762), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_836), .B(n_777), .Y(n_868) );
INVx2_ASAP7_75t_SL g869 ( .A(n_852), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g870 ( .A(n_860), .B(n_834), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_849), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_868), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_857), .Y(n_873) );
AOI332xp33_ASAP7_75t_L g874 ( .A1(n_861), .A2(n_821), .A3(n_825), .B1(n_835), .B2(n_820), .B3(n_803), .C1(n_840), .C2(n_818), .Y(n_874) );
NOR3xp33_ASAP7_75t_L g875 ( .A(n_853), .B(n_806), .C(n_829), .Y(n_875) );
AND2x2_ASAP7_75t_L g876 ( .A(n_858), .B(n_827), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_867), .B(n_844), .Y(n_877) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_867), .B(n_844), .Y(n_878) );
NAND2x1_ASAP7_75t_L g879 ( .A(n_856), .B(n_760), .Y(n_879) );
INVx2_ASAP7_75t_L g880 ( .A(n_863), .Y(n_880) );
NOR4xp25_ASAP7_75t_L g881 ( .A(n_869), .B(n_854), .C(n_866), .D(n_851), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_876), .B(n_864), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_873), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g884 ( .A1(n_875), .A2(n_865), .B1(n_854), .B2(n_818), .Y(n_884) );
AOI22xp5_ASAP7_75t_L g885 ( .A1(n_871), .A2(n_831), .B1(n_845), .B2(n_862), .Y(n_885) );
AOI211x1_ASAP7_75t_L g886 ( .A1(n_872), .A2(n_859), .B(n_855), .C(n_850), .Y(n_886) );
AOI21xp5_ASAP7_75t_L g887 ( .A1(n_881), .A2(n_879), .B(n_870), .Y(n_887) );
AOI211xp5_ASAP7_75t_SL g888 ( .A1(n_884), .A2(n_793), .B(n_760), .C(n_809), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g889 ( .A1(n_886), .A2(n_878), .B1(n_877), .B2(n_880), .C(n_874), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_883), .Y(n_890) );
NOR2x1_ASAP7_75t_L g891 ( .A(n_887), .B(n_766), .Y(n_891) );
NAND5xp2_ASAP7_75t_L g892 ( .A(n_888), .B(n_790), .C(n_885), .D(n_795), .E(n_799), .Y(n_892) );
NAND4xp75_ASAP7_75t_L g893 ( .A(n_891), .B(n_889), .C(n_890), .D(n_882), .Y(n_893) );
NAND4xp25_ASAP7_75t_L g894 ( .A(n_892), .B(n_793), .C(n_768), .D(n_786), .Y(n_894) );
OAI211xp5_ASAP7_75t_L g895 ( .A1(n_894), .A2(n_793), .B(n_768), .C(n_786), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_893), .B(n_828), .Y(n_896) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_896), .A2(n_778), .B1(n_828), .B2(n_827), .Y(n_897) );
BUFx2_ASAP7_75t_L g898 ( .A(n_895), .Y(n_898) );
OA22x2_ASAP7_75t_L g899 ( .A1(n_898), .A2(n_786), .B1(n_779), .B2(n_802), .Y(n_899) );
AND2x4_ASAP7_75t_L g900 ( .A(n_897), .B(n_848), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_899), .Y(n_901) );
OAI22x1_ASAP7_75t_L g902 ( .A1(n_901), .A2(n_900), .B1(n_779), .B2(n_798), .Y(n_902) );
AOI21xp5_ASAP7_75t_L g903 ( .A1(n_902), .A2(n_779), .B(n_783), .Y(n_903) );
OR2x6_ASAP7_75t_L g904 ( .A(n_903), .B(n_848), .Y(n_904) );
AOI22xp5_ASAP7_75t_SL g905 ( .A1(n_904), .A2(n_846), .B1(n_817), .B2(n_782), .Y(n_905) );
BUFx3_ASAP7_75t_L g906 ( .A(n_905), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g907 ( .A1(n_906), .A2(n_839), .B(n_823), .Y(n_907) );
endmodule