module fake_netlist_6_853_n_2400 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2400);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2400;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2382;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_1371;
wire n_1285;
wire n_383;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_322;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_2368;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_1141;
wire n_562;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_2374;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2373;
wire n_1472;
wire n_2050;
wire n_2120;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g230 ( 
.A(n_169),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_105),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_27),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_110),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_75),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_53),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_202),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_30),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_32),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_164),
.Y(n_242)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_55),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_97),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_97),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_119),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_217),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_186),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_209),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_41),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_178),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_43),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_175),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_6),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_65),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_112),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_204),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_224),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_35),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_64),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_74),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_142),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_54),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_69),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_5),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_143),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_8),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_191),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_64),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_2),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_199),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_170),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_36),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_188),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_155),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_90),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_19),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_121),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_30),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_115),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_141),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_105),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_29),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_212),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_208),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_226),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_162),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_45),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_203),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_88),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_71),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_223),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_221),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_150),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_136),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_126),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_190),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_51),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_4),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_61),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_116),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_55),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_44),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_177),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_108),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_139),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_78),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_70),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_147),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_3),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_104),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_92),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_195),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_69),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_7),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_102),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_78),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_137),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_99),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_86),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_98),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_182),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_15),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_1),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_218),
.Y(n_334)
);

BUFx8_ASAP7_75t_SL g335 ( 
.A(n_47),
.Y(n_335)
);

BUFx2_ASAP7_75t_SL g336 ( 
.A(n_98),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_8),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_154),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_125),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_146),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_216),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_213),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_181),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_54),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_153),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_32),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_24),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_163),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_201),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_72),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_40),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_7),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_90),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_91),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_27),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_120),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_46),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_87),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_193),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_159),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_228),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_86),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_144),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_2),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_28),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_165),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_149),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_160),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_48),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_134),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_41),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_176),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_24),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_72),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_198),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_106),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_87),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_103),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_171),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_63),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_0),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_67),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_84),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_50),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_100),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_11),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_104),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_63),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_82),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_219),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_52),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_167),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_4),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_14),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_100),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_205),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_80),
.Y(n_397)
);

BUFx3_ASAP7_75t_L g398 ( 
.A(n_23),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_174),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_75),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_225),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_58),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_94),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_151),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_38),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_93),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_118),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_94),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_1),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_183),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_34),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_88),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_9),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_92),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_5),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_66),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_43),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_227),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_21),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_185),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_180),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_81),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_77),
.Y(n_423)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_19),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_67),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_117),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_168),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_12),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_103),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_36),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g431 ( 
.A(n_140),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_12),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_47),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_135),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_122),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_66),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_197),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_15),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_194),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_189),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_80),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_152),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_114),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_109),
.Y(n_444)
);

BUFx2_ASAP7_75t_SL g445 ( 
.A(n_17),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_44),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_79),
.Y(n_447)
);

INVx2_ASAP7_75t_SL g448 ( 
.A(n_35),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_84),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_123),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_38),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_131),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_335),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_243),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_243),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_238),
.Y(n_456)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_409),
.B(n_6),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_243),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_264),
.B(n_9),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_240),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_248),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_244),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_243),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_249),
.Y(n_464)
);

BUFx6f_ASAP7_75t_SL g465 ( 
.A(n_290),
.Y(n_465)
);

NOR2xp67_ASAP7_75t_L g466 ( 
.A(n_409),
.B(n_10),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_243),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_255),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_283),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_258),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_243),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g472 ( 
.A(n_264),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_243),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_10),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_243),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_244),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_259),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_242),
.B(n_11),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g480 ( 
.A(n_246),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_243),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_292),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_424),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_260),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_424),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_424),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_424),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_424),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_339),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_334),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_424),
.B(n_13),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_339),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_424),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_399),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_231),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_424),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_271),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_246),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_250),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_262),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_273),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_381),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_250),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_235),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_380),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_242),
.B(n_13),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_278),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_280),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g511 ( 
.A(n_431),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_381),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_285),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_276),
.B(n_14),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_286),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_289),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_448),
.B(n_16),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_291),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_R g520 ( 
.A(n_295),
.B(n_107),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_381),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_381),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_301),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_311),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_313),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_381),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_237),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_381),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_388),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_320),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_265),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_388),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_388),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_388),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_338),
.Y(n_535)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_262),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_376),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_343),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_345),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_356),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_388),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_359),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_388),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_257),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_257),
.Y(n_545)
);

BUFx2_ASAP7_75t_SL g546 ( 
.A(n_276),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_368),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_306),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_277),
.B(n_16),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_239),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_277),
.B(n_18),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_360),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_342),
.B(n_18),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_306),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_364),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_363),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_407),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_364),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_371),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_372),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_375),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_371),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_390),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_392),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_374),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_245),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_396),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_374),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_232),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_232),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_342),
.B(n_20),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_427),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_241),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_288),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_247),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_504),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_504),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_456),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_460),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_476),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_480),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_531),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_512),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_512),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_522),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_461),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_546),
.B(n_479),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

CKINVDCx8_ASAP7_75t_R g589 ( 
.A(n_480),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_574),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_531),
.Y(n_591)
);

OA21x2_ASAP7_75t_L g592 ( 
.A1(n_492),
.A2(n_256),
.B(n_241),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_522),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_521),
.B(n_401),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_478),
.B(n_394),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_464),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_531),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_537),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_531),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_526),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_401),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_468),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_537),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_574),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_490),
.B(n_434),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_526),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_470),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_528),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_493),
.B(n_452),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_454),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_477),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_528),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_529),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_459),
.B(n_278),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_484),
.B(n_437),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_529),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_508),
.B(n_251),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_499),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_454),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_469),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_537),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_532),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_482),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_455),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_491),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_532),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_533),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

OA21x2_ASAP7_75t_L g631 ( 
.A1(n_492),
.A2(n_263),
.B(n_256),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_458),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_458),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_533),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_463),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_503),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_495),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_516),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_500),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_463),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_519),
.Y(n_642)
);

CKINVDCx16_ASAP7_75t_R g643 ( 
.A(n_465),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_534),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_467),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_541),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_467),
.Y(n_647)
);

INVxp67_ASAP7_75t_L g648 ( 
.A(n_496),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_541),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_511),
.B(n_288),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_471),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_543),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_471),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_457),
.B(n_466),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_543),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_569),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_473),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_525),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_501),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_517),
.B(n_319),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_530),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_475),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_505),
.Y(n_666)
);

OA21x2_ASAP7_75t_L g667 ( 
.A1(n_475),
.A2(n_267),
.B(n_263),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_466),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_474),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_481),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_538),
.Y(n_671)
);

CKINVDCx20_ASAP7_75t_R g672 ( 
.A(n_581),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_619),
.B(n_539),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_587),
.B(n_540),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_643),
.B(n_542),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_667),
.Y(n_676)
);

INVx5_ASAP7_75t_L g677 ( 
.A(n_599),
.Y(n_677)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_626),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_667),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_587),
.B(n_556),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_628),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_663),
.Y(n_682)
);

INVx8_ASAP7_75t_L g683 ( 
.A(n_594),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_667),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_599),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_617),
.Y(n_686)
);

OAI22xp33_ASAP7_75t_L g687 ( 
.A1(n_615),
.A2(n_472),
.B1(n_509),
.B2(n_486),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_667),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_643),
.B(n_561),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_663),
.B(n_517),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_667),
.Y(n_691)
);

AND2x2_ASAP7_75t_SL g692 ( 
.A(n_615),
.B(n_514),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_592),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_580),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_619),
.A2(n_668),
.B1(n_669),
.B2(n_616),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_617),
.B(n_564),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_590),
.B(n_605),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_667),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_630),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_663),
.B(n_517),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_594),
.B(n_567),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_592),
.Y(n_702)
);

INVxp67_ASAP7_75t_SL g703 ( 
.A(n_630),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_628),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_578),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_SL g706 ( 
.A(n_589),
.B(n_453),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_590),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_630),
.Y(n_708)
);

INVxp67_ASAP7_75t_SL g709 ( 
.A(n_630),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_630),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_650),
.B(n_502),
.Y(n_711)
);

AO21x2_ASAP7_75t_L g712 ( 
.A1(n_655),
.A2(n_233),
.B(n_230),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_633),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_579),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_599),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_648),
.B(n_572),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_628),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_606),
.B(n_510),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_646),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_605),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_599),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_580),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_648),
.B(n_509),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_599),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_671),
.B(n_513),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_650),
.B(n_536),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_650),
.B(n_230),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_592),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_599),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_594),
.B(n_547),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_594),
.B(n_557),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_633),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_606),
.B(n_515),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_616),
.B(n_507),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_646),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_599),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_599),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_668),
.B(n_507),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_626),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_600),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_633),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_600),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_669),
.B(n_544),
.Y(n_743)
);

INVx1_ASAP7_75t_SL g744 ( 
.A(n_639),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_595),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_646),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_589),
.B(n_523),
.Y(n_747)
);

BUFx3_ASAP7_75t_L g748 ( 
.A(n_592),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_655),
.B(n_336),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_L g750 ( 
.A1(n_581),
.A2(n_474),
.B1(n_518),
.B2(n_462),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_594),
.B(n_233),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_586),
.B(n_524),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_633),
.Y(n_753)
);

INVxp33_ASAP7_75t_SL g754 ( 
.A(n_596),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_611),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_595),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_611),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_610),
.B(n_535),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_481),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_611),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_603),
.B(n_552),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_610),
.B(n_560),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_602),
.B(n_483),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_633),
.B(n_265),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_608),
.B(n_563),
.Y(n_765)
);

OAI21xp33_ASAP7_75t_L g766 ( 
.A1(n_657),
.A2(n_551),
.B(n_549),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_635),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_626),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_611),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_621),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_657),
.B(n_658),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_658),
.B(n_234),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_612),
.A2(n_465),
.B1(n_527),
.B2(n_506),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_600),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_620),
.B(n_550),
.Y(n_775)
);

AND2x6_ASAP7_75t_L g776 ( 
.A(n_635),
.B(n_265),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_600),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_635),
.B(n_483),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_592),
.A2(n_571),
.B1(n_553),
.B2(n_518),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_592),
.B(n_544),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_635),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_631),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_631),
.B(n_566),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_636),
.B(n_575),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_639),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_638),
.B(n_465),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_662),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_635),
.Y(n_788)
);

NAND3x1_ASAP7_75t_L g789 ( 
.A(n_660),
.B(n_294),
.C(n_267),
.Y(n_789)
);

BUFx4f_ASAP7_75t_L g790 ( 
.A(n_631),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_645),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_234),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_645),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_626),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_600),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_589),
.A2(n_406),
.B1(n_252),
.B2(n_261),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_631),
.B(n_545),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_645),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_642),
.B(n_465),
.Y(n_799)
);

NOR2x1p5_ASAP7_75t_L g800 ( 
.A(n_661),
.B(n_319),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_645),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_664),
.B(n_645),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_L g803 ( 
.A(n_626),
.B(n_265),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_600),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_647),
.B(n_435),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_576),
.B(n_236),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_621),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_647),
.B(n_485),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_631),
.A2(n_398),
.B1(n_325),
.B2(n_296),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_647),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_621),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_647),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_631),
.A2(n_440),
.B1(n_442),
.B2(n_439),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_647),
.B(n_254),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_651),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_651),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_651),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_651),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_621),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_626),
.Y(n_820)
);

BUFx8_ASAP7_75t_SL g821 ( 
.A(n_622),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_651),
.B(n_268),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_632),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_632),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_576),
.B(n_269),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_626),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_577),
.B(n_270),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_632),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_577),
.B(n_545),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_632),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_670),
.B(n_485),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_654),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_597),
.B(n_236),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_805),
.B(n_626),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_673),
.B(n_640),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_690),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_759),
.B(n_640),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_692),
.A2(n_444),
.B1(n_279),
.B2(n_300),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_771),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_L g840 ( 
.A(n_683),
.B(n_265),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_692),
.A2(n_340),
.B1(n_366),
.B2(n_312),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_676),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_763),
.B(n_640),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_SL g844 ( 
.A1(n_672),
.A2(n_666),
.B1(n_662),
.B2(n_625),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_683),
.A2(n_597),
.B(n_670),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_814),
.B(n_640),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_693),
.A2(n_296),
.B1(n_310),
.B2(n_294),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_676),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_679),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_679),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_822),
.B(n_640),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_802),
.B(n_640),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_640),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_693),
.A2(n_315),
.B1(n_318),
.B2(n_310),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_690),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_680),
.B(n_640),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_771),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_682),
.B(n_730),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_790),
.A2(n_318),
.B(n_323),
.C(n_315),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_684),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_684),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_688),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_790),
.B(n_653),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_682),
.B(n_653),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_790),
.B(n_653),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_697),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_771),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_731),
.B(n_653),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_683),
.B(n_653),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_702),
.A2(n_328),
.B1(n_337),
.B2(n_323),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_818),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_683),
.B(n_751),
.Y(n_872)
);

NAND2x1_ASAP7_75t_L g873 ( 
.A(n_688),
.B(n_597),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_695),
.B(n_272),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_818),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_751),
.B(n_653),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_751),
.B(n_653),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_691),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_703),
.B(n_653),
.Y(n_879)
);

AO22x1_ASAP7_75t_L g880 ( 
.A1(n_756),
.A2(n_337),
.B1(n_344),
.B2(n_328),
.Y(n_880)
);

AND2x6_ASAP7_75t_SL g881 ( 
.A(n_775),
.B(n_344),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_709),
.B(n_654),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_691),
.B(n_654),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_718),
.A2(n_279),
.B1(n_300),
.B2(n_253),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_733),
.A2(n_302),
.B1(n_303),
.B2(n_253),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_783),
.B(n_265),
.Y(n_886)
);

O2A1O1Ixp5_ASAP7_75t_L g887 ( 
.A1(n_698),
.A2(n_659),
.B(n_665),
.C(n_654),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_698),
.B(n_659),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_701),
.B(n_659),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_702),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_783),
.B(n_274),
.Y(n_891)
);

NAND3xp33_ASAP7_75t_SL g892 ( 
.A(n_694),
.B(n_422),
.C(n_405),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_758),
.A2(n_303),
.B1(n_308),
.B2(n_302),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_707),
.B(n_278),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_734),
.B(n_336),
.Y(n_895)
);

INVx8_ASAP7_75t_L g896 ( 
.A(n_749),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_L g897 ( 
.A1(n_728),
.A2(n_352),
.B1(n_387),
.B2(n_347),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_681),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_707),
.B(n_278),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_779),
.B(n_700),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_700),
.B(n_659),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_712),
.B(n_665),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_681),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_704),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_829),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_711),
.B(n_281),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_762),
.B(n_275),
.Y(n_907)
);

NAND3xp33_ASAP7_75t_L g908 ( 
.A(n_711),
.B(n_284),
.C(n_282),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_704),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_829),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_782),
.A2(n_670),
.B(n_665),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_712),
.B(n_665),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_L g913 ( 
.A(n_687),
.B(n_293),
.C(n_287),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_749),
.B(n_297),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_780),
.Y(n_915)
);

A2O1A1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_780),
.A2(n_352),
.B(n_387),
.C(n_347),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_797),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_L g918 ( 
.A(n_686),
.B(n_734),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_726),
.B(n_281),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_717),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_SL g921 ( 
.A(n_722),
.B(n_666),
.C(n_625),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_749),
.A2(n_316),
.B1(n_327),
.B2(n_308),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_782),
.A2(n_670),
.B(n_400),
.C(n_403),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_749),
.A2(n_316),
.B1(n_331),
.B2(n_327),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_712),
.B(n_583),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_797),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_728),
.B(n_266),
.Y(n_927)
);

INVxp67_ASAP7_75t_L g928 ( 
.A(n_738),
.Y(n_928)
);

AND2x6_ASAP7_75t_L g929 ( 
.A(n_748),
.B(n_331),
.Y(n_929)
);

INVx2_ASAP7_75t_SL g930 ( 
.A(n_697),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_717),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_772),
.B(n_792),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_778),
.A2(n_597),
.B(n_600),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_748),
.Y(n_934)
);

INVxp67_ASAP7_75t_L g935 ( 
.A(n_738),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_699),
.B(n_583),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_808),
.A2(n_597),
.B(n_600),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_719),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_699),
.B(n_584),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_715),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_772),
.B(n_341),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_715),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_708),
.B(n_584),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_708),
.B(n_585),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_813),
.B(n_266),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_715),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_710),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_710),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_713),
.B(n_585),
.Y(n_949)
);

INVx3_ASAP7_75t_L g950 ( 
.A(n_772),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_715),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_713),
.Y(n_952)
);

OAI221xp5_ASAP7_75t_L g953 ( 
.A1(n_766),
.A2(n_400),
.B1(n_425),
.B2(n_429),
.C(n_414),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_727),
.A2(n_348),
.B1(n_349),
.B2(n_341),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_732),
.B(n_593),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_732),
.B(n_593),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_L g957 ( 
.A1(n_809),
.A2(n_403),
.B1(n_411),
.B2(n_393),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_741),
.B(n_601),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_715),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_741),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_719),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_753),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_753),
.B(n_767),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_726),
.B(n_304),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_716),
.B(n_305),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_727),
.B(n_307),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_735),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_767),
.B(n_601),
.Y(n_968)
);

OAI22xp33_ASAP7_75t_L g969 ( 
.A1(n_745),
.A2(n_349),
.B1(n_361),
.B2(n_348),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_781),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_781),
.B(n_607),
.Y(n_971)
);

OAI22xp33_ASAP7_75t_L g972 ( 
.A1(n_745),
.A2(n_367),
.B1(n_370),
.B2(n_361),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_788),
.B(n_607),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_727),
.B(n_309),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_720),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_686),
.B(n_266),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_833),
.B(n_266),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_735),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_750),
.B(n_314),
.Y(n_979)
);

NOR2x1p5_ASAP7_75t_L g980 ( 
.A(n_743),
.B(n_325),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_743),
.A2(n_800),
.B1(n_723),
.B2(n_696),
.Y(n_981)
);

AOI22xp33_ASAP7_75t_L g982 ( 
.A1(n_792),
.A2(n_411),
.B1(n_412),
.B2(n_393),
.Y(n_982)
);

BUFx8_ASAP7_75t_L g983 ( 
.A(n_720),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_773),
.A2(n_420),
.B1(n_312),
.B2(n_340),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_705),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_788),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_791),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_791),
.B(n_609),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_821),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_793),
.B(n_609),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_793),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_798),
.B(n_613),
.Y(n_992)
);

NOR2x1p5_ASAP7_75t_L g993 ( 
.A(n_706),
.B(n_398),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_798),
.B(n_613),
.Y(n_994)
);

AND2x4_ASAP7_75t_L g995 ( 
.A(n_792),
.B(n_806),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_796),
.B(n_317),
.Y(n_996)
);

NAND2x1_ASAP7_75t_L g997 ( 
.A(n_685),
.B(n_614),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_801),
.B(n_614),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_784),
.B(n_321),
.Y(n_999)
);

OR2x6_ASAP7_75t_L g1000 ( 
.A(n_725),
.B(n_445),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_801),
.B(n_618),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_787),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_721),
.Y(n_1003)
);

AOI221xp5_ASAP7_75t_L g1004 ( 
.A1(n_825),
.A2(n_414),
.B1(n_429),
.B2(n_425),
.C(n_412),
.Y(n_1004)
);

NAND2x1p5_ASAP7_75t_L g1005 ( 
.A(n_806),
.B(n_367),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_L g1006 ( 
.A(n_785),
.B(n_761),
.C(n_752),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_827),
.A2(n_450),
.B1(n_443),
.B2(n_426),
.Y(n_1007)
);

INVx2_ASAP7_75t_SL g1008 ( 
.A(n_806),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_810),
.B(n_618),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_947),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_948),
.Y(n_1011)
);

INVx2_ASAP7_75t_SL g1012 ( 
.A(n_836),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_907),
.B(n_981),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_SL g1014 ( 
.A(n_907),
.B(n_744),
.C(n_627),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_975),
.Y(n_1015)
);

AND2x6_ASAP7_75t_SL g1016 ( 
.A(n_996),
.B(n_765),
.Y(n_1016)
);

BUFx2_ASAP7_75t_L g1017 ( 
.A(n_983),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_898),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_844),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_952),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_900),
.A2(n_833),
.B1(n_786),
.B2(n_799),
.Y(n_1021)
);

BUFx8_ASAP7_75t_L g1022 ( 
.A(n_1002),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_960),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_858),
.B(n_810),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_905),
.B(n_705),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_898),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_983),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_926),
.B(n_812),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_890),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_903),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_836),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_928),
.B(n_754),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_903),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_989),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_921),
.B(n_622),
.Y(n_1035)
);

INVx8_ASAP7_75t_L g1036 ( 
.A(n_896),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_894),
.Y(n_1037)
);

INVx6_ASAP7_75t_L g1038 ( 
.A(n_932),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_962),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_904),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_899),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_866),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_855),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_930),
.B(n_675),
.Y(n_1044)
);

BUFx2_ASAP7_75t_L g1045 ( 
.A(n_983),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_985),
.B(n_627),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_855),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_890),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_932),
.B(n_995),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_890),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_890),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_904),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_985),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_926),
.B(n_812),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_935),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_932),
.B(n_995),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_915),
.B(n_815),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_995),
.B(n_747),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_996),
.B(n_754),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_895),
.B(n_906),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_R g1061 ( 
.A(n_892),
.B(n_637),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_839),
.B(n_689),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_934),
.Y(n_1063)
);

NOR2xp67_ASAP7_75t_L g1064 ( 
.A(n_908),
.B(n_965),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_1000),
.Y(n_1065)
);

OR2x2_ASAP7_75t_L g1066 ( 
.A(n_919),
.B(n_445),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_970),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_917),
.B(n_815),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_891),
.B(n_816),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_909),
.Y(n_1070)
);

NAND2xp33_ASAP7_75t_SL g1071 ( 
.A(n_934),
.B(n_672),
.Y(n_1071)
);

CKINVDCx20_ASAP7_75t_R g1072 ( 
.A(n_896),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_857),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_986),
.Y(n_1074)
);

BUFx3_ASAP7_75t_L g1075 ( 
.A(n_867),
.Y(n_1075)
);

INVxp33_ASAP7_75t_SL g1076 ( 
.A(n_1006),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_891),
.B(n_816),
.Y(n_1077)
);

OAI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_838),
.A2(n_833),
.B1(n_370),
.B2(n_410),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_945),
.A2(n_817),
.B1(n_420),
.B2(n_366),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_934),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_910),
.B(n_705),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_964),
.B(n_714),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_987),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_934),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_896),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_991),
.Y(n_1086)
);

HB1xp67_ASAP7_75t_L g1087 ( 
.A(n_980),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_835),
.B(n_817),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_993),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_950),
.B(n_637),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_1008),
.B(n_379),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_929),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_SL g1093 ( 
.A(n_999),
.B(n_714),
.Y(n_1093)
);

INVx5_ASAP7_75t_L g1094 ( 
.A(n_929),
.Y(n_1094)
);

INVx5_ASAP7_75t_L g1095 ( 
.A(n_929),
.Y(n_1095)
);

INVx3_ASAP7_75t_L g1096 ( 
.A(n_871),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_964),
.B(n_714),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_942),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1000),
.B(n_874),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_909),
.Y(n_1100)
);

AOI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_950),
.A2(n_824),
.B1(n_828),
.B2(n_823),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_942),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_889),
.B(n_823),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_842),
.B(n_824),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_1005),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_963),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_920),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_942),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_842),
.B(n_828),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_871),
.Y(n_1110)
);

AO22x1_ASAP7_75t_L g1111 ( 
.A1(n_929),
.A2(n_410),
.B1(n_418),
.B2(n_379),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_941),
.B(n_418),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_1000),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_966),
.B(n_755),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_966),
.B(n_755),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_875),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_931),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_941),
.B(n_421),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_931),
.Y(n_1119)
);

NOR2x1_ASAP7_75t_SL g1120 ( 
.A(n_942),
.B(n_678),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_848),
.B(n_832),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_938),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_938),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_929),
.A2(n_832),
.B1(n_739),
.B2(n_768),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_961),
.Y(n_1125)
);

NAND2xp33_ASAP7_75t_SL g1126 ( 
.A(n_847),
.B(n_787),
.Y(n_1126)
);

NOR3xp33_ASAP7_75t_SL g1127 ( 
.A(n_874),
.B(n_324),
.C(n_322),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_961),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_SL g1129 ( 
.A(n_979),
.B(n_329),
.C(n_326),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_875),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1005),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_941),
.Y(n_1132)
);

BUFx10_ASAP7_75t_L g1133 ( 
.A(n_965),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_945),
.A2(n_426),
.B1(n_443),
.B2(n_421),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_967),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_967),
.Y(n_1136)
);

OR2x2_ASAP7_75t_SL g1137 ( 
.A(n_881),
.B(n_438),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_848),
.B(n_849),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_849),
.B(n_757),
.Y(n_1139)
);

BUFx3_ASAP7_75t_L g1140 ( 
.A(n_901),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_850),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_850),
.B(n_757),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_978),
.Y(n_1143)
);

BUFx3_ASAP7_75t_L g1144 ( 
.A(n_860),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_914),
.B(n_721),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_978),
.Y(n_1146)
);

NAND2xp33_ASAP7_75t_SL g1147 ( 
.A(n_847),
.B(n_450),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_860),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_R g1149 ( 
.A(n_999),
.B(n_685),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_914),
.B(n_979),
.Y(n_1150)
);

NOR3xp33_ASAP7_75t_SL g1151 ( 
.A(n_969),
.B(n_332),
.C(n_330),
.Y(n_1151)
);

BUFx4f_ASAP7_75t_L g1152 ( 
.A(n_946),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_861),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_861),
.B(n_760),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_884),
.B(n_721),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_862),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_885),
.B(n_721),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_862),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_SL g1159 ( 
.A(n_913),
.B(n_520),
.C(n_346),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_SL g1160 ( 
.A(n_972),
.B(n_350),
.C(n_333),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_872),
.B(n_918),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_878),
.B(n_760),
.Y(n_1162)
);

OR2x6_ASAP7_75t_L g1163 ( 
.A(n_880),
.B(n_789),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_916),
.Y(n_1164)
);

OR2x2_ASAP7_75t_SL g1165 ( 
.A(n_922),
.B(n_438),
.Y(n_1165)
);

AOI221xp5_ASAP7_75t_L g1166 ( 
.A1(n_1004),
.A2(n_441),
.B1(n_449),
.B2(n_432),
.C(n_428),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_974),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_878),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_946),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1009),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_887),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_976),
.B(n_974),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_946),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_976),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_883),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_946),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_893),
.B(n_721),
.Y(n_1177)
);

INVx4_ASAP7_75t_L g1178 ( 
.A(n_951),
.Y(n_1178)
);

AOI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_886),
.A2(n_678),
.B1(n_739),
.B2(n_826),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_936),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_951),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_939),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_957),
.B(n_769),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_916),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_886),
.B(n_854),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_957),
.B(n_769),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_951),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_854),
.B(n_770),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_951),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_943),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_841),
.Y(n_1191)
);

NOR3xp33_ASAP7_75t_SL g1192 ( 
.A(n_953),
.B(n_353),
.C(n_351),
.Y(n_1192)
);

AND3x2_ASAP7_75t_SL g1193 ( 
.A(n_859),
.B(n_789),
.C(n_382),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1003),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_924),
.B(n_678),
.Y(n_1195)
);

NOR3xp33_ASAP7_75t_SL g1196 ( 
.A(n_984),
.B(n_355),
.C(n_354),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_864),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_944),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_870),
.B(n_770),
.Y(n_1199)
);

HB1xp67_ASAP7_75t_L g1200 ( 
.A(n_954),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_870),
.B(n_807),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_897),
.B(n_807),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_897),
.B(n_811),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_949),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1106),
.B(n_868),
.Y(n_1205)
);

AO21x1_ASAP7_75t_L g1206 ( 
.A1(n_1013),
.A2(n_927),
.B(n_852),
.Y(n_1206)
);

NAND2x1_ASAP7_75t_L g1207 ( 
.A(n_1029),
.B(n_1003),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1152),
.A2(n_840),
.B(n_911),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1198),
.B(n_853),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1059),
.B(n_927),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1082),
.B(n_1097),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1171),
.A2(n_865),
.B(n_863),
.Y(n_1212)
);

O2A1O1Ixp5_ASAP7_75t_L g1213 ( 
.A1(n_1172),
.A2(n_846),
.B(n_851),
.C(n_977),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1171),
.A2(n_865),
.B(n_863),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1139),
.A2(n_1154),
.B(n_1142),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1069),
.A2(n_912),
.B(n_902),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1133),
.B(n_1082),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1152),
.A2(n_840),
.B(n_869),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1077),
.A2(n_925),
.B(n_888),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1170),
.B(n_856),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1162),
.A2(n_879),
.B(n_877),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1170),
.B(n_982),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1053),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1152),
.A2(n_959),
.B(n_940),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1185),
.A2(n_876),
.B1(n_834),
.B2(n_843),
.Y(n_1225)
);

OAI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1183),
.A2(n_882),
.B(n_837),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1060),
.B(n_955),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1104),
.A2(n_958),
.B(n_956),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1144),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1088),
.A2(n_959),
.B(n_940),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1147),
.A2(n_982),
.B1(n_1007),
.B2(n_977),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1060),
.B(n_968),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1144),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1156),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1164),
.A2(n_859),
.A3(n_1001),
.B(n_998),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1120),
.A2(n_845),
.B(n_1003),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1015),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1141),
.Y(n_1238)
);

NAND2xp33_ASAP7_75t_L g1239 ( 
.A(n_1094),
.B(n_1003),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1120),
.A2(n_873),
.B(n_768),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1186),
.A2(n_923),
.B(n_971),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1097),
.B(n_281),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1109),
.A2(n_988),
.B(n_973),
.Y(n_1243)
);

NOR2x1_ASAP7_75t_SL g1244 ( 
.A(n_1094),
.B(n_990),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1121),
.A2(n_994),
.B(n_992),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1180),
.B(n_811),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1180),
.B(n_819),
.Y(n_1247)
);

CKINVDCx6p67_ASAP7_75t_R g1248 ( 
.A(n_1053),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1182),
.B(n_819),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1047),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1094),
.A2(n_768),
.B(n_739),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1028),
.A2(n_937),
.B(n_933),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1185),
.A2(n_449),
.B(n_441),
.C(n_573),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1156),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1182),
.B(n_830),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1158),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1029),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1094),
.A2(n_820),
.B(n_794),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1158),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1022),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1188),
.A2(n_997),
.B(n_830),
.Y(n_1261)
);

OR2x2_ASAP7_75t_L g1262 ( 
.A(n_1066),
.B(n_570),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1034),
.B(n_290),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1029),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1054),
.A2(n_729),
.B(n_685),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1047),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1190),
.B(n_729),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1168),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1201),
.A2(n_1203),
.B(n_1202),
.Y(n_1269)
);

AO22x2_ASAP7_75t_L g1270 ( 
.A1(n_1099),
.A2(n_573),
.B1(n_281),
.B2(n_382),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1147),
.A2(n_1166),
.B(n_1064),
.C(n_1190),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1029),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1204),
.B(n_729),
.Y(n_1273)
);

INVxp67_ASAP7_75t_SL g1274 ( 
.A(n_1029),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1168),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1048),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1018),
.A2(n_740),
.B(n_737),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1204),
.B(n_737),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1140),
.B(n_737),
.Y(n_1279)
);

NAND3xp33_ASAP7_75t_SL g1280 ( 
.A(n_1150),
.B(n_358),
.C(n_357),
.Y(n_1280)
);

AOI21x1_ASAP7_75t_SL g1281 ( 
.A1(n_1114),
.A2(n_831),
.B(n_803),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1140),
.B(n_740),
.Y(n_1282)
);

AO32x2_ASAP7_75t_L g1283 ( 
.A1(n_1021),
.A2(n_826),
.A3(n_820),
.B1(n_794),
.B2(n_803),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1025),
.B(n_382),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1018),
.A2(n_742),
.B(n_740),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1026),
.A2(n_774),
.B(n_742),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1025),
.B(n_382),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1094),
.A2(n_820),
.B(n_794),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1095),
.A2(n_826),
.B(n_777),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1095),
.A2(n_777),
.B(n_736),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1175),
.B(n_1012),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1175),
.B(n_742),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1095),
.A2(n_777),
.B(n_736),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1095),
.A2(n_777),
.B(n_736),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1095),
.A2(n_777),
.B(n_736),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1138),
.A2(n_804),
.B(n_774),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1012),
.B(n_774),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1026),
.A2(n_804),
.B(n_746),
.Y(n_1298)
);

AO31x2_ASAP7_75t_L g1299 ( 
.A1(n_1164),
.A2(n_746),
.A3(n_488),
.B(n_489),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1133),
.B(n_736),
.Y(n_1300)
);

NAND3x1_ASAP7_75t_L g1301 ( 
.A(n_1032),
.B(n_554),
.C(n_548),
.Y(n_1301)
);

AOI211x1_ASAP7_75t_L g1302 ( 
.A1(n_1010),
.A2(n_1023),
.B(n_1039),
.C(n_1011),
.Y(n_1302)
);

BUFx4f_ASAP7_75t_SL g1303 ( 
.A(n_1022),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1141),
.A2(n_804),
.B(n_629),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1022),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1031),
.B(n_624),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1030),
.A2(n_588),
.B(n_582),
.Y(n_1307)
);

O2A1O1Ixp5_ASAP7_75t_L g1308 ( 
.A1(n_1145),
.A2(n_634),
.B(n_624),
.C(n_629),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1030),
.A2(n_588),
.B(n_582),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1103),
.A2(n_795),
.B(n_724),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1031),
.B(n_634),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1078),
.A2(n_644),
.B(n_641),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1184),
.A2(n_487),
.A3(n_488),
.B(n_489),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1081),
.B(n_548),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1036),
.B(n_376),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1024),
.A2(n_795),
.B(n_724),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1033),
.A2(n_588),
.B(n_582),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1114),
.A2(n_776),
.B(n_764),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1191),
.A2(n_795),
.B1(n_266),
.B2(n_298),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1033),
.A2(n_1052),
.B(n_1040),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1048),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1167),
.B(n_362),
.Y(n_1322)
);

BUFx10_ASAP7_75t_L g1323 ( 
.A(n_1034),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_1141),
.Y(n_1324)
);

A2O1A1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1184),
.A2(n_430),
.B(n_386),
.C(n_389),
.Y(n_1325)
);

AO31x2_ASAP7_75t_L g1326 ( 
.A1(n_1148),
.A2(n_487),
.A3(n_494),
.B(n_497),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1115),
.B(n_641),
.Y(n_1327)
);

AND2x6_ASAP7_75t_L g1328 ( 
.A(n_1199),
.B(n_795),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1197),
.A2(n_724),
.B(n_677),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1049),
.A2(n_724),
.B(n_677),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1063),
.A2(n_677),
.B(n_588),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1048),
.A2(n_376),
.B(n_298),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_SL g1333 ( 
.A(n_1133),
.B(n_1048),
.Y(n_1333)
);

AO31x2_ASAP7_75t_L g1334 ( 
.A1(n_1153),
.A2(n_1195),
.A3(n_1067),
.B(n_1020),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_SL g1335 ( 
.A1(n_1063),
.A2(n_497),
.B(n_494),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1080),
.B(n_677),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1115),
.A2(n_776),
.B(n_764),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1174),
.B(n_644),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1040),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1052),
.A2(n_591),
.B(n_582),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1155),
.A2(n_677),
.B(n_591),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1036),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1037),
.B(n_649),
.Y(n_1343)
);

AO21x1_ASAP7_75t_L g1344 ( 
.A1(n_1093),
.A2(n_656),
.B(n_652),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1041),
.B(n_649),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1020),
.B(n_652),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1070),
.A2(n_591),
.B(n_656),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1157),
.A2(n_591),
.B(n_623),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1048),
.A2(n_376),
.B(n_298),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1070),
.A2(n_598),
.B(n_604),
.Y(n_1350)
);

OA21x2_ASAP7_75t_L g1351 ( 
.A1(n_1079),
.A2(n_498),
.B(n_598),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1067),
.B(n_365),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1074),
.B(n_369),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1083),
.B(n_373),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1057),
.A2(n_498),
.A3(n_598),
.B(n_604),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1055),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1177),
.A2(n_623),
.B(n_376),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1086),
.B(n_377),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1126),
.A2(n_417),
.B(n_451),
.C(n_447),
.Y(n_1359)
);

AO21x1_ASAP7_75t_L g1360 ( 
.A1(n_1099),
.A2(n_555),
.B(n_568),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1117),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1056),
.B(n_111),
.Y(n_1362)
);

O2A1O1Ixp5_ASAP7_75t_L g1363 ( 
.A1(n_1111),
.A2(n_1068),
.B(n_1123),
.C(n_1122),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1100),
.A2(n_604),
.B(n_554),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1092),
.A2(n_266),
.B1(n_298),
.B2(n_299),
.Y(n_1365)
);

NAND3xp33_ASAP7_75t_L g1366 ( 
.A(n_1126),
.B(n_415),
.C(n_446),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1100),
.A2(n_565),
.B(n_558),
.Y(n_1367)
);

INVx4_ASAP7_75t_L g1368 ( 
.A(n_1051),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1110),
.A2(n_623),
.B(n_299),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1192),
.A2(n_413),
.B(n_436),
.C(n_433),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1076),
.B(n_1200),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1076),
.B(n_378),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1304),
.A2(n_1119),
.B(n_1107),
.Y(n_1373)
);

INVx2_ASAP7_75t_SL g1374 ( 
.A(n_1223),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_1305),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1339),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1333),
.B(n_1051),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1339),
.Y(n_1378)
);

OAI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1210),
.A2(n_1134),
.B(n_1101),
.Y(n_1379)
);

NOR2x1_ASAP7_75t_SL g1380 ( 
.A(n_1257),
.B(n_1051),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_SL g1381 ( 
.A(n_1371),
.B(n_1090),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1304),
.A2(n_1119),
.B(n_1107),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1234),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1254),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1250),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1333),
.B(n_1051),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1296),
.A2(n_1143),
.B(n_1128),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1210),
.A2(n_1199),
.B(n_1058),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1372),
.A2(n_1132),
.B1(n_1014),
.B2(n_1159),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1211),
.B(n_1227),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1320),
.Y(n_1391)
);

NAND2xp33_ASAP7_75t_R g1392 ( 
.A(n_1371),
.B(n_1046),
.Y(n_1392)
);

INVx5_ASAP7_75t_L g1393 ( 
.A(n_1328),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1361),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1263),
.A2(n_1065),
.B1(n_1113),
.B2(n_1044),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1256),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1296),
.A2(n_1143),
.B(n_1128),
.Y(n_1397)
);

HB1xp67_ASAP7_75t_L g1398 ( 
.A(n_1250),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1208),
.A2(n_1084),
.B(n_1051),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1259),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1362),
.B(n_1056),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1268),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_SL g1403 ( 
.A1(n_1360),
.A2(n_1206),
.B(n_1344),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1363),
.A2(n_1135),
.B(n_1125),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1275),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1372),
.A2(n_1071),
.B1(n_1113),
.B2(n_1081),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1356),
.Y(n_1407)
);

AOI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1225),
.A2(n_1111),
.B(n_1136),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1366),
.A2(n_1132),
.B1(n_1071),
.B2(n_1062),
.Y(n_1409)
);

NAND2x1p5_ASAP7_75t_L g1410 ( 
.A(n_1212),
.B(n_1084),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1227),
.B(n_1043),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1302),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1362),
.B(n_1056),
.Y(n_1413)
);

AO21x1_ASAP7_75t_L g1414 ( 
.A1(n_1319),
.A2(n_1118),
.B(n_1112),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1216),
.A2(n_1149),
.B(n_1179),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1232),
.B(n_1205),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1281),
.A2(n_1096),
.B(n_1146),
.Y(n_1417)
);

INVxp33_ASAP7_75t_L g1418 ( 
.A(n_1242),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1226),
.A2(n_1124),
.B(n_1196),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1281),
.A2(n_1096),
.B(n_1169),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1363),
.A2(n_1091),
.B(n_1112),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1238),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1291),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1214),
.B(n_1084),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1213),
.A2(n_1091),
.B(n_1112),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1265),
.A2(n_1096),
.B(n_1169),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1260),
.A2(n_1019),
.B1(n_1137),
.B2(n_1065),
.Y(n_1427)
);

AO21x2_ASAP7_75t_L g1428 ( 
.A1(n_1269),
.A2(n_1118),
.B(n_1091),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1347),
.A2(n_1298),
.B(n_1307),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1239),
.A2(n_1084),
.B(n_1092),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1237),
.B(n_1016),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1305),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1309),
.A2(n_1194),
.B(n_1169),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1317),
.A2(n_1194),
.B(n_1050),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1232),
.B(n_1042),
.Y(n_1435)
);

OR2x6_ASAP7_75t_L g1436 ( 
.A(n_1217),
.B(n_1036),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1257),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1223),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1229),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1340),
.A2(n_1194),
.B(n_1050),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1241),
.A2(n_1118),
.B(n_1129),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1217),
.A2(n_1161),
.B1(n_1062),
.B2(n_1089),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1280),
.A2(n_1062),
.B1(n_1043),
.B2(n_1075),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1239),
.A2(n_1084),
.B(n_1108),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1362),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1233),
.Y(n_1446)
);

INVxp67_ASAP7_75t_L g1447 ( 
.A(n_1266),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1322),
.B(n_1044),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1271),
.A2(n_1066),
.B(n_1110),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1257),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1314),
.Y(n_1451)
);

AOI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1300),
.A2(n_1080),
.B(n_1116),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1271),
.A2(n_1116),
.B(n_1151),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1213),
.A2(n_558),
.B(n_555),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1238),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1342),
.B(n_1073),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1219),
.A2(n_1127),
.B(n_1160),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1277),
.A2(n_1050),
.B(n_1105),
.Y(n_1458)
);

CKINVDCx12_ASAP7_75t_R g1459 ( 
.A(n_1315),
.Y(n_1459)
);

AO31x2_ASAP7_75t_L g1460 ( 
.A1(n_1253),
.A2(n_1193),
.A3(n_1131),
.B(n_1187),
.Y(n_1460)
);

AO21x1_ASAP7_75t_L g1461 ( 
.A1(n_1365),
.A2(n_1300),
.B(n_1220),
.Y(n_1461)
);

NAND2x1_ASAP7_75t_L g1462 ( 
.A(n_1328),
.B(n_1108),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1324),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1222),
.A2(n_1131),
.B1(n_1075),
.B2(n_1073),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1285),
.A2(n_559),
.B(n_562),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1209),
.B(n_1161),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1338),
.Y(n_1467)
);

AO31x2_ASAP7_75t_L g1468 ( 
.A1(n_1253),
.A2(n_1193),
.A3(n_1108),
.B(n_1187),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1324),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1236),
.A2(n_1178),
.B(n_1187),
.Y(n_1470)
);

AO31x2_ASAP7_75t_L g1471 ( 
.A1(n_1312),
.A2(n_1193),
.A3(n_1178),
.B(n_559),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1346),
.Y(n_1472)
);

OAI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1231),
.A2(n_1038),
.B1(n_1130),
.B2(n_1085),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1262),
.B(n_1161),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1248),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1286),
.A2(n_568),
.B(n_565),
.Y(n_1476)
);

NAND2x1p5_ASAP7_75t_L g1477 ( 
.A(n_1342),
.B(n_1178),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1322),
.A2(n_1061),
.B1(n_1035),
.B2(n_1087),
.C(n_1019),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1315),
.B(n_1036),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1306),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1266),
.B(n_1165),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1311),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1303),
.A2(n_1045),
.B1(n_1017),
.B2(n_1027),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1261),
.A2(n_562),
.B(n_1181),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1252),
.A2(n_1181),
.B(n_1173),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1350),
.A2(n_1181),
.B(n_1173),
.Y(n_1486)
);

HB1xp67_ASAP7_75t_L g1487 ( 
.A(n_1284),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1357),
.A2(n_1098),
.B(n_1181),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1287),
.A2(n_1163),
.B1(n_1038),
.B2(n_1130),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1303),
.A2(n_1045),
.B1(n_1017),
.B2(n_1027),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1343),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1231),
.A2(n_1163),
.B1(n_1038),
.B2(n_1072),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1367),
.Y(n_1493)
);

BUFx2_ASAP7_75t_R g1494 ( 
.A(n_1353),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1257),
.B(n_1098),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1221),
.A2(n_1181),
.B(n_1173),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1364),
.A2(n_1215),
.B(n_1240),
.Y(n_1497)
);

NAND3xp33_ASAP7_75t_L g1498 ( 
.A(n_1359),
.B(n_1163),
.C(n_385),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1218),
.A2(n_1173),
.B(n_1098),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1323),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1334),
.B(n_1165),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1230),
.A2(n_1173),
.B(n_1102),
.Y(n_1502)
);

AOI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1348),
.A2(n_1163),
.B(n_1102),
.Y(n_1503)
);

AO31x2_ASAP7_75t_L g1504 ( 
.A1(n_1325),
.A2(n_1102),
.A3(n_1098),
.B(n_1189),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1323),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1299),
.Y(n_1506)
);

AOI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1327),
.A2(n_1102),
.B(n_1098),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1345),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1352),
.B(n_1359),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1274),
.A2(n_1038),
.B1(n_1085),
.B2(n_1072),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1341),
.A2(n_1102),
.B(n_1189),
.Y(n_1511)
);

OAI21x1_ASAP7_75t_L g1512 ( 
.A1(n_1329),
.A2(n_1176),
.B(n_776),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1228),
.A2(n_1245),
.B(n_1243),
.Y(n_1513)
);

AOI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1354),
.A2(n_1176),
.B1(n_383),
.B2(n_384),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1308),
.A2(n_776),
.B(n_764),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1299),
.Y(n_1516)
);

OAI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1274),
.A2(n_1137),
.B1(n_408),
.B2(n_391),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1323),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1246),
.A2(n_419),
.B1(n_397),
.B2(n_416),
.Y(n_1519)
);

AOI221x1_ASAP7_75t_L g1520 ( 
.A1(n_1270),
.A2(n_404),
.B1(n_299),
.B2(n_298),
.C(n_623),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1264),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1358),
.B(n_395),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1299),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1325),
.B(n_423),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1276),
.B(n_1368),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1308),
.A2(n_776),
.B(n_764),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1335),
.A2(n_776),
.B(n_764),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1247),
.B(n_764),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_L g1529 ( 
.A1(n_1310),
.A2(n_404),
.B(n_299),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1299),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1251),
.A2(n_404),
.B(n_299),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1264),
.Y(n_1532)
);

CKINVDCx6p67_ASAP7_75t_R g1533 ( 
.A(n_1260),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_SL g1534 ( 
.A(n_1370),
.B(n_290),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1258),
.A2(n_404),
.B(n_299),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1264),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1288),
.A2(n_404),
.B(n_298),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1289),
.A2(n_404),
.B(n_623),
.Y(n_1538)
);

BUFx12f_ASAP7_75t_L g1539 ( 
.A(n_1315),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1326),
.Y(n_1540)
);

AOI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1224),
.A2(n_623),
.B(n_172),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1270),
.A2(n_623),
.B1(n_21),
.B2(n_22),
.Y(n_1542)
);

OA21x2_ASAP7_75t_L g1543 ( 
.A1(n_1369),
.A2(n_1249),
.B(n_1255),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1334),
.B(n_113),
.Y(n_1544)
);

A2O1A1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1370),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1326),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1326),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1331),
.A2(n_229),
.B(n_220),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1267),
.A2(n_25),
.B(n_26),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1290),
.A2(n_214),
.B(n_211),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1334),
.B(n_25),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1301),
.A2(n_1328),
.B1(n_1279),
.B2(n_1282),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1293),
.A2(n_1294),
.B(n_1295),
.Y(n_1553)
);

O2A1O1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1273),
.A2(n_26),
.B(n_28),
.C(n_29),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1316),
.A2(n_210),
.B(n_206),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1264),
.Y(n_1556)
);

NAND2xp33_ASAP7_75t_L g1557 ( 
.A(n_1416),
.B(n_1328),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1376),
.Y(n_1558)
);

AO31x2_ASAP7_75t_L g1559 ( 
.A1(n_1461),
.A2(n_1244),
.A3(n_1283),
.B(n_1278),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1383),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1384),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1385),
.Y(n_1562)
);

INVx3_ASAP7_75t_SL g1563 ( 
.A(n_1518),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1415),
.A2(n_1470),
.B(n_1393),
.Y(n_1564)
);

INVx6_ASAP7_75t_L g1565 ( 
.A(n_1500),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1475),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_R g1567 ( 
.A(n_1392),
.B(n_1272),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1390),
.B(n_1334),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1542),
.A2(n_1328),
.B1(n_1292),
.B2(n_1301),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1406),
.A2(n_1297),
.B1(n_1276),
.B2(n_1368),
.Y(n_1570)
);

NAND2x1p5_ASAP7_75t_L g1571 ( 
.A(n_1393),
.B(n_1272),
.Y(n_1571)
);

NOR2xp33_ASAP7_75t_L g1572 ( 
.A(n_1448),
.B(n_1321),
.Y(n_1572)
);

INVx2_ASAP7_75t_SL g1573 ( 
.A(n_1475),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1436),
.B(n_1332),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1394),
.Y(n_1575)
);

OAI21xp33_ASAP7_75t_L g1576 ( 
.A1(n_1435),
.A2(n_1349),
.B(n_1337),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1518),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1509),
.A2(n_1318),
.B(n_1330),
.Y(n_1578)
);

OAI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1520),
.A2(n_1272),
.B1(n_1207),
.B2(n_1336),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1451),
.B(n_1313),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1407),
.Y(n_1581)
);

OAI21x1_ASAP7_75t_SL g1582 ( 
.A1(n_1453),
.A2(n_1351),
.B(n_1313),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1418),
.B(n_1313),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1400),
.Y(n_1584)
);

OAI222xp33_ASAP7_75t_L g1585 ( 
.A1(n_1492),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.C1(n_37),
.C2(n_39),
.Y(n_1585)
);

AOI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1478),
.A2(n_1235),
.B1(n_1313),
.B2(n_1283),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1418),
.B(n_1487),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1481),
.B(n_1235),
.Y(n_1588)
);

CKINVDCx8_ASAP7_75t_R g1589 ( 
.A(n_1375),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1415),
.A2(n_1283),
.B(n_1235),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1481),
.B(n_1235),
.Y(n_1591)
);

NAND2xp33_ASAP7_75t_R g1592 ( 
.A(n_1425),
.B(n_1283),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1402),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1405),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1398),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1389),
.A2(n_1355),
.B1(n_33),
.B2(n_37),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1379),
.A2(n_31),
.B(n_39),
.C(n_40),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1376),
.Y(n_1598)
);

OAI21x1_ASAP7_75t_L g1599 ( 
.A1(n_1496),
.A2(n_1355),
.B(n_200),
.Y(n_1599)
);

INVx2_ASAP7_75t_SL g1600 ( 
.A(n_1505),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_L g1601 ( 
.A1(n_1467),
.A2(n_42),
.B1(n_46),
.B2(n_48),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1411),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1491),
.B(n_1355),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1388),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1396),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_R g1606 ( 
.A(n_1425),
.B(n_196),
.Y(n_1606)
);

BUFx6f_ASAP7_75t_L g1607 ( 
.A(n_1556),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1443),
.A2(n_1355),
.B1(n_57),
.B2(n_59),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1508),
.B(n_56),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1401),
.B(n_187),
.Y(n_1610)
);

AO31x2_ASAP7_75t_L g1611 ( 
.A1(n_1461),
.A2(n_56),
.A3(n_57),
.B(n_59),
.Y(n_1611)
);

AOI221xp5_ASAP7_75t_L g1612 ( 
.A1(n_1395),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.C(n_65),
.Y(n_1612)
);

BUFx6f_ASAP7_75t_L g1613 ( 
.A(n_1556),
.Y(n_1613)
);

AOI221xp5_ASAP7_75t_L g1614 ( 
.A1(n_1554),
.A2(n_60),
.B1(n_62),
.B2(n_68),
.C(n_70),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1472),
.A2(n_68),
.B1(n_71),
.B2(n_73),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1436),
.B(n_1479),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1415),
.A2(n_184),
.B(n_179),
.Y(n_1617)
);

AO21x2_ASAP7_75t_L g1618 ( 
.A1(n_1403),
.A2(n_173),
.B(n_166),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1498),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1378),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1449),
.B(n_76),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1375),
.Y(n_1622)
);

BUFx3_ASAP7_75t_L g1623 ( 
.A(n_1505),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_SL g1624 ( 
.A1(n_1427),
.A2(n_77),
.B1(n_79),
.B2(n_81),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1474),
.B(n_82),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1378),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1422),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1422),
.Y(n_1628)
);

NAND2x1p5_ASAP7_75t_L g1629 ( 
.A(n_1393),
.B(n_127),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1455),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1428),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1496),
.A2(n_124),
.B(n_158),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1480),
.A2(n_83),
.B1(n_85),
.B2(n_89),
.Y(n_1633)
);

OAI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1482),
.A2(n_83),
.B1(n_85),
.B2(n_89),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1439),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1446),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1457),
.A2(n_91),
.B1(n_93),
.B2(n_95),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1374),
.Y(n_1638)
);

NOR2xp67_ASAP7_75t_SL g1639 ( 
.A(n_1500),
.B(n_95),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1545),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.C(n_102),
.Y(n_1640)
);

INVx4_ASAP7_75t_L g1641 ( 
.A(n_1456),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1457),
.A2(n_96),
.B1(n_101),
.B2(n_161),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1423),
.B(n_128),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1457),
.A2(n_156),
.B1(n_130),
.B2(n_132),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1466),
.B(n_129),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1428),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1463),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1525),
.Y(n_1648)
);

OR2x6_ASAP7_75t_L g1649 ( 
.A(n_1436),
.B(n_133),
.Y(n_1649)
);

OAI22xp33_ASAP7_75t_L g1650 ( 
.A1(n_1501),
.A2(n_1442),
.B1(n_1393),
.B2(n_1445),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1469),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1522),
.A2(n_145),
.B1(n_148),
.B2(n_1524),
.C(n_1545),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1381),
.B(n_1401),
.Y(n_1653)
);

AO21x2_ASAP7_75t_L g1654 ( 
.A1(n_1403),
.A2(n_1513),
.B(n_1408),
.Y(n_1654)
);

INVx4_ASAP7_75t_L g1655 ( 
.A(n_1456),
.Y(n_1655)
);

AND2x4_ASAP7_75t_L g1656 ( 
.A(n_1401),
.B(n_1413),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1489),
.B(n_1409),
.C(n_1514),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1393),
.A2(n_1399),
.B(n_1430),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1445),
.A2(n_1473),
.B1(n_1431),
.B2(n_1494),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_SL g1660 ( 
.A(n_1534),
.B(n_1483),
.C(n_1490),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1417),
.Y(n_1661)
);

CKINVDCx16_ASAP7_75t_R g1662 ( 
.A(n_1539),
.Y(n_1662)
);

INVx1_ASAP7_75t_SL g1663 ( 
.A(n_1374),
.Y(n_1663)
);

INVx3_ASAP7_75t_L g1664 ( 
.A(n_1525),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1441),
.A2(n_1551),
.B1(n_1501),
.B2(n_1414),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1445),
.A2(n_1552),
.B1(n_1510),
.B2(n_1413),
.Y(n_1666)
);

OR2x6_ASAP7_75t_L g1667 ( 
.A(n_1436),
.B(n_1479),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1413),
.B(n_1447),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1445),
.A2(n_1464),
.B1(n_1456),
.B2(n_1438),
.Y(n_1669)
);

INVx4_ASAP7_75t_L g1670 ( 
.A(n_1556),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1412),
.Y(n_1671)
);

NAND2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1438),
.B(n_1432),
.Y(n_1672)
);

INVx4_ASAP7_75t_SL g1673 ( 
.A(n_1460),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1551),
.Y(n_1674)
);

A2O1A1Ixp33_ASAP7_75t_L g1675 ( 
.A1(n_1544),
.A2(n_1541),
.B(n_1550),
.C(n_1444),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1556),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1517),
.B(n_1519),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1441),
.B(n_1544),
.Y(n_1678)
);

INVx4_ASAP7_75t_L g1679 ( 
.A(n_1556),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1441),
.B(n_1428),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1506),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1513),
.A2(n_1408),
.B(n_1497),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1414),
.B(n_1377),
.Y(n_1683)
);

NAND3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1432),
.B(n_1386),
.C(n_1377),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1419),
.A2(n_1549),
.B1(n_1539),
.B2(n_1533),
.Y(n_1685)
);

BUFx3_ASAP7_75t_L g1686 ( 
.A(n_1525),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1419),
.A2(n_1546),
.B1(n_1547),
.B2(n_1540),
.C(n_1530),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1533),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_SL g1689 ( 
.A1(n_1419),
.A2(n_1549),
.B1(n_1425),
.B2(n_1479),
.Y(n_1689)
);

OAI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1499),
.A2(n_1417),
.B(n_1502),
.Y(n_1690)
);

AOI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1549),
.A2(n_1421),
.B1(n_1530),
.B2(n_1516),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1479),
.A2(n_1377),
.B1(n_1386),
.B2(n_1421),
.C(n_1528),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1462),
.B(n_1386),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1495),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1516),
.Y(n_1695)
);

OR2x2_ASAP7_75t_L g1696 ( 
.A(n_1437),
.B(n_1536),
.Y(n_1696)
);

AOI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1421),
.A2(n_1523),
.B1(n_1540),
.B2(n_1404),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_L g1698 ( 
.A(n_1477),
.B(n_1532),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1468),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1477),
.A2(n_1462),
.B1(n_1503),
.B2(n_1495),
.Y(n_1700)
);

OAI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1477),
.A2(n_1503),
.B1(n_1495),
.B2(n_1437),
.Y(n_1701)
);

OAI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1543),
.A2(n_1404),
.B1(n_1521),
.B2(n_1450),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1536),
.B(n_1532),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1404),
.Y(n_1704)
);

BUFx12f_ASAP7_75t_L g1705 ( 
.A(n_1450),
.Y(n_1705)
);

AOI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1543),
.A2(n_1484),
.B1(n_1548),
.B2(n_1454),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1521),
.B(n_1380),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1460),
.B(n_1468),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1460),
.B(n_1504),
.Y(n_1709)
);

NAND2xp33_ASAP7_75t_R g1710 ( 
.A(n_1543),
.B(n_1454),
.Y(n_1710)
);

AOI22xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1550),
.A2(n_1548),
.B1(n_1555),
.B2(n_1484),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1484),
.A2(n_1493),
.B1(n_1391),
.B2(n_1410),
.C(n_1424),
.Y(n_1712)
);

AND2x2_ASAP7_75t_SL g1713 ( 
.A(n_1454),
.B(n_1459),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1420),
.Y(n_1714)
);

OAI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1452),
.A2(n_1391),
.B1(n_1459),
.B2(n_1507),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1458),
.B(n_1468),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1507),
.A2(n_1452),
.B1(n_1424),
.B2(n_1410),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1460),
.B(n_1504),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1504),
.B(n_1471),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1420),
.Y(n_1720)
);

CKINVDCx5p33_ASAP7_75t_R g1721 ( 
.A(n_1493),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1488),
.B(n_1527),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1458),
.Y(n_1723)
);

OAI21xp33_ASAP7_75t_L g1724 ( 
.A1(n_1555),
.A2(n_1424),
.B(n_1410),
.Y(n_1724)
);

BUFx10_ASAP7_75t_L g1725 ( 
.A(n_1471),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_SL g1726 ( 
.A1(n_1531),
.A2(n_1537),
.B1(n_1535),
.B2(n_1527),
.Y(n_1726)
);

OR2x6_ASAP7_75t_L g1727 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1488),
.A2(n_1527),
.B1(n_1387),
.B2(n_1397),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1468),
.B(n_1504),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1504),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1468),
.A2(n_1471),
.B1(n_1485),
.B2(n_1488),
.Y(n_1731)
);

INVx6_ASAP7_75t_L g1732 ( 
.A(n_1511),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1471),
.B(n_1529),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1387),
.A2(n_1397),
.B1(n_1373),
.B2(n_1382),
.Y(n_1734)
);

AND2x2_ASAP7_75t_SL g1735 ( 
.A(n_1471),
.B(n_1537),
.Y(n_1735)
);

INVx4_ASAP7_75t_L g1736 ( 
.A(n_1434),
.Y(n_1736)
);

BUFx12f_ASAP7_75t_L g1737 ( 
.A(n_1529),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1512),
.A2(n_1553),
.B1(n_1426),
.B2(n_1434),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1433),
.Y(n_1739)
);

NAND2x1_ASAP7_75t_L g1740 ( 
.A(n_1433),
.B(n_1440),
.Y(n_1740)
);

OAI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1512),
.A2(n_1526),
.B1(n_1515),
.B2(n_1531),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1465),
.B(n_1476),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1426),
.B(n_1440),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1465),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1476),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_1553),
.Y(n_1746)
);

INVx3_ASAP7_75t_L g1747 ( 
.A(n_1486),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1535),
.A2(n_1497),
.B1(n_1515),
.B2(n_1526),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1612),
.A2(n_1429),
.B1(n_1486),
.B2(n_1538),
.C(n_1602),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1668),
.B(n_1538),
.Y(n_1750)
);

AOI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1660),
.A2(n_1657),
.B1(n_1659),
.B2(n_1677),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1605),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1653),
.B(n_1583),
.Y(n_1753)
);

OR2x6_ASAP7_75t_L g1754 ( 
.A(n_1616),
.B(n_1667),
.Y(n_1754)
);

OA21x2_ASAP7_75t_L g1755 ( 
.A1(n_1590),
.A2(n_1706),
.B(n_1734),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1624),
.A2(n_1604),
.B1(n_1619),
.B2(n_1572),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1561),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1621),
.A2(n_1614),
.B1(n_1604),
.B2(n_1637),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1619),
.A2(n_1572),
.B1(n_1637),
.B2(n_1642),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1588),
.B(n_1591),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1625),
.A2(n_1639),
.B1(n_1666),
.B2(n_1610),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1575),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1625),
.A2(n_1610),
.B1(n_1672),
.B2(n_1602),
.Y(n_1763)
);

OAI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1597),
.A2(n_1569),
.B1(n_1563),
.B2(n_1601),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1631),
.Y(n_1765)
);

AO31x2_ASAP7_75t_L g1766 ( 
.A1(n_1731),
.A2(n_1717),
.A3(n_1564),
.B(n_1745),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1634),
.A2(n_1649),
.B1(n_1606),
.B2(n_1596),
.Y(n_1767)
);

INVx2_ASAP7_75t_SL g1768 ( 
.A(n_1565),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1584),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_SL g1770 ( 
.A1(n_1608),
.A2(n_1649),
.B1(n_1678),
.B2(n_1567),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1569),
.A2(n_1563),
.B1(n_1601),
.B2(n_1644),
.Y(n_1771)
);

AOI22xp33_ASAP7_75t_L g1772 ( 
.A1(n_1615),
.A2(n_1633),
.B1(n_1634),
.B2(n_1644),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1627),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1615),
.A2(n_1633),
.B1(n_1609),
.B2(n_1649),
.Y(n_1774)
);

OAI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1606),
.A2(n_1586),
.B1(n_1585),
.B2(n_1650),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1640),
.A2(n_1675),
.B1(n_1576),
.B2(n_1617),
.C(n_1645),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1631),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1581),
.A2(n_1674),
.B1(n_1595),
.B2(n_1568),
.Y(n_1778)
);

NAND3xp33_ASAP7_75t_L g1779 ( 
.A(n_1685),
.B(n_1675),
.C(n_1643),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1567),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1646),
.Y(n_1781)
);

OAI21xp33_ASAP7_75t_L g1782 ( 
.A1(n_1665),
.A2(n_1685),
.B(n_1680),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1593),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1594),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_SL g1785 ( 
.A1(n_1688),
.A2(n_1577),
.B1(n_1623),
.B2(n_1662),
.Y(n_1785)
);

AOI222xp33_ASAP7_75t_L g1786 ( 
.A1(n_1562),
.A2(n_1650),
.B1(n_1665),
.B2(n_1580),
.C1(n_1635),
.C2(n_1636),
.Y(n_1786)
);

AOI221xp5_ASAP7_75t_L g1787 ( 
.A1(n_1578),
.A2(n_1570),
.B1(n_1683),
.B2(n_1669),
.C(n_1692),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1656),
.B(n_1641),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1658),
.A2(n_1579),
.B(n_1698),
.Y(n_1789)
);

AOI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1740),
.A2(n_1700),
.B(n_1701),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1557),
.A2(n_1656),
.B1(n_1618),
.B2(n_1671),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1589),
.A2(n_1573),
.B1(n_1566),
.B2(n_1565),
.Y(n_1792)
);

INVx2_ASAP7_75t_SL g1793 ( 
.A(n_1565),
.Y(n_1793)
);

AOI222xp33_ASAP7_75t_L g1794 ( 
.A1(n_1622),
.A2(n_1663),
.B1(n_1683),
.B2(n_1651),
.C1(n_1566),
.C2(n_1603),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1623),
.A2(n_1600),
.B1(n_1638),
.B2(n_1655),
.Y(n_1795)
);

AOI33xp33_ASAP7_75t_L g1796 ( 
.A1(n_1689),
.A2(n_1719),
.A3(n_1691),
.B1(n_1702),
.B2(n_1709),
.B3(n_1715),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1628),
.Y(n_1797)
);

OAI21x1_ASAP7_75t_L g1798 ( 
.A1(n_1690),
.A2(n_1599),
.B(n_1632),
.Y(n_1798)
);

OAI222xp33_ASAP7_75t_L g1799 ( 
.A1(n_1616),
.A2(n_1667),
.B1(n_1629),
.B2(n_1574),
.C1(n_1641),
.C2(n_1655),
.Y(n_1799)
);

OAI22xp5_ASAP7_75t_L g1800 ( 
.A1(n_1721),
.A2(n_1667),
.B1(n_1616),
.B2(n_1570),
.Y(n_1800)
);

A2O1A1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1724),
.A2(n_1746),
.B(n_1684),
.C(n_1711),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1618),
.A2(n_1582),
.B1(n_1629),
.B2(n_1574),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1574),
.A2(n_1626),
.B1(n_1664),
.B2(n_1648),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1664),
.B(n_1630),
.Y(n_1804)
);

INVx3_ASAP7_75t_SL g1805 ( 
.A(n_1703),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_L g1806 ( 
.A1(n_1734),
.A2(n_1739),
.B(n_1744),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1706),
.A2(n_1687),
.B(n_1691),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1696),
.B(n_1647),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_1705),
.Y(n_1809)
);

AO31x2_ASAP7_75t_L g1810 ( 
.A1(n_1744),
.A2(n_1661),
.A3(n_1704),
.B(n_1723),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1558),
.B(n_1620),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1558),
.A2(n_1620),
.B1(n_1598),
.B2(n_1735),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1598),
.A2(n_1735),
.B1(n_1737),
.B2(n_1730),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_1607),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1646),
.A2(n_1699),
.B1(n_1713),
.B2(n_1695),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1693),
.A2(n_1571),
.B1(n_1718),
.B2(n_1707),
.Y(n_1816)
);

INVx3_ASAP7_75t_L g1817 ( 
.A(n_1670),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1693),
.A2(n_1571),
.B1(n_1707),
.B2(n_1708),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1726),
.A2(n_1738),
.B1(n_1748),
.B2(n_1712),
.C(n_1733),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1613),
.B(n_1676),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1748),
.A2(n_1722),
.B1(n_1728),
.B2(n_1729),
.C(n_1693),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1681),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1694),
.A2(n_1699),
.B1(n_1697),
.B2(n_1679),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1670),
.B(n_1679),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1613),
.B(n_1676),
.Y(n_1825)
);

BUFx4f_ASAP7_75t_SL g1826 ( 
.A(n_1613),
.Y(n_1826)
);

AOI22xp33_ASAP7_75t_SL g1827 ( 
.A1(n_1732),
.A2(n_1694),
.B1(n_1716),
.B2(n_1613),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1695),
.A2(n_1694),
.B1(n_1725),
.B2(n_1654),
.Y(n_1828)
);

O2A1O1Ixp33_ASAP7_75t_SL g1829 ( 
.A1(n_1715),
.A2(n_1741),
.B(n_1720),
.C(n_1702),
.Y(n_1829)
);

OR2x6_ASAP7_75t_L g1830 ( 
.A(n_1716),
.B(n_1727),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1741),
.A2(n_1697),
.B1(n_1728),
.B2(n_1704),
.C(n_1743),
.Y(n_1831)
);

OAI211xp5_ASAP7_75t_SL g1832 ( 
.A1(n_1739),
.A2(n_1714),
.B(n_1747),
.C(n_1611),
.Y(n_1832)
);

OAI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1732),
.A2(n_1736),
.B1(n_1727),
.B2(n_1710),
.C(n_1592),
.Y(n_1833)
);

OAI211xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1747),
.A2(n_1611),
.B(n_1725),
.C(n_1673),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1694),
.A2(n_1732),
.B1(n_1676),
.B2(n_1727),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1736),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1654),
.A2(n_1673),
.B1(n_1742),
.B2(n_1743),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1682),
.A2(n_1710),
.B(n_1592),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1611),
.B(n_1559),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1611),
.Y(n_1840)
);

OAI221xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1673),
.A2(n_1059),
.B1(n_687),
.B2(n_1619),
.C(n_1099),
.Y(n_1841)
);

A2O1A1Ixp33_ASAP7_75t_L g1842 ( 
.A1(n_1559),
.A2(n_1059),
.B(n_907),
.C(n_1210),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1559),
.A2(n_1682),
.B1(n_1059),
.B2(n_1624),
.Y(n_1843)
);

CKINVDCx5p33_ASAP7_75t_R g1844 ( 
.A(n_1577),
.Y(n_1844)
);

BUFx12f_ASAP7_75t_L g1845 ( 
.A(n_1688),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1657),
.A2(n_1059),
.B1(n_1093),
.B2(n_1150),
.Y(n_1847)
);

AOI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1660),
.A2(n_1059),
.B1(n_907),
.B2(n_1093),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1849)
);

AOI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1560),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1581),
.Y(n_1852)
);

AOI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1612),
.A2(n_874),
.B1(n_907),
.B2(n_1059),
.C(n_687),
.Y(n_1853)
);

AOI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1658),
.A2(n_1013),
.B(n_1239),
.Y(n_1854)
);

AO31x2_ASAP7_75t_L g1855 ( 
.A1(n_1731),
.A2(n_1520),
.A3(n_1717),
.B(n_1461),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1560),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1560),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1659),
.B(n_1133),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1657),
.A2(n_1059),
.B1(n_1371),
.B2(n_1406),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1577),
.Y(n_1860)
);

OAI21xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1624),
.A2(n_1059),
.B(n_907),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1625),
.B(n_1371),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1641),
.Y(n_1864)
);

NAND3xp33_ASAP7_75t_L g1865 ( 
.A(n_1619),
.B(n_1059),
.C(n_907),
.Y(n_1865)
);

OAI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1652),
.A2(n_907),
.B(n_1059),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1625),
.B(n_1390),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1868)
);

OA21x2_ASAP7_75t_L g1869 ( 
.A1(n_1590),
.A2(n_1706),
.B(n_1513),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1577),
.Y(n_1871)
);

OAI211xp5_ASAP7_75t_L g1872 ( 
.A1(n_1637),
.A2(n_1059),
.B(n_907),
.C(n_673),
.Y(n_1872)
);

AOI22xp33_ASAP7_75t_L g1873 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1873)
);

NAND2x1p5_ASAP7_75t_L g1874 ( 
.A(n_1621),
.B(n_1393),
.Y(n_1874)
);

OAI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1657),
.A2(n_1059),
.B1(n_1371),
.B2(n_1406),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1612),
.A2(n_874),
.B1(n_907),
.B2(n_1059),
.C(n_687),
.Y(n_1876)
);

NAND4xp25_ASAP7_75t_L g1877 ( 
.A(n_1637),
.B(n_615),
.C(n_874),
.D(n_1059),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1674),
.B(n_1588),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1625),
.B(n_1371),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1650),
.B(n_1210),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1560),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1883)
);

AOI22xp33_ASAP7_75t_L g1884 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1612),
.A2(n_874),
.B1(n_907),
.B2(n_1059),
.C(n_687),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1625),
.B(n_1390),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1658),
.A2(n_1013),
.B(n_1239),
.Y(n_1888)
);

OAI211xp5_ASAP7_75t_L g1889 ( 
.A1(n_1637),
.A2(n_1059),
.B(n_907),
.C(n_673),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1631),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1560),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_L g1892 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1560),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1657),
.A2(n_1059),
.B1(n_1093),
.B2(n_1150),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1895)
);

AOI221xp5_ASAP7_75t_L g1896 ( 
.A1(n_1612),
.A2(n_874),
.B1(n_907),
.B2(n_1059),
.C(n_687),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1686),
.B(n_1648),
.Y(n_1897)
);

INVx2_ASAP7_75t_SL g1898 ( 
.A(n_1565),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_SL g1899 ( 
.A1(n_1657),
.A2(n_1059),
.B1(n_1093),
.B2(n_1150),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_L g1900 ( 
.A1(n_1658),
.A2(n_1013),
.B(n_1239),
.Y(n_1900)
);

OAI21x1_ASAP7_75t_L g1901 ( 
.A1(n_1564),
.A2(n_1513),
.B(n_1497),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1660),
.A2(n_1059),
.B1(n_907),
.B2(n_1093),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1560),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1905)
);

BUFx12f_ASAP7_75t_L g1906 ( 
.A(n_1688),
.Y(n_1906)
);

AOI221xp5_ASAP7_75t_L g1907 ( 
.A1(n_1612),
.A2(n_874),
.B1(n_907),
.B2(n_1059),
.C(n_687),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_L g1908 ( 
.A1(n_1621),
.A2(n_1150),
.B1(n_1126),
.B2(n_1059),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1668),
.B(n_1587),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1863),
.B(n_1868),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1810),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1810),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1822),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1810),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1805),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1760),
.B(n_1753),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1879),
.B(n_1878),
.Y(n_1918)
);

INVx2_ASAP7_75t_SL g1919 ( 
.A(n_1805),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1765),
.B(n_1777),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1865),
.A2(n_1853),
.B1(n_1896),
.B2(n_1885),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1895),
.B(n_1909),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1779),
.B(n_1836),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1810),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1910),
.Y(n_1925)
);

AO21x2_ASAP7_75t_L g1926 ( 
.A1(n_1842),
.A2(n_1838),
.B(n_1840),
.Y(n_1926)
);

INVx3_ASAP7_75t_SL g1927 ( 
.A(n_1785),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1830),
.B(n_1815),
.Y(n_1928)
);

BUFx2_ASAP7_75t_L g1929 ( 
.A(n_1830),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1830),
.B(n_1815),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1806),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1808),
.B(n_1867),
.Y(n_1932)
);

AO21x2_ASAP7_75t_L g1933 ( 
.A1(n_1829),
.A2(n_1789),
.B(n_1901),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1765),
.B(n_1777),
.Y(n_1934)
);

AOI222xp33_ASAP7_75t_L g1935 ( 
.A1(n_1876),
.A2(n_1907),
.B1(n_1756),
.B2(n_1759),
.C1(n_1758),
.C2(n_1772),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1886),
.B(n_1862),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1781),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1757),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1812),
.B(n_1762),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1862),
.B(n_1880),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1754),
.B(n_1836),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1754),
.B(n_1790),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1769),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1880),
.B(n_1778),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1812),
.B(n_1783),
.Y(n_1945)
);

OAI21xp33_ASAP7_75t_SL g1946 ( 
.A1(n_1881),
.A2(n_1877),
.B(n_1772),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1784),
.B(n_1851),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1856),
.B(n_1857),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1882),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1891),
.B(n_1893),
.Y(n_1950)
);

BUFx2_ASAP7_75t_L g1951 ( 
.A(n_1754),
.Y(n_1951)
);

HB1xp67_ASAP7_75t_L g1952 ( 
.A(n_1781),
.Y(n_1952)
);

INVx2_ASAP7_75t_L g1953 ( 
.A(n_1903),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1796),
.B(n_1837),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1837),
.B(n_1813),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1813),
.B(n_1782),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1807),
.B(n_1828),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1798),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1807),
.B(n_1828),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1778),
.B(n_1752),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1890),
.Y(n_1961)
);

INVx2_ASAP7_75t_L g1962 ( 
.A(n_1869),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1869),
.Y(n_1963)
);

BUFx8_ASAP7_75t_L g1964 ( 
.A(n_1845),
.Y(n_1964)
);

BUFx2_ASAP7_75t_L g1965 ( 
.A(n_1835),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1839),
.B(n_1833),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1807),
.B(n_1750),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1831),
.B(n_1755),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1766),
.B(n_1755),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1755),
.B(n_1787),
.Y(n_1970)
);

OAI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1758),
.A2(n_1774),
.B1(n_1905),
.B2(n_1887),
.Y(n_1971)
);

OR2x2_ASAP7_75t_L g1972 ( 
.A(n_1766),
.B(n_1821),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1811),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1855),
.B(n_1786),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1751),
.B(n_1852),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1766),
.B(n_1801),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1855),
.B(n_1766),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1859),
.B(n_1875),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1855),
.B(n_1820),
.Y(n_1979)
);

AOI22xp33_ASAP7_75t_SL g1980 ( 
.A1(n_1872),
.A2(n_1889),
.B1(n_1771),
.B2(n_1764),
.Y(n_1980)
);

A2O1A1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1861),
.A2(n_1848),
.B(n_1902),
.C(n_1866),
.Y(n_1981)
);

HB1xp67_ASAP7_75t_L g1982 ( 
.A(n_1804),
.Y(n_1982)
);

INVx2_ASAP7_75t_L g1983 ( 
.A(n_1869),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1794),
.B(n_1881),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1773),
.B(n_1797),
.Y(n_1985)
);

CKINVDCx5p33_ASAP7_75t_R g1986 ( 
.A(n_1844),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1855),
.B(n_1823),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1803),
.B(n_1802),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1832),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1803),
.B(n_1802),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1834),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1818),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1816),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1827),
.B(n_1874),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1897),
.B(n_1791),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1874),
.B(n_1791),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1819),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1800),
.B(n_1897),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1825),
.Y(n_1999)
);

INVxp67_ASAP7_75t_L g2000 ( 
.A(n_1780),
.Y(n_2000)
);

OAI322xp33_ASAP7_75t_L g2001 ( 
.A1(n_1767),
.A2(n_1775),
.A3(n_1763),
.B1(n_1761),
.B2(n_1843),
.C1(n_1776),
.C2(n_1858),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1795),
.B(n_1775),
.Y(n_2002)
);

OR2x2_ASAP7_75t_SL g2003 ( 
.A(n_1841),
.B(n_1799),
.Y(n_2003)
);

AO21x2_ASAP7_75t_L g2004 ( 
.A1(n_1854),
.A2(n_1900),
.B(n_1888),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1940),
.B(n_1793),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1938),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1979),
.B(n_1770),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1979),
.B(n_1788),
.Y(n_2008)
);

AOI22xp33_ASAP7_75t_L g2009 ( 
.A1(n_1980),
.A2(n_1894),
.B1(n_1847),
.B2(n_1899),
.Y(n_2009)
);

AOI222xp33_ASAP7_75t_L g2010 ( 
.A1(n_1921),
.A2(n_1908),
.B1(n_1870),
.B2(n_1905),
.C1(n_1850),
.C2(n_1849),
.Y(n_2010)
);

BUFx2_ASAP7_75t_SL g2011 ( 
.A(n_1916),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1967),
.B(n_1814),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1923),
.B(n_1864),
.Y(n_2013)
);

AOI211xp5_ASAP7_75t_L g2014 ( 
.A1(n_1981),
.A2(n_1767),
.B(n_1792),
.C(n_1904),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1937),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1967),
.B(n_1749),
.Y(n_2016)
);

AOI222xp33_ASAP7_75t_L g2017 ( 
.A1(n_1946),
.A2(n_1870),
.B1(n_1904),
.B2(n_1892),
.C1(n_1887),
.C2(n_1884),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1978),
.A2(n_1908),
.B1(n_1850),
.B2(n_1892),
.Y(n_2018)
);

OAI211xp5_ASAP7_75t_L g2019 ( 
.A1(n_1946),
.A2(n_1883),
.B(n_1873),
.C(n_1849),
.Y(n_2019)
);

NOR4xp25_ASAP7_75t_SL g2020 ( 
.A(n_1997),
.B(n_1860),
.C(n_1871),
.D(n_1809),
.Y(n_2020)
);

AOI21xp5_ASAP7_75t_L g2021 ( 
.A1(n_1935),
.A2(n_1884),
.B(n_1883),
.Y(n_2021)
);

AOI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1935),
.A2(n_1846),
.B1(n_1873),
.B2(n_1774),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1928),
.B(n_1768),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_1997),
.B(n_1846),
.C(n_1898),
.Y(n_2024)
);

OAI211xp5_ASAP7_75t_SL g2025 ( 
.A1(n_1984),
.A2(n_1975),
.B(n_1944),
.C(n_1936),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1920),
.B(n_1817),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_1971),
.B(n_1864),
.C(n_1817),
.Y(n_2027)
);

OAI211xp5_ASAP7_75t_SL g2028 ( 
.A1(n_2000),
.A2(n_1906),
.B(n_1826),
.C(n_1824),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1929),
.Y(n_2029)
);

OAI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_1971),
.A2(n_1824),
.B1(n_1826),
.B2(n_1927),
.C(n_2002),
.Y(n_2030)
);

AOI211xp5_ASAP7_75t_L g2031 ( 
.A1(n_2001),
.A2(n_1927),
.B(n_1954),
.C(n_1956),
.Y(n_2031)
);

INVx4_ASAP7_75t_R g2032 ( 
.A(n_1916),
.Y(n_2032)
);

AND2x4_ASAP7_75t_L g2033 ( 
.A(n_1942),
.B(n_1941),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1951),
.Y(n_2034)
);

BUFx2_ASAP7_75t_L g2035 ( 
.A(n_1929),
.Y(n_2035)
);

OAI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_1927),
.A2(n_2002),
.B1(n_1923),
.B2(n_1954),
.C(n_1991),
.Y(n_2036)
);

NAND4xp25_ASAP7_75t_SL g2037 ( 
.A(n_1974),
.B(n_1956),
.C(n_1970),
.D(n_1968),
.Y(n_2037)
);

NAND3xp33_ASAP7_75t_L g2038 ( 
.A(n_1970),
.B(n_1974),
.C(n_1991),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1928),
.B(n_1930),
.Y(n_2039)
);

NOR2x1_ASAP7_75t_L g2040 ( 
.A(n_1989),
.B(n_1976),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1953),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_1952),
.Y(n_2042)
);

OR2x6_ASAP7_75t_L g2043 ( 
.A(n_1942),
.B(n_1951),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1953),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1961),
.Y(n_2045)
);

AO21x2_ASAP7_75t_L g2046 ( 
.A1(n_1962),
.A2(n_1983),
.B(n_1963),
.Y(n_2046)
);

AND2x2_ASAP7_75t_L g2047 ( 
.A(n_1930),
.B(n_1968),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1957),
.B(n_1959),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1920),
.B(n_1934),
.Y(n_2049)
);

OAI321xp33_ASAP7_75t_L g2050 ( 
.A1(n_1972),
.A2(n_1992),
.A3(n_1993),
.B1(n_1966),
.B2(n_1989),
.C(n_1955),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1982),
.B(n_1999),
.Y(n_2051)
);

INVx2_ASAP7_75t_SL g2052 ( 
.A(n_1919),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2003),
.A2(n_1919),
.B1(n_1992),
.B2(n_1925),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1934),
.Y(n_2054)
);

AOI21xp33_ASAP7_75t_SL g2055 ( 
.A1(n_1986),
.A2(n_1976),
.B(n_1966),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_2001),
.A2(n_1993),
.B1(n_1988),
.B2(n_1990),
.Y(n_2056)
);

AOI22xp33_ASAP7_75t_L g2057 ( 
.A1(n_1988),
.A2(n_1990),
.B1(n_1955),
.B2(n_1995),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1957),
.B(n_1959),
.Y(n_2058)
);

BUFx3_ASAP7_75t_L g2059 ( 
.A(n_1964),
.Y(n_2059)
);

AOI22xp5_ASAP7_75t_L g2060 ( 
.A1(n_1976),
.A2(n_1996),
.B1(n_1995),
.B2(n_1960),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_1941),
.Y(n_2061)
);

NAND3xp33_ASAP7_75t_SL g2062 ( 
.A(n_1972),
.B(n_1965),
.C(n_1996),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1943),
.Y(n_2063)
);

AO31x2_ASAP7_75t_L g2064 ( 
.A1(n_1912),
.A2(n_1913),
.A3(n_1915),
.B(n_1924),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1999),
.B(n_1918),
.Y(n_2065)
);

OAI211xp5_ASAP7_75t_L g2066 ( 
.A1(n_1987),
.A2(n_1965),
.B(n_1977),
.C(n_1969),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_2003),
.A2(n_1976),
.B1(n_1922),
.B2(n_1911),
.Y(n_2067)
);

OA21x2_ASAP7_75t_L g2068 ( 
.A1(n_1962),
.A2(n_1963),
.B(n_1983),
.Y(n_2068)
);

AOI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_1995),
.A2(n_1994),
.B1(n_1998),
.B2(n_1941),
.Y(n_2069)
);

NAND3xp33_ASAP7_75t_L g2070 ( 
.A(n_1987),
.B(n_1977),
.C(n_1969),
.Y(n_2070)
);

AO21x2_ASAP7_75t_L g2071 ( 
.A1(n_1962),
.A2(n_1983),
.B(n_1963),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1949),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1918),
.B(n_1932),
.Y(n_2073)
);

BUFx2_ASAP7_75t_L g2074 ( 
.A(n_1941),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2006),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2048),
.B(n_1926),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2048),
.B(n_1926),
.Y(n_2077)
);

OR2x2_ASAP7_75t_L g2078 ( 
.A(n_2070),
.B(n_1926),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2006),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_L g2080 ( 
.A(n_2025),
.B(n_1917),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2058),
.B(n_1926),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2047),
.B(n_1931),
.Y(n_2082)
);

INVx2_ASAP7_75t_L g2083 ( 
.A(n_2068),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2047),
.B(n_1942),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2012),
.B(n_1942),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_2016),
.B(n_1948),
.Y(n_2086)
);

BUFx3_ASAP7_75t_L g2087 ( 
.A(n_2013),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2016),
.B(n_2038),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_2043),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2046),
.B(n_1913),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2046),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_2070),
.B(n_1915),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_2071),
.Y(n_2093)
);

AND2x2_ASAP7_75t_L g2094 ( 
.A(n_2071),
.B(n_2012),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_2064),
.Y(n_2095)
);

NAND2x1p5_ASAP7_75t_L g2096 ( 
.A(n_2040),
.B(n_1958),
.Y(n_2096)
);

AND2x2_ASAP7_75t_L g2097 ( 
.A(n_2039),
.B(n_1933),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2039),
.B(n_2033),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2033),
.B(n_1933),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2033),
.B(n_1933),
.Y(n_2100)
);

OR2x2_ASAP7_75t_L g2101 ( 
.A(n_2049),
.B(n_1973),
.Y(n_2101)
);

NAND4xp25_ASAP7_75t_L g2102 ( 
.A(n_2031),
.B(n_1945),
.C(n_1939),
.D(n_1985),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2049),
.B(n_1973),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2033),
.B(n_1958),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_2043),
.B(n_2064),
.Y(n_2105)
);

BUFx2_ASAP7_75t_L g2106 ( 
.A(n_2043),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2043),
.B(n_1933),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2043),
.B(n_1924),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2064),
.B(n_2004),
.Y(n_2109)
);

AND2x2_ASAP7_75t_L g2110 ( 
.A(n_2041),
.B(n_2004),
.Y(n_2110)
);

NOR2xp67_ASAP7_75t_L g2111 ( 
.A(n_2066),
.B(n_1958),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2044),
.B(n_2004),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2038),
.B(n_1950),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2063),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2008),
.B(n_1945),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2063),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2054),
.B(n_1947),
.Y(n_2117)
);

AND2x4_ASAP7_75t_L g2118 ( 
.A(n_2061),
.B(n_1958),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2072),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2015),
.B(n_1914),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2072),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_2008),
.B(n_2004),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2114),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2114),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2114),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2088),
.B(n_2042),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_2090),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2116),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2116),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2098),
.B(n_2061),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2090),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2116),
.Y(n_2132)
);

NAND3xp33_ASAP7_75t_L g2133 ( 
.A(n_2102),
.B(n_2031),
.C(n_2014),
.Y(n_2133)
);

INVx1_ASAP7_75t_SL g2134 ( 
.A(n_2113),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2102),
.A2(n_2014),
.B1(n_2022),
.B2(n_2019),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2119),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2088),
.B(n_2062),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_2111),
.A2(n_2021),
.B(n_2036),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2098),
.B(n_2074),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2098),
.B(n_2084),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_2098),
.B(n_2074),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2119),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2119),
.Y(n_2143)
);

OAI211xp5_ASAP7_75t_SL g2144 ( 
.A1(n_2078),
.A2(n_2009),
.B(n_2056),
.C(n_2022),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_2111),
.A2(n_2018),
.B(n_2024),
.Y(n_2145)
);

OAI31xp33_ASAP7_75t_L g2146 ( 
.A1(n_2078),
.A2(n_2037),
.A3(n_2067),
.B(n_2053),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_2111),
.B(n_2055),
.Y(n_2147)
);

INVxp67_ASAP7_75t_SL g2148 ( 
.A(n_2113),
.Y(n_2148)
);

AOI32xp33_ASAP7_75t_L g2149 ( 
.A1(n_2080),
.A2(n_2007),
.A3(n_2050),
.B1(n_2057),
.B2(n_2040),
.Y(n_2149)
);

OAI21xp5_ASAP7_75t_SL g2150 ( 
.A1(n_2080),
.A2(n_2010),
.B(n_2017),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2121),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2121),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_2084),
.B(n_2023),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2084),
.B(n_2023),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2086),
.B(n_2029),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2121),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2089),
.B(n_2029),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2075),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_2086),
.B(n_2059),
.Y(n_2159)
);

NOR3xp33_ASAP7_75t_L g2160 ( 
.A(n_2078),
.B(n_2024),
.C(n_2030),
.Y(n_2160)
);

AOI22xp33_ASAP7_75t_L g2161 ( 
.A1(n_2089),
.A2(n_2007),
.B1(n_2027),
.B2(n_1995),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2075),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2075),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2089),
.B(n_2035),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2079),
.Y(n_2165)
);

AND2x2_ASAP7_75t_L g2166 ( 
.A(n_2106),
.B(n_2035),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2092),
.B(n_2051),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2106),
.B(n_2052),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2106),
.B(n_2085),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_2115),
.B(n_2065),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2085),
.B(n_2082),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2115),
.B(n_2052),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2079),
.Y(n_2173)
);

OR2x2_ASAP7_75t_L g2174 ( 
.A(n_2092),
.B(n_2026),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_2087),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2115),
.B(n_2073),
.Y(n_2176)
);

AND2x2_ASAP7_75t_L g2177 ( 
.A(n_2085),
.B(n_2034),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_2096),
.Y(n_2178)
);

AND2x4_ASAP7_75t_L g2179 ( 
.A(n_2105),
.B(n_2034),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2122),
.B(n_2060),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2140),
.B(n_2122),
.Y(n_2181)
);

OAI31xp33_ASAP7_75t_L g2182 ( 
.A1(n_2133),
.A2(n_2027),
.A3(n_2081),
.B(n_2076),
.Y(n_2182)
);

NOR2xp33_ASAP7_75t_SL g2183 ( 
.A(n_2133),
.B(n_2059),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2145),
.B(n_2122),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_2140),
.B(n_2122),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2150),
.B(n_2076),
.Y(n_2186)
);

OR2x2_ASAP7_75t_L g2187 ( 
.A(n_2167),
.B(n_2092),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2123),
.Y(n_2188)
);

AND3x2_ASAP7_75t_L g2189 ( 
.A(n_2138),
.B(n_2020),
.C(n_1964),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2123),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_2171),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2124),
.Y(n_2192)
);

OR2x2_ASAP7_75t_L g2193 ( 
.A(n_2167),
.B(n_2101),
.Y(n_2193)
);

NAND2x1_ASAP7_75t_L g2194 ( 
.A(n_2178),
.B(n_2032),
.Y(n_2194)
);

NAND4xp25_ASAP7_75t_L g2195 ( 
.A(n_2135),
.B(n_2005),
.C(n_2060),
.D(n_2069),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_2160),
.B(n_2076),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2124),
.Y(n_2197)
);

NAND2xp33_ASAP7_75t_SL g2198 ( 
.A(n_2147),
.B(n_2020),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2125),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2169),
.B(n_2076),
.Y(n_2200)
);

HB1xp67_ASAP7_75t_L g2201 ( 
.A(n_2155),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2125),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2174),
.B(n_2101),
.Y(n_2203)
);

INVx1_ASAP7_75t_SL g2204 ( 
.A(n_2157),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2171),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_2128),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2135),
.A2(n_1994),
.B1(n_2077),
.B2(n_2081),
.Y(n_2207)
);

OR2x2_ASAP7_75t_L g2208 ( 
.A(n_2174),
.B(n_2101),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_2144),
.B(n_1964),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_2128),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2169),
.B(n_2077),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2149),
.B(n_2077),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_2178),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2149),
.B(n_2077),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2157),
.B(n_2081),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2129),
.Y(n_2216)
);

NAND3xp33_ASAP7_75t_L g2217 ( 
.A(n_2146),
.B(n_2055),
.C(n_2109),
.Y(n_2217)
);

INVxp67_ASAP7_75t_SL g2218 ( 
.A(n_2164),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2129),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2126),
.B(n_2081),
.Y(n_2220)
);

NOR2x1p5_ASAP7_75t_L g2221 ( 
.A(n_2137),
.B(n_2087),
.Y(n_2221)
);

AND2x4_ASAP7_75t_SL g2222 ( 
.A(n_2164),
.B(n_2105),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_2134),
.B(n_2148),
.Y(n_2223)
);

AND2x4_ASAP7_75t_L g2224 ( 
.A(n_2179),
.B(n_2105),
.Y(n_2224)
);

AO21x2_ASAP7_75t_L g2225 ( 
.A1(n_2158),
.A2(n_2093),
.B(n_2091),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_L g2226 ( 
.A(n_2159),
.B(n_2082),
.Y(n_2226)
);

AND2x2_ASAP7_75t_SL g2227 ( 
.A(n_2137),
.B(n_2109),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_2155),
.Y(n_2228)
);

OR2x2_ASAP7_75t_L g2229 ( 
.A(n_2180),
.B(n_2103),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_2166),
.B(n_2104),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2170),
.B(n_2103),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_2132),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2132),
.Y(n_2233)
);

NAND4xp75_ASAP7_75t_L g2234 ( 
.A(n_2166),
.B(n_2109),
.C(n_2107),
.D(n_2097),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_2222),
.Y(n_2235)
);

NAND4xp75_ASAP7_75t_SL g2236 ( 
.A(n_2182),
.B(n_2107),
.C(n_2168),
.D(n_2109),
.Y(n_2236)
);

OAI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2198),
.A2(n_2161),
.B1(n_2175),
.B2(n_2178),
.C(n_2096),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2188),
.Y(n_2238)
);

OR2x2_ASAP7_75t_L g2239 ( 
.A(n_2229),
.B(n_2176),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2188),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2209),
.B(n_2172),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2229),
.B(n_2136),
.Y(n_2242)
);

AOI32xp33_ASAP7_75t_L g2243 ( 
.A1(n_2183),
.A2(n_2179),
.A3(n_2168),
.B1(n_2107),
.B2(n_2097),
.Y(n_2243)
);

AOI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_2186),
.A2(n_2097),
.B1(n_2105),
.B2(n_2179),
.C(n_2107),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2199),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2217),
.A2(n_2096),
.B(n_2013),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2199),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2218),
.B(n_2175),
.Y(n_2248)
);

XNOR2xp5_ASAP7_75t_L g2249 ( 
.A(n_2195),
.B(n_1998),
.Y(n_2249)
);

INVx2_ASAP7_75t_L g2250 ( 
.A(n_2210),
.Y(n_2250)
);

INVxp67_ASAP7_75t_L g2251 ( 
.A(n_2201),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2219),
.Y(n_2252)
);

NOR2xp33_ASAP7_75t_L g2253 ( 
.A(n_2196),
.B(n_2177),
.Y(n_2253)
);

AOI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2198),
.A2(n_2028),
.B(n_2096),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2221),
.B(n_2179),
.Y(n_2255)
);

AOI22xp33_ASAP7_75t_L g2256 ( 
.A1(n_2212),
.A2(n_2087),
.B1(n_2097),
.B2(n_2104),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_SL g2257 ( 
.A(n_2227),
.B(n_2087),
.Y(n_2257)
);

INVxp67_ASAP7_75t_L g2258 ( 
.A(n_2228),
.Y(n_2258)
);

INVxp67_ASAP7_75t_SL g2259 ( 
.A(n_2223),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2219),
.Y(n_2260)
);

OAI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2214),
.A2(n_2013),
.B1(n_2177),
.B2(n_2130),
.Y(n_2261)
);

INVxp67_ASAP7_75t_L g2262 ( 
.A(n_2223),
.Y(n_2262)
);

AOI221xp5_ASAP7_75t_L g2263 ( 
.A1(n_2184),
.A2(n_2105),
.B1(n_2131),
.B2(n_2127),
.C(n_2156),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2190),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2204),
.Y(n_2265)
);

AND2x2_ASAP7_75t_L g2266 ( 
.A(n_2222),
.B(n_2130),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2210),
.Y(n_2267)
);

NAND2xp5_ASAP7_75t_L g2268 ( 
.A(n_2207),
.B(n_2227),
.Y(n_2268)
);

NOR2xp33_ASAP7_75t_L g2269 ( 
.A(n_2226),
.B(n_2153),
.Y(n_2269)
);

OAI22xp5_ASAP7_75t_L g2270 ( 
.A1(n_2234),
.A2(n_2139),
.B1(n_2141),
.B2(n_2096),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2193),
.B(n_2153),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2193),
.B(n_2154),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2192),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_2191),
.B(n_2154),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2197),
.Y(n_2275)
);

AOI222xp33_ASAP7_75t_L g2276 ( 
.A1(n_2220),
.A2(n_1964),
.B1(n_2112),
.B2(n_2110),
.C1(n_2099),
.C2(n_2100),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2202),
.Y(n_2277)
);

O2A1O1Ixp5_ASAP7_75t_R g2278 ( 
.A1(n_2268),
.A2(n_2272),
.B(n_2271),
.C(n_2274),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2259),
.B(n_2191),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2249),
.B(n_2205),
.Y(n_2280)
);

NAND2x1_ASAP7_75t_SL g2281 ( 
.A(n_2255),
.B(n_2213),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2266),
.B(n_2230),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2238),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_L g2284 ( 
.A1(n_2254),
.A2(n_2194),
.B(n_2187),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2240),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_2266),
.B(n_2230),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2245),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2265),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2251),
.B(n_2205),
.Y(n_2289)
);

OAI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2237),
.A2(n_2234),
.B1(n_2194),
.B2(n_2224),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_2248),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2247),
.Y(n_2292)
);

OR2x2_ASAP7_75t_L g2293 ( 
.A(n_2258),
.B(n_2203),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2252),
.Y(n_2294)
);

AOI22xp5_ASAP7_75t_L g2295 ( 
.A1(n_2270),
.A2(n_2189),
.B1(n_2224),
.B2(n_2099),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2260),
.Y(n_2296)
);

OAI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_2235),
.A2(n_2224),
.B1(n_2231),
.B2(n_2200),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2262),
.B(n_2203),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_2264),
.Y(n_2299)
);

OA21x2_ASAP7_75t_L g2300 ( 
.A1(n_2246),
.A2(n_2232),
.B(n_2216),
.Y(n_2300)
);

NOR4xp25_ASAP7_75t_L g2301 ( 
.A(n_2257),
.B(n_2244),
.C(n_2275),
.D(n_2273),
.Y(n_2301)
);

AOI22xp5_ASAP7_75t_L g2302 ( 
.A1(n_2253),
.A2(n_2099),
.B1(n_2100),
.B2(n_2215),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2253),
.B(n_2215),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2255),
.B(n_2200),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2235),
.B(n_2211),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2248),
.B(n_2211),
.Y(n_2306)
);

OAI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2257),
.A2(n_2231),
.B1(n_2208),
.B2(n_2187),
.Y(n_2307)
);

AOI21xp33_ASAP7_75t_L g2308 ( 
.A1(n_2241),
.A2(n_2208),
.B(n_2206),
.Y(n_2308)
);

INVx1_ASAP7_75t_SL g2309 ( 
.A(n_2291),
.Y(n_2309)
);

NOR2x1_ASAP7_75t_SL g2310 ( 
.A(n_2298),
.B(n_2277),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_L g2311 ( 
.A(n_2288),
.B(n_2269),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_2288),
.B(n_2269),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_2293),
.B(n_2239),
.Y(n_2313)
);

XNOR2x2_ASAP7_75t_L g2314 ( 
.A(n_2278),
.B(n_2263),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2282),
.B(n_2241),
.Y(n_2315)
);

INVx1_ASAP7_75t_SL g2316 ( 
.A(n_2281),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2293),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2301),
.B(n_2239),
.Y(n_2318)
);

OR2x2_ASAP7_75t_L g2319 ( 
.A(n_2298),
.B(n_2242),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_2279),
.Y(n_2320)
);

AND2x2_ASAP7_75t_L g2321 ( 
.A(n_2282),
.B(n_2286),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2286),
.B(n_2256),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2280),
.B(n_2242),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2283),
.Y(n_2324)
);

BUFx2_ASAP7_75t_L g2325 ( 
.A(n_2305),
.Y(n_2325)
);

AOI221x1_ASAP7_75t_L g2326 ( 
.A1(n_2308),
.A2(n_2261),
.B1(n_2267),
.B2(n_2250),
.C(n_2233),
.Y(n_2326)
);

NOR2xp33_ASAP7_75t_L g2327 ( 
.A(n_2289),
.B(n_2139),
.Y(n_2327)
);

NAND2xp33_ASAP7_75t_SL g2328 ( 
.A(n_2307),
.B(n_2236),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2285),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2304),
.B(n_2181),
.Y(n_2330)
);

NAND2x1_ASAP7_75t_L g2331 ( 
.A(n_2305),
.B(n_2250),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2325),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2325),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2331),
.Y(n_2334)
);

BUFx6f_ASAP7_75t_L g2335 ( 
.A(n_2331),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2310),
.Y(n_2336)
);

NAND4xp25_ASAP7_75t_L g2337 ( 
.A(n_2318),
.B(n_2295),
.C(n_2284),
.D(n_2299),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2309),
.B(n_2305),
.Y(n_2338)
);

AOI21xp33_ASAP7_75t_L g2339 ( 
.A1(n_2316),
.A2(n_2312),
.B(n_2311),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2310),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2319),
.Y(n_2341)
);

OAI22xp5_ASAP7_75t_L g2342 ( 
.A1(n_2313),
.A2(n_2303),
.B1(n_2290),
.B2(n_2306),
.Y(n_2342)
);

NOR2x1_ASAP7_75t_L g2343 ( 
.A(n_2317),
.B(n_2287),
.Y(n_2343)
);

NOR3xp33_ASAP7_75t_L g2344 ( 
.A(n_2320),
.B(n_2297),
.C(n_2292),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2319),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_SL g2346 ( 
.A(n_2313),
.B(n_2243),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2338),
.B(n_2315),
.Y(n_2347)
);

O2A1O1Ixp33_ASAP7_75t_L g2348 ( 
.A1(n_2336),
.A2(n_2329),
.B(n_2324),
.C(n_2314),
.Y(n_2348)
);

AOI21xp5_ASAP7_75t_L g2349 ( 
.A1(n_2346),
.A2(n_2328),
.B(n_2326),
.Y(n_2349)
);

AOI211xp5_ASAP7_75t_L g2350 ( 
.A1(n_2337),
.A2(n_2328),
.B(n_2314),
.C(n_2323),
.Y(n_2350)
);

AOI32xp33_ASAP7_75t_L g2351 ( 
.A1(n_2340),
.A2(n_2321),
.A3(n_2315),
.B1(n_2322),
.B2(n_2327),
.Y(n_2351)
);

AOI211xp5_ASAP7_75t_L g2352 ( 
.A1(n_2337),
.A2(n_2321),
.B(n_2322),
.C(n_2294),
.Y(n_2352)
);

NOR2xp67_ASAP7_75t_L g2353 ( 
.A(n_2334),
.B(n_2296),
.Y(n_2353)
);

NAND3xp33_ASAP7_75t_L g2354 ( 
.A(n_2343),
.B(n_2326),
.C(n_2300),
.Y(n_2354)
);

OAI211xp5_ASAP7_75t_L g2355 ( 
.A1(n_2339),
.A2(n_2300),
.B(n_2276),
.C(n_2302),
.Y(n_2355)
);

NAND4xp25_ASAP7_75t_SL g2356 ( 
.A(n_2344),
.B(n_2304),
.C(n_2330),
.D(n_2267),
.Y(n_2356)
);

OAI221xp5_ASAP7_75t_L g2357 ( 
.A1(n_2342),
.A2(n_2300),
.B1(n_2330),
.B2(n_2213),
.C(n_2011),
.Y(n_2357)
);

AOI21xp33_ASAP7_75t_SL g2358 ( 
.A1(n_2341),
.A2(n_2213),
.B(n_2232),
.Y(n_2358)
);

OAI21xp33_ASAP7_75t_SL g2359 ( 
.A1(n_2345),
.A2(n_2185),
.B(n_2181),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2332),
.A2(n_2011),
.B1(n_2185),
.B2(n_2105),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2347),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2349),
.Y(n_2362)
);

NAND2xp33_ASAP7_75t_SL g2363 ( 
.A(n_2354),
.B(n_2335),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2353),
.Y(n_2364)
);

INVx1_ASAP7_75t_SL g2365 ( 
.A(n_2356),
.Y(n_2365)
);

O2A1O1Ixp33_ASAP7_75t_L g2366 ( 
.A1(n_2348),
.A2(n_2333),
.B(n_2335),
.C(n_2131),
.Y(n_2366)
);

OAI22xp5_ASAP7_75t_L g2367 ( 
.A1(n_2350),
.A2(n_2335),
.B1(n_2127),
.B2(n_2151),
.Y(n_2367)
);

NAND2xp33_ASAP7_75t_SL g2368 ( 
.A(n_2360),
.B(n_2141),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2361),
.Y(n_2369)
);

NAND3x1_ASAP7_75t_L g2370 ( 
.A(n_2364),
.B(n_2352),
.C(n_2351),
.Y(n_2370)
);

NOR2x1_ASAP7_75t_L g2371 ( 
.A(n_2366),
.B(n_2357),
.Y(n_2371)
);

CKINVDCx5p33_ASAP7_75t_R g2372 ( 
.A(n_2362),
.Y(n_2372)
);

NOR3xp33_ASAP7_75t_SL g2373 ( 
.A(n_2363),
.B(n_2355),
.C(n_2359),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2367),
.Y(n_2374)
);

HB1xp67_ASAP7_75t_L g2375 ( 
.A(n_2365),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_2368),
.B(n_2358),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2361),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2361),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2375),
.Y(n_2379)
);

OAI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2373),
.A2(n_2142),
.B1(n_2143),
.B2(n_2151),
.Y(n_2380)
);

O2A1O1Ixp33_ASAP7_75t_L g2381 ( 
.A1(n_2375),
.A2(n_2225),
.B(n_2083),
.C(n_2095),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2371),
.A2(n_2376),
.B(n_2372),
.Y(n_2382)
);

NAND5xp2_ASAP7_75t_L g2383 ( 
.A(n_2373),
.B(n_2099),
.C(n_2100),
.D(n_2108),
.E(n_2094),
.Y(n_2383)
);

AO22x2_ASAP7_75t_L g2384 ( 
.A1(n_2374),
.A2(n_2136),
.B1(n_2142),
.B2(n_2143),
.Y(n_2384)
);

NAND4xp25_ASAP7_75t_SL g2385 ( 
.A(n_2369),
.B(n_2094),
.C(n_2108),
.D(n_2152),
.Y(n_2385)
);

NAND3xp33_ASAP7_75t_SL g2386 ( 
.A(n_2382),
.B(n_2378),
.C(n_2377),
.Y(n_2386)
);

AOI221xp5_ASAP7_75t_L g2387 ( 
.A1(n_2383),
.A2(n_2370),
.B1(n_2225),
.B2(n_2156),
.C(n_2152),
.Y(n_2387)
);

NAND4xp25_ASAP7_75t_L g2388 ( 
.A(n_2379),
.B(n_2034),
.C(n_2104),
.D(n_2108),
.Y(n_2388)
);

OAI322xp33_ASAP7_75t_L g2389 ( 
.A1(n_2380),
.A2(n_2158),
.A3(n_2173),
.B1(n_2165),
.B2(n_2163),
.C1(n_2162),
.C2(n_2083),
.Y(n_2389)
);

OAI322xp33_ASAP7_75t_L g2390 ( 
.A1(n_2387),
.A2(n_2381),
.A3(n_2384),
.B1(n_2385),
.B2(n_2162),
.C1(n_2173),
.C2(n_2165),
.Y(n_2390)
);

NAND2xp5_ASAP7_75t_L g2391 ( 
.A(n_2390),
.B(n_2386),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_2391),
.A2(n_2388),
.B1(n_2389),
.B2(n_2225),
.Y(n_2392)
);

INVx4_ASAP7_75t_L g2393 ( 
.A(n_2391),
.Y(n_2393)
);

OAI222xp33_ASAP7_75t_L g2394 ( 
.A1(n_2392),
.A2(n_2163),
.B1(n_2120),
.B2(n_2091),
.C1(n_2093),
.C2(n_2083),
.Y(n_2394)
);

OAI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_2393),
.A2(n_2120),
.B1(n_2095),
.B2(n_2091),
.Y(n_2395)
);

OAI21xp33_ASAP7_75t_L g2396 ( 
.A1(n_2395),
.A2(n_2094),
.B(n_2108),
.Y(n_2396)
);

XNOR2xp5_ASAP7_75t_L g2397 ( 
.A(n_2394),
.B(n_2104),
.Y(n_2397)
);

AOI322xp5_ASAP7_75t_L g2398 ( 
.A1(n_2396),
.A2(n_2094),
.A3(n_2095),
.B1(n_2118),
.B2(n_2093),
.C1(n_2091),
.C2(n_2083),
.Y(n_2398)
);

OAI221xp5_ASAP7_75t_L g2399 ( 
.A1(n_2398),
.A2(n_2397),
.B1(n_2120),
.B2(n_2093),
.C(n_2117),
.Y(n_2399)
);

AOI211xp5_ASAP7_75t_L g2400 ( 
.A1(n_2399),
.A2(n_2104),
.B(n_2118),
.C(n_2045),
.Y(n_2400)
);


endmodule