module fake_jpeg_15057_n_217 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_217);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_36),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_18),
.B(n_0),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_44),
.Y(n_49)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_22),
.B(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_54),
.B1(n_39),
.B2(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_50),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_17),
.B1(n_30),
.B2(n_31),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_51),
.A2(n_29),
.B1(n_35),
.B2(n_43),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_17),
.B1(n_42),
.B2(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_33),
.B(n_28),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_63),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_35),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_28),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_72),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_80),
.B1(n_56),
.B2(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_49),
.Y(n_72)
);

OA22x2_ASAP7_75t_SL g73 ( 
.A1(n_61),
.A2(n_34),
.B1(n_44),
.B2(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_78),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_16),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_59),
.B(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_83),
.B(n_62),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_49),
.B(n_62),
.C(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_98),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g89 ( 
.A(n_82),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_93),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_77),
.Y(n_107)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_34),
.Y(n_95)
);

OR2x4_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_96),
.A2(n_97),
.B1(n_70),
.B2(n_68),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_66),
.A2(n_56),
.B1(n_59),
.B2(n_60),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_50),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_101),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_46),
.Y(n_101)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_27),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_112),
.B(n_38),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_107),
.B(n_109),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_SL g108 ( 
.A1(n_95),
.A2(n_88),
.B(n_94),
.C(n_98),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_103),
.B1(n_89),
.B2(n_92),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

OA21x2_ASAP7_75t_L g111 ( 
.A1(n_95),
.A2(n_73),
.B(n_76),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_123),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_88),
.A2(n_95),
.B(n_97),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_83),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_114),
.C(n_122),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_94),
.C(n_90),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_76),
.B1(n_68),
.B2(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_124),
.B1(n_28),
.B2(n_21),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_76),
.C(n_75),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_101),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_84),
.A2(n_64),
.B1(n_81),
.B2(n_78),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_87),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_140),
.C(n_125),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

NOR4xp25_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_102),
.C(n_99),
.D(n_104),
.Y(n_129)
);

OAI322xp33_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_120),
.A3(n_116),
.B1(n_111),
.B2(n_27),
.C1(n_21),
.C2(n_23),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_117),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_115),
.B(n_99),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_134),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_82),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_106),
.B1(n_111),
.B2(n_108),
.Y(n_148)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_93),
.Y(n_139)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_38),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_142),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_47),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_144),
.Y(n_155)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_149),
.C(n_152),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_156),
.B(n_130),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_113),
.C(n_107),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_15),
.C(n_13),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_53),
.C(n_20),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_20),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_160),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_22),
.Y(n_158)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_158),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_20),
.C(n_24),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_145),
.B(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_132),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_174),
.C(n_26),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_168),
.A2(n_172),
.B1(n_26),
.B2(n_24),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_126),
.B1(n_135),
.B2(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_171),
.B1(n_173),
.B2(n_175),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_143),
.B(n_133),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_159),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_159),
.A2(n_138),
.B1(n_142),
.B2(n_128),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_147),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_22),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_153),
.B1(n_161),
.B2(n_160),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_177),
.A2(n_182),
.B1(n_184),
.B2(n_173),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_170),
.B(n_149),
.C(n_152),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_179),
.C(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_157),
.C(n_156),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_167),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_136),
.B1(n_15),
.B2(n_12),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_183),
.B(n_1),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_26),
.C(n_24),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_22),
.C(n_2),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_179),
.C(n_178),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_190),
.C(n_192),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_176),
.B1(n_4),
.B2(n_5),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_169),
.B1(n_167),
.B2(n_4),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_181),
.B(n_1),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_195),
.A2(n_22),
.B(n_7),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_3),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_196),
.A2(n_8),
.B(n_9),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_195),
.A2(n_3),
.B(n_4),
.Y(n_198)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_199),
.B(n_192),
.C(n_194),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_194),
.A2(n_3),
.B(n_7),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_201),
.A2(n_10),
.B(n_8),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_206),
.Y(n_214)
);

NAND3xp33_ASAP7_75t_SL g211 ( 
.A(n_208),
.B(n_203),
.C(n_200),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_10),
.Y(n_216)
);

AOI322xp5_ASAP7_75t_L g215 ( 
.A1(n_213),
.A2(n_210),
.A3(n_212),
.B1(n_203),
.B2(n_10),
.C1(n_8),
.C2(n_9),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_216),
.Y(n_217)
);


endmodule