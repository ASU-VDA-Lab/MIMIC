module fake_jpeg_21352_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_21),
.Y(n_26)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_18),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_38),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_11),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_37),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_37),
.B(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_44),
.A2(n_28),
.B1(n_23),
.B2(n_33),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_50),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_23),
.B1(n_21),
.B2(n_28),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_33),
.B(n_13),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_53),
.C(n_55),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_33),
.C(n_22),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

AO22x1_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_22),
.B1(n_34),
.B2(n_12),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_41),
.C(n_32),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_60),
.C(n_55),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_34),
.C(n_14),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_51),
.B(n_52),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_13),
.C(n_12),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_61),
.A2(n_40),
.B1(n_12),
.B2(n_38),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_62),
.Y(n_70)
);

BUFx24_ASAP7_75t_SL g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_3),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_6),
.C(n_8),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_71),
.B(n_8),
.Y(n_75)
);

INVxp33_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

AO21x1_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_74),
.B(n_70),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_6),
.Y(n_78)
);


endmodule