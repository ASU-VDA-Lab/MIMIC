module real_aes_7276_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_241;
wire n_168;
wire n_175;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g111 ( .A(n_0), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_1), .A2(n_160), .B(n_163), .C(n_243), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_2), .A2(n_189), .B(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g489 ( .A(n_3), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_4), .B(n_219), .Y(n_218) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_5), .A2(n_189), .B(n_473), .Y(n_472) );
AND2x6_ASAP7_75t_L g160 ( .A(n_6), .B(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g256 ( .A(n_7), .Y(n_256) );
INVx1_ASAP7_75t_L g108 ( .A(n_8), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g128 ( .A(n_8), .B(n_41), .Y(n_128) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_9), .A2(n_188), .B(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_10), .B(n_172), .Y(n_245) );
INVx1_ASAP7_75t_L g477 ( .A(n_11), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_12), .B(n_213), .Y(n_512) );
INVx1_ASAP7_75t_L g152 ( .A(n_13), .Y(n_152) );
INVx1_ASAP7_75t_L g524 ( .A(n_14), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_15), .A2(n_77), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_15), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_16), .A2(n_197), .B(n_278), .C(n_280), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_17), .B(n_219), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_18), .B(n_455), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_19), .B(n_189), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_20), .B(n_203), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_21), .A2(n_213), .B(n_264), .C(n_266), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_22), .B(n_219), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_23), .B(n_172), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_24), .A2(n_199), .B(n_280), .C(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_25), .B(n_172), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g154 ( .A(n_26), .Y(n_154) );
INVx1_ASAP7_75t_L g226 ( .A(n_27), .Y(n_226) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_28), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_29), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_30), .B(n_172), .Y(n_490) );
INVx1_ASAP7_75t_L g195 ( .A(n_31), .Y(n_195) );
INVx1_ASAP7_75t_L g467 ( .A(n_32), .Y(n_467) );
INVx2_ASAP7_75t_L g158 ( .A(n_33), .Y(n_158) );
AOI222xp33_ASAP7_75t_SL g130 ( .A1(n_34), .A2(n_131), .B1(n_134), .B2(n_727), .C1(n_728), .C2(n_730), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_35), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_36), .A2(n_213), .B(n_214), .C(n_216), .Y(n_212) );
INVxp67_ASAP7_75t_L g198 ( .A(n_37), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g211 ( .A(n_38), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_39), .A2(n_163), .B(n_225), .C(n_229), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_40), .A2(n_160), .B(n_163), .C(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_41), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g466 ( .A(n_42), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_43), .A2(n_174), .B(n_254), .C(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g533 ( .A(n_44), .B(n_172), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_45), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_46), .Y(n_191) );
INVx1_ASAP7_75t_L g262 ( .A(n_47), .Y(n_262) );
CKINVDCx16_ASAP7_75t_R g468 ( .A(n_48), .Y(n_468) );
OAI22xp5_ASAP7_75t_SL g738 ( .A1(n_49), .A2(n_59), .B1(n_739), .B2(n_740), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_49), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_50), .B(n_189), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_51), .A2(n_163), .B1(n_266), .B2(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_52), .Y(n_504) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_53), .Y(n_486) );
CKINVDCx14_ASAP7_75t_R g252 ( .A(n_54), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_55), .A2(n_216), .B(n_254), .C(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_56), .Y(n_129) );
INVx1_ASAP7_75t_L g474 ( .A(n_57), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_58), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_59), .Y(n_740) );
INVx1_ASAP7_75t_L g161 ( .A(n_60), .Y(n_161) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
INVx1_ASAP7_75t_SL g215 ( .A(n_62), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_63), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_64), .B(n_219), .Y(n_268) );
INVx1_ASAP7_75t_L g167 ( .A(n_65), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_SL g454 ( .A1(n_66), .A2(n_216), .B(n_455), .C(n_456), .Y(n_454) );
INVxp67_ASAP7_75t_L g457 ( .A(n_67), .Y(n_457) );
INVx1_ASAP7_75t_L g115 ( .A(n_68), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_69), .A2(n_189), .B(n_251), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_70), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_71), .A2(n_189), .B(n_275), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_72), .Y(n_470) );
INVx1_ASAP7_75t_L g530 ( .A(n_73), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_74), .A2(n_188), .B(n_190), .Y(n_187) );
CKINVDCx16_ASAP7_75t_R g223 ( .A(n_75), .Y(n_223) );
INVx1_ASAP7_75t_L g276 ( .A(n_76), .Y(n_276) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_77), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_78), .A2(n_160), .B(n_163), .C(n_532), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_79), .A2(n_189), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g279 ( .A(n_80), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_81), .B(n_196), .Y(n_501) );
INVx2_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
INVx1_ASAP7_75t_L g244 ( .A(n_83), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_84), .B(n_455), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_85), .A2(n_102), .B1(n_116), .B2(n_743), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_86), .A2(n_160), .B(n_163), .C(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g112 ( .A(n_87), .Y(n_112) );
OR2x2_ASAP7_75t_L g125 ( .A(n_87), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g442 ( .A(n_87), .B(n_127), .Y(n_442) );
A2O1A1Ixp33_ASAP7_75t_L g162 ( .A1(n_88), .A2(n_163), .B(n_166), .C(n_176), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_89), .B(n_181), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_90), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_91), .A2(n_160), .B(n_163), .C(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_92), .Y(n_516) );
INVx1_ASAP7_75t_L g453 ( .A(n_93), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g521 ( .A(n_94), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_95), .B(n_196), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_96), .B(n_147), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_97), .B(n_147), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_98), .B(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g265 ( .A(n_99), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_100), .A2(n_189), .B(n_452), .Y(n_451) );
BUFx4f_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx2_ASAP7_75t_L g745 ( .A(n_105), .Y(n_745) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_111), .B(n_112), .C(n_113), .Y(n_110) );
AND2x2_ASAP7_75t_L g127 ( .A(n_111), .B(n_128), .Y(n_127) );
OR2x2_ASAP7_75t_L g726 ( .A(n_112), .B(n_127), .Y(n_726) );
NOR2x2_ASAP7_75t_L g732 ( .A(n_112), .B(n_126), .Y(n_732) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_130), .B1(n_733), .B2(n_735), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_122), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g734 ( .A(n_120), .Y(n_734) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_122), .A2(n_736), .B(n_741), .Y(n_735) );
NOR2xp33_ASAP7_75t_SL g122 ( .A(n_123), .B(n_129), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g742 ( .A(n_125), .Y(n_742) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g727 ( .A(n_131), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_442), .B1(n_443), .B2(n_724), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g736 ( .A1(n_135), .A2(n_136), .B1(n_737), .B2(n_738), .Y(n_736) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_136), .A2(n_442), .B1(n_724), .B2(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_376), .Y(n_136) );
NAND5xp2_ASAP7_75t_L g137 ( .A(n_138), .B(n_305), .C(n_335), .D(n_356), .E(n_362), .Y(n_137) );
AOI221xp5_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_235), .B1(n_269), .B2(n_271), .C(n_282), .Y(n_138) );
INVxp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_232), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g141 ( .A(n_142), .B(n_204), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_SL g356 ( .A1(n_143), .A2(n_220), .B(n_357), .C(n_360), .Y(n_356) );
AND2x2_ASAP7_75t_L g426 ( .A(n_143), .B(n_221), .Y(n_426) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_182), .Y(n_143) );
AND2x2_ASAP7_75t_L g284 ( .A(n_144), .B(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g288 ( .A(n_144), .B(n_285), .Y(n_288) );
OR2x2_ASAP7_75t_L g314 ( .A(n_144), .B(n_221), .Y(n_314) );
AND2x2_ASAP7_75t_L g316 ( .A(n_144), .B(n_207), .Y(n_316) );
AND2x2_ASAP7_75t_L g334 ( .A(n_144), .B(n_206), .Y(n_334) );
INVx1_ASAP7_75t_L g367 ( .A(n_144), .Y(n_367) );
INVx2_ASAP7_75t_SL g144 ( .A(n_145), .Y(n_144) );
BUFx2_ASAP7_75t_L g234 ( .A(n_145), .Y(n_234) );
AND2x2_ASAP7_75t_L g270 ( .A(n_145), .B(n_207), .Y(n_270) );
AND2x2_ASAP7_75t_L g423 ( .A(n_145), .B(n_221), .Y(n_423) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_153), .B(n_178), .Y(n_145) );
INVx3_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_146), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_146), .B(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_SL g503 ( .A(n_146), .B(n_504), .Y(n_503) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_147), .Y(n_208) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_147), .A2(n_451), .B(n_458), .Y(n_450) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g185 ( .A(n_148), .Y(n_185) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_SL g181 ( .A(n_149), .B(n_150), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_162), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_155), .A2(n_181), .B(n_223), .C(n_224), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_155), .A2(n_241), .B(n_242), .Y(n_240) );
OAI22xp33_ASAP7_75t_L g463 ( .A1(n_155), .A2(n_177), .B1(n_464), .B2(n_468), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_155), .A2(n_486), .B(n_487), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_155), .A2(n_530), .B(n_531), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g155 ( .A(n_156), .B(n_160), .Y(n_155) );
AND2x4_ASAP7_75t_L g189 ( .A(n_156), .B(n_160), .Y(n_189) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx1_ASAP7_75t_L g200 ( .A(n_157), .Y(n_200) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g164 ( .A(n_158), .Y(n_164) );
INVx1_ASAP7_75t_L g267 ( .A(n_158), .Y(n_267) );
INVx1_ASAP7_75t_L g165 ( .A(n_159), .Y(n_165) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_159), .Y(n_170) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_159), .Y(n_172) );
INVx3_ASAP7_75t_L g197 ( .A(n_159), .Y(n_197) );
INVx1_ASAP7_75t_L g455 ( .A(n_159), .Y(n_455) );
INVx4_ASAP7_75t_SL g177 ( .A(n_160), .Y(n_177) );
BUFx3_ASAP7_75t_L g229 ( .A(n_160), .Y(n_229) );
INVx5_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
AND2x6_ASAP7_75t_L g163 ( .A(n_164), .B(n_165), .Y(n_163) );
BUFx3_ASAP7_75t_L g175 ( .A(n_164), .Y(n_175) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_164), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_168), .B(n_171), .C(n_173), .Y(n_166) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_168), .A2(n_173), .B(n_244), .C(n_245), .Y(n_243) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OAI22xp5_ASAP7_75t_SL g465 ( .A1(n_169), .A2(n_170), .B1(n_466), .B2(n_467), .Y(n_465) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx4_ASAP7_75t_L g199 ( .A(n_170), .Y(n_199) );
INVx4_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
INVx2_ASAP7_75t_L g254 ( .A(n_172), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_173), .A2(n_501), .B(n_502), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_173), .A2(n_533), .B(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g280 ( .A(n_175), .Y(n_280) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_177), .A2(n_191), .B(n_192), .C(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g210 ( .A1(n_177), .A2(n_192), .B(n_211), .C(n_212), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_SL g251 ( .A1(n_177), .A2(n_192), .B(n_252), .C(n_253), .Y(n_251) );
O2A1O1Ixp33_ASAP7_75t_SL g261 ( .A1(n_177), .A2(n_192), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_SL g275 ( .A1(n_177), .A2(n_192), .B(n_276), .C(n_277), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_L g452 ( .A1(n_177), .A2(n_192), .B(n_453), .C(n_454), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_177), .A2(n_192), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_177), .A2(n_192), .B(n_521), .C(n_522), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_180), .A2(n_508), .B(n_515), .Y(n_507) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g239 ( .A(n_181), .Y(n_239) );
OA21x2_ASAP7_75t_L g249 ( .A1(n_181), .A2(n_250), .B(n_257), .Y(n_249) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_181), .A2(n_519), .B(n_525), .Y(n_518) );
AND2x2_ASAP7_75t_L g304 ( .A(n_182), .B(n_205), .Y(n_304) );
OR2x2_ASAP7_75t_L g308 ( .A(n_182), .B(n_221), .Y(n_308) );
AND2x2_ASAP7_75t_L g333 ( .A(n_182), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g380 ( .A(n_182), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_182), .B(n_342), .Y(n_428) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_186), .B(n_201), .Y(n_182) );
INVx1_ASAP7_75t_L g286 ( .A(n_183), .Y(n_286) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_183), .A2(n_529), .B(n_535), .Y(n_528) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AOI21xp5_ASAP7_75t_SL g497 ( .A1(n_184), .A2(n_498), .B(n_499), .Y(n_497) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_185), .A2(n_463), .B(n_469), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_185), .B(n_470), .Y(n_469) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_185), .A2(n_485), .B(n_492), .Y(n_484) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_187), .A2(n_202), .B(n_286), .Y(n_285) );
BUFx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_194), .B(n_200), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_198), .B2(n_199), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_196), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_196), .A2(n_489), .B(n_490), .C(n_491), .Y(n_488) );
INVx5_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_197), .B(n_256), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_197), .B(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_197), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_199), .B(n_265), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_199), .B(n_279), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_199), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g228 ( .A(n_200), .Y(n_228) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OAI322xp33_ASAP7_75t_L g429 ( .A1(n_204), .A2(n_365), .A3(n_388), .B1(n_409), .B2(n_430), .C1(n_432), .C2(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_205), .B(n_285), .Y(n_432) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_220), .Y(n_205) );
AND2x2_ASAP7_75t_L g233 ( .A(n_206), .B(n_234), .Y(n_233) );
AND2x4_ASAP7_75t_L g301 ( .A(n_206), .B(n_221), .Y(n_301) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g342 ( .A(n_207), .B(n_221), .Y(n_342) );
AND2x2_ASAP7_75t_L g386 ( .A(n_207), .B(n_220), .Y(n_386) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_218), .Y(n_207) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_208), .A2(n_260), .B(n_268), .Y(n_259) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_208), .A2(n_274), .B(n_281), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_213), .B(n_215), .Y(n_214) );
INVx3_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_217), .Y(n_513) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_219), .A2(n_472), .B(n_478), .Y(n_471) );
AND2x2_ASAP7_75t_L g269 ( .A(n_220), .B(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g287 ( .A(n_220), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_220), .B(n_316), .Y(n_440) );
INVx3_ASAP7_75t_SL g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g232 ( .A(n_221), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_221), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g354 ( .A(n_221), .B(n_285), .Y(n_354) );
AND2x2_ASAP7_75t_L g381 ( .A(n_221), .B(n_316), .Y(n_381) );
OR2x2_ASAP7_75t_L g437 ( .A(n_221), .B(n_288), .Y(n_437) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_230), .Y(n_221) );
INVx1_ASAP7_75t_SL g323 ( .A(n_232), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_233), .B(n_354), .Y(n_355) );
AND2x2_ASAP7_75t_L g389 ( .A(n_233), .B(n_379), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_233), .B(n_312), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_233), .B(n_434), .Y(n_433) );
OAI31xp33_ASAP7_75t_L g407 ( .A1(n_235), .A2(n_269), .A3(n_408), .B(n_410), .Y(n_407) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_236), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g390 ( .A(n_236), .B(n_325), .Y(n_390) );
OR2x2_ASAP7_75t_L g397 ( .A(n_236), .B(n_398), .Y(n_397) );
OR2x2_ASAP7_75t_L g409 ( .A(n_236), .B(n_298), .Y(n_409) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g343 ( .A(n_237), .B(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g271 ( .A(n_238), .B(n_272), .Y(n_271) );
INVx4_ASAP7_75t_L g292 ( .A(n_238), .Y(n_292) );
AND2x2_ASAP7_75t_L g329 ( .A(n_238), .B(n_273), .Y(n_329) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_246), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_239), .B(n_493), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_239), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_239), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g328 ( .A(n_248), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_SL g398 ( .A(n_248), .Y(n_398) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_258), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_249), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g298 ( .A(n_249), .B(n_259), .Y(n_298) );
INVx2_ASAP7_75t_L g318 ( .A(n_249), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_249), .B(n_259), .Y(n_332) );
AND2x2_ASAP7_75t_L g339 ( .A(n_249), .B(n_295), .Y(n_339) );
BUFx3_ASAP7_75t_L g349 ( .A(n_249), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_249), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
AND2x2_ASAP7_75t_L g302 ( .A(n_258), .B(n_292), .Y(n_302) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g272 ( .A(n_259), .B(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_259), .Y(n_326) );
INVx2_ASAP7_75t_L g491 ( .A(n_266), .Y(n_491) );
INVx3_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_SL g309 ( .A(n_270), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_270), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_270), .B(n_379), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_271), .B(n_349), .Y(n_402) );
INVx1_ASAP7_75t_SL g436 ( .A(n_271), .Y(n_436) );
INVx1_ASAP7_75t_SL g344 ( .A(n_272), .Y(n_344) );
INVx1_ASAP7_75t_SL g295 ( .A(n_273), .Y(n_295) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_273), .Y(n_306) );
OR2x2_ASAP7_75t_L g317 ( .A(n_273), .B(n_292), .Y(n_317) );
AND2x2_ASAP7_75t_L g331 ( .A(n_273), .B(n_292), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_273), .B(n_321), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_287), .B(n_289), .C(n_300), .Y(n_282) );
AOI31xp33_ASAP7_75t_L g399 ( .A1(n_283), .A2(n_400), .A3(n_401), .B(n_402), .Y(n_399) );
AND2x2_ASAP7_75t_L g372 ( .A(n_284), .B(n_301), .Y(n_372) );
BUFx3_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_285), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g348 ( .A(n_285), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_285), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g303 ( .A(n_288), .Y(n_303) );
OAI222xp33_ASAP7_75t_L g412 ( .A1(n_288), .A2(n_413), .B1(n_416), .B2(n_417), .C1(n_418), .C2(n_419), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g418 ( .A(n_290), .Y(n_418) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_292), .B(n_295), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_292), .B(n_318), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_292), .B(n_293), .Y(n_388) );
INVx1_ASAP7_75t_L g439 ( .A(n_292), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g369 ( .A(n_293), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g441 ( .A(n_293), .Y(n_441) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
AOI32xp33_ASAP7_75t_L g300 ( .A1(n_296), .A2(n_301), .A3(n_302), .B1(n_303), .B2(n_304), .Y(n_300) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_298), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g375 ( .A(n_298), .Y(n_375) );
OR2x2_ASAP7_75t_L g416 ( .A(n_298), .B(n_317), .Y(n_416) );
INVx1_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_301), .B(n_312), .Y(n_337) );
INVx3_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
AOI322xp5_ASAP7_75t_L g362 ( .A1(n_301), .A2(n_346), .A3(n_363), .B1(n_365), .B2(n_368), .C1(n_372), .C2(n_373), .Y(n_362) );
AND2x2_ASAP7_75t_L g338 ( .A(n_302), .B(n_339), .Y(n_338) );
INVxp67_ASAP7_75t_L g415 ( .A(n_302), .Y(n_415) );
A2O1A1O1Ixp25_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_310), .C(n_318), .D(n_319), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_306), .B(n_349), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_308), .A2(n_320), .B1(n_323), .B2(n_324), .C(n_327), .Y(n_319) );
INVx1_ASAP7_75t_SL g434 ( .A(n_308), .Y(n_434) );
AOI21xp33_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_315), .B(n_317), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_312), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_314), .A2(n_398), .B1(n_405), .B2(n_406), .C(n_407), .Y(n_404) );
OAI222xp33_ASAP7_75t_L g435 ( .A1(n_315), .A2(n_436), .B1(n_437), .B2(n_438), .C1(n_440), .C2(n_441), .Y(n_435) );
AND2x2_ASAP7_75t_L g393 ( .A(n_316), .B(n_379), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_316), .A2(n_331), .B(n_378), .Y(n_405) );
INVx1_ASAP7_75t_L g419 ( .A(n_316), .Y(n_419) );
INVx2_ASAP7_75t_SL g322 ( .A(n_317), .Y(n_322) );
AND2x2_ASAP7_75t_L g325 ( .A(n_318), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_SL g359 ( .A(n_321), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_321), .B(n_331), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_322), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_322), .B(n_332), .Y(n_361) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI21xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_330), .B(n_333), .Y(n_327) );
INVx1_ASAP7_75t_SL g345 ( .A(n_329), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_329), .B(n_375), .Y(n_392) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
AND2x2_ASAP7_75t_L g431 ( .A(n_331), .B(n_349), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_332), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_SL g417 ( .A(n_333), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B1(n_340), .B2(n_347), .C(n_350), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_343), .B1(n_345), .B2(n_346), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI22xp33_ASAP7_75t_L g350 ( .A1(n_344), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_350) );
OR2x2_ASAP7_75t_L g421 ( .A(n_345), .B(n_349), .Y(n_421) );
OR2x2_ASAP7_75t_L g424 ( .A(n_345), .B(n_359), .Y(n_424) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g420 ( .A1(n_366), .A2(n_421), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND3xp33_ASAP7_75t_SL g376 ( .A(n_377), .B(n_391), .C(n_403), .Y(n_376) );
AOI222xp33_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B1(n_384), .B2(n_387), .C1(n_389), .C2(n_390), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_379), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g401 ( .A(n_381), .Y(n_401) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B1(n_394), .B2(n_396), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g406 ( .A(n_392), .Y(n_406) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_426), .B(n_427), .Y(n_425) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
NOR5xp2_ASAP7_75t_L g403 ( .A(n_404), .B(n_412), .C(n_420), .D(n_429), .E(n_435), .Y(n_403) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g729 ( .A(n_443), .Y(n_729) );
AND2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_661), .Y(n_443) );
NOR4xp25_ASAP7_75t_L g444 ( .A(n_445), .B(n_591), .C(n_622), .D(n_641), .Y(n_444) );
NAND4xp25_ASAP7_75t_L g445 ( .A(n_446), .B(n_549), .C(n_564), .D(n_582), .Y(n_445) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_494), .B1(n_526), .B2(n_537), .C1(n_542), .C2(n_544), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_479), .Y(n_447) );
INVx1_ASAP7_75t_L g605 ( .A(n_448), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_459), .Y(n_448) );
AND2x2_ASAP7_75t_L g480 ( .A(n_449), .B(n_471), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_449), .B(n_483), .Y(n_634) );
INVx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g541 ( .A(n_450), .B(n_461), .Y(n_541) );
AND2x2_ASAP7_75t_L g550 ( .A(n_450), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g576 ( .A(n_450), .Y(n_576) );
AND2x2_ASAP7_75t_L g597 ( .A(n_450), .B(n_461), .Y(n_597) );
BUFx2_ASAP7_75t_L g620 ( .A(n_450), .Y(n_620) );
AND2x2_ASAP7_75t_L g644 ( .A(n_450), .B(n_462), .Y(n_644) );
AND2x2_ASAP7_75t_L g708 ( .A(n_450), .B(n_471), .Y(n_708) );
AND2x2_ASAP7_75t_L g609 ( .A(n_459), .B(n_540), .Y(n_609) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_460), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_471), .Y(n_460) );
OR2x2_ASAP7_75t_L g569 ( .A(n_461), .B(n_484), .Y(n_569) );
AND2x2_ASAP7_75t_L g581 ( .A(n_461), .B(n_540), .Y(n_581) );
BUFx2_ASAP7_75t_L g713 ( .A(n_461), .Y(n_713) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g482 ( .A(n_462), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g563 ( .A(n_462), .B(n_484), .Y(n_563) );
AND2x2_ASAP7_75t_L g616 ( .A(n_462), .B(n_471), .Y(n_616) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_462), .Y(n_652) );
AND2x2_ASAP7_75t_L g539 ( .A(n_471), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_SL g551 ( .A(n_471), .Y(n_551) );
INVx2_ASAP7_75t_L g562 ( .A(n_471), .Y(n_562) );
BUFx2_ASAP7_75t_L g586 ( .A(n_471), .Y(n_586) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_471), .B(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AOI332xp33_ASAP7_75t_L g564 ( .A1(n_480), .A2(n_565), .A3(n_569), .B1(n_570), .B2(n_574), .B3(n_577), .C1(n_578), .C2(n_580), .Y(n_564) );
NAND2x1_ASAP7_75t_L g649 ( .A(n_480), .B(n_540), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_480), .B(n_554), .Y(n_700) );
A2O1A1Ixp33_ASAP7_75t_SL g582 ( .A1(n_481), .A2(n_583), .B(n_586), .C(n_587), .Y(n_582) );
AND2x2_ASAP7_75t_L g721 ( .A(n_481), .B(n_562), .Y(n_721) );
INVx3_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OR2x2_ASAP7_75t_L g618 ( .A(n_482), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g623 ( .A(n_482), .B(n_620), .Y(n_623) );
INVx1_ASAP7_75t_L g554 ( .A(n_483), .Y(n_554) );
AND2x2_ASAP7_75t_L g657 ( .A(n_483), .B(n_616), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_483), .B(n_597), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_483), .B(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_483), .B(n_575), .Y(n_683) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g540 ( .A(n_484), .Y(n_540) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_494), .A2(n_643), .A3(n_650), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_505), .Y(n_494) );
AND2x2_ASAP7_75t_L g526 ( .A(n_495), .B(n_527), .Y(n_526) );
NAND2x1_ASAP7_75t_SL g545 ( .A(n_495), .B(n_546), .Y(n_545) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_495), .Y(n_632) );
AND2x2_ASAP7_75t_L g637 ( .A(n_495), .B(n_548), .Y(n_637) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_496), .A2(n_550), .B(n_552), .C(n_555), .Y(n_549) );
OR2x2_ASAP7_75t_L g566 ( .A(n_496), .B(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g579 ( .A(n_496), .Y(n_579) );
AND2x2_ASAP7_75t_L g585 ( .A(n_496), .B(n_528), .Y(n_585) );
INVx2_ASAP7_75t_L g603 ( .A(n_496), .Y(n_603) );
AND2x2_ASAP7_75t_L g614 ( .A(n_496), .B(n_568), .Y(n_614) );
AND2x2_ASAP7_75t_L g646 ( .A(n_496), .B(n_604), .Y(n_646) );
AND2x2_ASAP7_75t_L g650 ( .A(n_496), .B(n_573), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_496), .B(n_505), .Y(n_655) );
AND2x2_ASAP7_75t_L g689 ( .A(n_496), .B(n_690), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_496), .B(n_592), .Y(n_723) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_505), .B(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g631 ( .A(n_505), .Y(n_631) );
AND2x2_ASAP7_75t_L g693 ( .A(n_505), .B(n_614), .Y(n_693) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_517), .Y(n_505) );
OR2x2_ASAP7_75t_L g547 ( .A(n_506), .B(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g557 ( .A(n_506), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_506), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g665 ( .A(n_506), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_506), .B(n_528), .Y(n_682) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x2_ASAP7_75t_L g573 ( .A(n_507), .B(n_517), .Y(n_573) );
AND2x2_ASAP7_75t_L g602 ( .A(n_507), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g613 ( .A(n_507), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_507), .B(n_568), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_514), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g527 ( .A(n_518), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g548 ( .A(n_518), .Y(n_548) );
AND2x2_ASAP7_75t_L g604 ( .A(n_518), .B(n_568), .Y(n_604) );
INVx1_ASAP7_75t_L g706 ( .A(n_526), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_527), .Y(n_710) );
INVx2_ASAP7_75t_L g568 ( .A(n_528), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_539), .B(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_539), .B(n_644), .Y(n_702) );
OR2x2_ASAP7_75t_L g543 ( .A(n_540), .B(n_541), .Y(n_543) );
INVx1_ASAP7_75t_SL g595 ( .A(n_540), .Y(n_595) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AOI221xp5_ASAP7_75t_L g598 ( .A1(n_546), .A2(n_599), .B1(n_601), .B2(n_605), .C(n_606), .Y(n_598) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g626 ( .A(n_547), .B(n_590), .Y(n_626) );
INVx2_ASAP7_75t_L g558 ( .A(n_548), .Y(n_558) );
INVx1_ASAP7_75t_L g584 ( .A(n_548), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_548), .B(n_568), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_548), .B(n_571), .Y(n_678) );
INVx1_ASAP7_75t_L g686 ( .A(n_548), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_550), .B(n_554), .Y(n_600) );
AND2x4_ASAP7_75t_L g575 ( .A(n_551), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g688 ( .A(n_554), .B(n_644), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_556), .B(n_559), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_557), .B(n_589), .Y(n_588) );
INVxp67_ASAP7_75t_L g696 ( .A(n_558), .Y(n_696) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g596 ( .A(n_562), .B(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g668 ( .A(n_562), .B(n_644), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_562), .B(n_581), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g628 ( .A1(n_563), .A2(n_597), .A3(n_604), .B1(n_629), .B2(n_632), .C1(n_633), .C2(n_635), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_563), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g694 ( .A(n_566), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g640 ( .A(n_567), .Y(n_640) );
INVx2_ASAP7_75t_L g571 ( .A(n_568), .Y(n_571) );
INVx1_ASAP7_75t_L g630 ( .A(n_568), .Y(n_630) );
CKINVDCx16_ASAP7_75t_R g577 ( .A(n_569), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x2_ASAP7_75t_L g666 ( .A(n_571), .B(n_579), .Y(n_666) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g578 ( .A(n_573), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g621 ( .A(n_573), .B(n_614), .Y(n_621) );
AND2x2_ASAP7_75t_L g625 ( .A(n_573), .B(n_585), .Y(n_625) );
OAI21xp33_ASAP7_75t_SL g635 ( .A1(n_574), .A2(n_636), .B(n_638), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g705 ( .A1(n_574), .A2(n_706), .B1(n_707), .B2(n_709), .Y(n_705) );
INVx3_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g580 ( .A(n_575), .B(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_575), .B(n_595), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_577), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g717 ( .A(n_584), .Y(n_717) );
INVx4_ASAP7_75t_L g590 ( .A(n_585), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_585), .B(n_612), .Y(n_660) );
INVx1_ASAP7_75t_SL g672 ( .A(n_586), .Y(n_672) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp67_ASAP7_75t_L g685 ( .A(n_590), .B(n_686), .Y(n_685) );
OAI211xp5_ASAP7_75t_SL g591 ( .A1(n_592), .A2(n_593), .B(n_598), .C(n_615), .Y(n_591) );
OAI221xp5_ASAP7_75t_SL g711 ( .A1(n_593), .A2(n_631), .B1(n_710), .B2(n_712), .C(n_714), .Y(n_711) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_595), .B(n_708), .Y(n_707) );
OAI31xp33_ASAP7_75t_L g687 ( .A1(n_596), .A2(n_673), .A3(n_688), .B(n_689), .Y(n_687) );
INVx1_ASAP7_75t_L g627 ( .A(n_597), .Y(n_627) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g677 ( .A(n_602), .Y(n_677) );
AND2x2_ASAP7_75t_L g690 ( .A(n_604), .B(n_613), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_610), .Y(n_606) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_614), .B(n_717), .Y(n_716) );
OAI21xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B(n_621), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_624), .B1(n_626), .B2(n_627), .C(n_628), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g691 ( .A1(n_623), .A2(n_692), .B(n_694), .C(n_697), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_626), .B(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx1_ASAP7_75t_L g653 ( .A(n_634), .Y(n_653) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g639 ( .A(n_637), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g681 ( .A(n_637), .B(n_682), .Y(n_681) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_645), .B(n_647), .C(n_656), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
OAI221xp5_ASAP7_75t_L g718 ( .A1(n_645), .A2(n_655), .B1(n_719), .B2(n_720), .C(n_722), .Y(n_718) );
INVx1_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B1(n_651), .B2(n_654), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OAI21xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_658), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_SL g719 ( .A(n_658), .Y(n_719) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NOR4xp25_ASAP7_75t_L g661 ( .A(n_662), .B(n_691), .C(n_711), .D(n_718), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_667), .B(n_669), .C(n_687), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_666), .Y(n_663) );
INVxp67_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_673), .B(n_675), .C(n_679), .Y(n_669) );
INVx1_ASAP7_75t_SL g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_SL g698 ( .A(n_676), .Y(n_698) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
OR2x2_ASAP7_75t_L g709 ( .A(n_677), .B(n_710), .Y(n_709) );
OAI21xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_683), .B(n_684), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B1(n_701), .B2(n_703), .C(n_705), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_708), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g733 ( .A(n_734), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
endmodule