module real_aes_1170_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_776, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_776;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g154 ( .A(n_0), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_1), .B(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_2), .B(n_160), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_3), .B(n_157), .Y(n_504) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_4), .A2(n_99), .B1(n_739), .B2(n_750), .C1(n_762), .C2(n_766), .Y(n_98) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_4), .A2(n_102), .B1(n_103), .B2(n_753), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_4), .Y(n_753) );
INVx1_ASAP7_75t_L g120 ( .A(n_5), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_6), .B(n_160), .Y(n_182) );
NAND2xp33_ASAP7_75t_SL g140 ( .A(n_7), .B(n_141), .Y(n_140) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g746 ( .A(n_9), .Y(n_746) );
AND2x2_ASAP7_75t_L g180 ( .A(n_10), .B(n_163), .Y(n_180) );
AND2x2_ASAP7_75t_L g455 ( .A(n_11), .B(n_136), .Y(n_455) );
AND2x2_ASAP7_75t_L g506 ( .A(n_12), .B(n_191), .Y(n_506) );
INVx2_ASAP7_75t_L g114 ( .A(n_13), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_14), .B(n_157), .Y(n_479) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_15), .Y(n_428) );
AOI221x1_ASAP7_75t_L g132 ( .A1(n_16), .A2(n_133), .B1(n_135), .B2(n_136), .C(n_139), .Y(n_132) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_17), .B(n_160), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_18), .B(n_160), .Y(n_511) );
INVx1_ASAP7_75t_L g431 ( .A(n_19), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_20), .A2(n_87), .B1(n_115), .B2(n_160), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_21), .A2(n_135), .B(n_184), .Y(n_183) );
AOI221xp5_ASAP7_75t_SL g227 ( .A1(n_22), .A2(n_35), .B1(n_135), .B2(n_160), .C(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_23), .B(n_155), .Y(n_185) );
OR2x2_ASAP7_75t_L g113 ( .A(n_24), .B(n_86), .Y(n_113) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_24), .A2(n_86), .B(n_114), .Y(n_138) );
INVxp67_ASAP7_75t_L g131 ( .A(n_25), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_26), .B(n_157), .Y(n_222) );
AND2x2_ASAP7_75t_L g174 ( .A(n_27), .B(n_162), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_28), .A2(n_135), .B(n_153), .Y(n_152) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_29), .A2(n_136), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_30), .B(n_157), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_31), .A2(n_135), .B(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_32), .B(n_157), .Y(n_487) );
AND2x2_ASAP7_75t_L g122 ( .A(n_33), .B(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g126 ( .A(n_33), .Y(n_126) );
AND2x2_ASAP7_75t_L g141 ( .A(n_33), .B(n_120), .Y(n_141) );
OR2x6_ASAP7_75t_L g429 ( .A(n_34), .B(n_430), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_36), .B(n_160), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_37), .A2(n_78), .B1(n_124), .B2(n_135), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_38), .B(n_157), .Y(n_470) );
INVx1_ASAP7_75t_L g732 ( .A(n_39), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_40), .B(n_160), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_41), .B(n_155), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_42), .A2(n_135), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g161 ( .A(n_43), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_44), .B(n_155), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_45), .B(n_162), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_46), .B(n_160), .Y(n_476) );
INVx1_ASAP7_75t_L g118 ( .A(n_47), .Y(n_118) );
INVx1_ASAP7_75t_L g145 ( .A(n_47), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_48), .B(n_157), .Y(n_453) );
AND2x2_ASAP7_75t_L g465 ( .A(n_49), .B(n_162), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_50), .B(n_160), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_51), .B(n_155), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_52), .B(n_155), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_53), .A2(n_732), .B1(n_734), .B2(n_737), .Y(n_733) );
AND2x2_ASAP7_75t_L g203 ( .A(n_54), .B(n_162), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g454 ( .A(n_55), .B(n_160), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_56), .B(n_157), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_57), .B(n_160), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_58), .A2(n_135), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_59), .B(n_155), .Y(n_201) );
AND2x2_ASAP7_75t_SL g223 ( .A(n_60), .B(n_163), .Y(n_223) );
AND2x2_ASAP7_75t_L g517 ( .A(n_61), .B(n_163), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_62), .A2(n_135), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_63), .B(n_157), .Y(n_186) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_64), .B(n_191), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_65), .B(n_155), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_66), .B(n_155), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_67), .A2(n_89), .B1(n_124), .B2(n_135), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_68), .B(n_157), .Y(n_514) );
INVx1_ASAP7_75t_L g123 ( .A(n_69), .Y(n_123) );
INVx1_ASAP7_75t_L g147 ( .A(n_69), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_70), .B(n_155), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_71), .A2(n_135), .B(n_469), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_72), .A2(n_135), .B(n_443), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_73), .A2(n_135), .B(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g489 ( .A(n_74), .B(n_163), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_75), .B(n_162), .Y(n_457) );
AOI22xp5_ASAP7_75t_L g193 ( .A1(n_76), .A2(n_81), .B1(n_115), .B2(n_160), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_77), .B(n_160), .Y(n_202) );
INVx1_ASAP7_75t_L g432 ( .A(n_79), .Y(n_432) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_80), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_82), .B(n_155), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_83), .B(n_155), .Y(n_230) );
AND2x2_ASAP7_75t_L g446 ( .A(n_84), .B(n_191), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_85), .A2(n_135), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_88), .B(n_157), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_90), .A2(n_135), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_91), .B(n_157), .Y(n_444) );
INVxp67_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_93), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_94), .B(n_157), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_95), .A2(n_135), .B(n_220), .Y(n_219) );
BUFx2_ASAP7_75t_L g516 ( .A(n_96), .Y(n_516) );
BUFx2_ASAP7_75t_L g747 ( .A(n_97), .Y(n_747) );
BUFx2_ASAP7_75t_SL g772 ( .A(n_97), .Y(n_772) );
OAI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_732), .B(n_733), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_426), .B1(n_433), .B2(n_728), .Y(n_101) );
INVx3_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OA22x2_ASAP7_75t_L g735 ( .A1(n_103), .A2(n_426), .B1(n_434), .B2(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_303), .Y(n_103) );
NOR4xp25_ASAP7_75t_L g104 ( .A(n_105), .B(n_246), .C(n_285), .D(n_292), .Y(n_104) );
OAI221xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_164), .B1(n_204), .B2(n_213), .C(n_232), .Y(n_105) );
OR2x2_ASAP7_75t_L g376 ( .A(n_106), .B(n_238), .Y(n_376) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g291 ( .A(n_107), .B(n_216), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_107), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_107), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g107 ( .A(n_108), .B(n_148), .Y(n_107) );
AND2x4_ASAP7_75t_SL g215 ( .A(n_108), .B(n_216), .Y(n_215) );
INVx3_ASAP7_75t_L g237 ( .A(n_108), .Y(n_237) );
AND2x2_ASAP7_75t_L g272 ( .A(n_108), .B(n_245), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_108), .B(n_149), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_108), .B(n_239), .Y(n_324) );
OR2x2_ASAP7_75t_L g402 ( .A(n_108), .B(n_216), .Y(n_402) );
AND2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_132), .Y(n_108) );
AOI22xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_115), .B1(n_124), .B2(n_130), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g130 ( .A(n_112), .B(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_112), .B(n_134), .Y(n_133) );
NOR3xp33_ASAP7_75t_L g139 ( .A(n_112), .B(n_140), .C(n_142), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_112), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_112), .A2(n_467), .B(n_468), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_112), .A2(n_476), .B(n_477), .Y(n_475) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AND2x2_ASAP7_75t_SL g163 ( .A(n_113), .B(n_114), .Y(n_163) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_121), .Y(n_115) );
AND2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_119), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g129 ( .A(n_118), .B(n_120), .Y(n_129) );
AND2x4_ASAP7_75t_L g157 ( .A(n_118), .B(n_146), .Y(n_157) );
HB1xp67_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AND2x6_ASAP7_75t_L g135 ( .A(n_122), .B(n_129), .Y(n_135) );
INVx2_ASAP7_75t_L g128 ( .A(n_123), .Y(n_128) );
AND2x6_ASAP7_75t_L g155 ( .A(n_123), .B(n_144), .Y(n_155) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
NOR2x1p5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx3_ASAP7_75t_L g482 ( .A(n_136), .Y(n_482) );
INVx4_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21x1_ASAP7_75t_L g150 ( .A1(n_137), .A2(n_151), .B(n_161), .Y(n_150) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_137), .A2(n_449), .B(n_455), .Y(n_448) );
INVx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx4f_ASAP7_75t_L g191 ( .A(n_138), .Y(n_191) );
INVx5_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
AND2x4_ASAP7_75t_L g160 ( .A(n_141), .B(n_143), .Y(n_160) );
INVx1_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AND2x2_ASAP7_75t_L g224 ( .A(n_149), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_149), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g250 ( .A(n_149), .Y(n_250) );
OR2x2_ASAP7_75t_L g255 ( .A(n_149), .B(n_239), .Y(n_255) );
AND2x2_ASAP7_75t_L g268 ( .A(n_149), .B(n_226), .Y(n_268) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_149), .Y(n_271) );
INVx1_ASAP7_75t_L g283 ( .A(n_149), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_149), .B(n_237), .Y(n_348) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_159), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_156), .B(n_158), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_155), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_158), .A2(n_170), .B(n_171), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_158), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_221), .B(n_222), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_158), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_158), .A2(n_444), .B(n_445), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_158), .A2(n_452), .B(n_453), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_158), .A2(n_470), .B(n_471), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_158), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_158), .A2(n_486), .B(n_487), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_158), .A2(n_503), .B(n_504), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_158), .A2(n_514), .B(n_515), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_162), .Y(n_173) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_162), .A2(n_227), .B(n_231), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_162), .A2(n_441), .B(n_442), .Y(n_440) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_162), .A2(n_459), .B(n_460), .Y(n_458) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_165), .B(n_175), .Y(n_164) );
HB1xp67_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OR2x2_ASAP7_75t_L g212 ( .A(n_166), .B(n_196), .Y(n_212) );
AND2x4_ASAP7_75t_L g242 ( .A(n_166), .B(n_179), .Y(n_242) );
INVx2_ASAP7_75t_L g276 ( .A(n_166), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_166), .B(n_196), .Y(n_334) );
AND2x2_ASAP7_75t_L g381 ( .A(n_166), .B(n_210), .Y(n_381) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_173), .B(n_174), .Y(n_166) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_167), .A2(n_173), .B(n_174), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_168), .B(n_172), .Y(n_167) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_173), .A2(n_197), .B(n_203), .Y(n_196) );
AOI21x1_ASAP7_75t_L g499 ( .A1(n_173), .A2(n_500), .B(n_506), .Y(n_499) );
AOI222xp33_ASAP7_75t_L g369 ( .A1(n_175), .A2(n_241), .B1(n_284), .B2(n_344), .C1(n_370), .C2(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_177), .B(n_187), .Y(n_176) );
AND2x2_ASAP7_75t_L g288 ( .A(n_177), .B(n_208), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_177), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g417 ( .A(n_177), .B(n_257), .Y(n_417) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_178), .A2(n_248), .B(n_252), .Y(n_247) );
AND2x2_ASAP7_75t_L g328 ( .A(n_178), .B(n_211), .Y(n_328) );
OR2x2_ASAP7_75t_L g353 ( .A(n_178), .B(n_212), .Y(n_353) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx5_ASAP7_75t_L g207 ( .A(n_179), .Y(n_207) );
AND2x2_ASAP7_75t_L g294 ( .A(n_179), .B(n_276), .Y(n_294) );
AND2x2_ASAP7_75t_L g320 ( .A(n_179), .B(n_196), .Y(n_320) );
OR2x2_ASAP7_75t_L g323 ( .A(n_179), .B(n_210), .Y(n_323) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_179), .Y(n_341) );
AND2x4_ASAP7_75t_SL g398 ( .A(n_179), .B(n_275), .Y(n_398) );
OR2x2_ASAP7_75t_L g407 ( .A(n_179), .B(n_234), .Y(n_407) );
OR2x6_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
INVx1_ASAP7_75t_L g240 ( .A(n_187), .Y(n_240) );
AOI221xp5_ASAP7_75t_SL g358 ( .A1(n_187), .A2(n_242), .B1(n_359), .B2(n_361), .C(n_362), .Y(n_358) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_196), .Y(n_187) );
OR2x2_ASAP7_75t_L g297 ( .A(n_188), .B(n_267), .Y(n_297) );
OR2x2_ASAP7_75t_L g307 ( .A(n_188), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g333 ( .A(n_188), .B(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g339 ( .A(n_188), .B(n_258), .Y(n_339) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_188), .B(n_322), .Y(n_351) );
INVx2_ASAP7_75t_L g364 ( .A(n_188), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_188), .B(n_242), .Y(n_385) );
AND2x2_ASAP7_75t_L g389 ( .A(n_188), .B(n_211), .Y(n_389) );
AND2x2_ASAP7_75t_L g397 ( .A(n_188), .B(n_398), .Y(n_397) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
AOI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B(n_195), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_191), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_191), .A2(n_511), .B(n_512), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_196), .B(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g241 ( .A(n_196), .B(n_210), .Y(n_241) );
INVx2_ASAP7_75t_L g258 ( .A(n_196), .Y(n_258) );
AND2x4_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_196), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g387 ( .A(n_206), .B(n_209), .Y(n_387) );
AND2x4_ASAP7_75t_L g233 ( .A(n_207), .B(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g274 ( .A(n_207), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g301 ( .A(n_207), .B(n_241), .Y(n_301) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_211), .Y(n_208) );
AND2x2_ASAP7_75t_L g405 ( .A(n_209), .B(n_406), .Y(n_405) );
BUFx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g257 ( .A(n_210), .B(n_258), .Y(n_257) );
OAI21xp5_ASAP7_75t_SL g277 ( .A1(n_211), .A2(n_278), .B(n_284), .Y(n_277) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_SL g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_224), .Y(n_214) );
INVx1_ASAP7_75t_SL g331 ( .A(n_215), .Y(n_331) );
AND2x2_ASAP7_75t_L g361 ( .A(n_215), .B(n_271), .Y(n_361) );
AND2x4_ASAP7_75t_L g372 ( .A(n_215), .B(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g238 ( .A(n_216), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g245 ( .A(n_216), .Y(n_245) );
AND2x4_ASAP7_75t_L g251 ( .A(n_216), .B(n_237), .Y(n_251) );
INVx2_ASAP7_75t_L g262 ( .A(n_216), .Y(n_262) );
INVx1_ASAP7_75t_L g311 ( .A(n_216), .Y(n_311) );
OR2x2_ASAP7_75t_L g332 ( .A(n_216), .B(n_316), .Y(n_332) );
OR2x2_ASAP7_75t_L g346 ( .A(n_216), .B(n_226), .Y(n_346) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_216), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_216), .B(n_268), .Y(n_418) );
OR2x6_ASAP7_75t_L g216 ( .A(n_217), .B(n_223), .Y(n_216) );
INVx1_ASAP7_75t_L g263 ( .A(n_224), .Y(n_263) );
AND2x2_ASAP7_75t_L g396 ( .A(n_224), .B(n_262), .Y(n_396) );
AND2x2_ASAP7_75t_L g421 ( .A(n_224), .B(n_251), .Y(n_421) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g239 ( .A(n_226), .Y(n_239) );
BUFx3_ASAP7_75t_L g281 ( .A(n_226), .Y(n_281) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_226), .Y(n_308) );
INVx1_ASAP7_75t_L g317 ( .A(n_226), .Y(n_317) );
AOI33xp33_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_235), .A3(n_240), .B1(n_241), .B2(n_242), .B3(n_243), .Y(n_232) );
AOI21x1_ASAP7_75t_SL g335 ( .A1(n_233), .A2(n_257), .B(n_319), .Y(n_335) );
INVx2_ASAP7_75t_L g365 ( .A(n_233), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_233), .B(n_364), .Y(n_371) );
AND2x2_ASAP7_75t_L g319 ( .A(n_234), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g282 ( .A(n_237), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g383 ( .A(n_238), .Y(n_383) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_239), .Y(n_373) );
OAI32xp33_ASAP7_75t_L g422 ( .A1(n_240), .A2(n_242), .A3(n_418), .B1(n_423), .B2(n_425), .Y(n_422) );
AND2x2_ASAP7_75t_L g340 ( .A(n_241), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g330 ( .A(n_242), .Y(n_330) );
AND2x2_ASAP7_75t_L g395 ( .A(n_242), .B(n_339), .Y(n_395) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
OAI221xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_256), .B1(n_259), .B2(n_273), .C(n_277), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_250), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_251), .B(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_251), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_251), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g300 ( .A(n_255), .Y(n_300) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NOR3xp33_ASAP7_75t_L g259 ( .A(n_260), .B(n_264), .C(n_269), .Y(n_259) );
INVx1_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g362 ( .A1(n_261), .A2(n_323), .B1(n_363), .B2(n_366), .Y(n_362) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx1_ASAP7_75t_L g266 ( .A(n_262), .Y(n_266) );
NOR2x1p5_ASAP7_75t_L g280 ( .A(n_262), .B(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_262), .Y(n_302) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OAI322xp33_ASAP7_75t_L g329 ( .A1(n_265), .A2(n_307), .A3(n_330), .B1(n_331), .B2(n_332), .C1(n_333), .C2(n_335), .Y(n_329) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
A2O1A1Ixp33_ASAP7_75t_L g285 ( .A1(n_267), .A2(n_286), .B(n_287), .C(n_289), .Y(n_285) );
OR2x2_ASAP7_75t_L g377 ( .A(n_267), .B(n_331), .Y(n_377) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g284 ( .A(n_268), .B(n_272), .Y(n_284) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g290 ( .A(n_274), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_SL g322 ( .A(n_275), .Y(n_322) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_279), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx1_ASAP7_75t_SL g326 ( .A(n_282), .Y(n_326) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_283), .Y(n_368) );
OR2x6_ASAP7_75t_SL g423 ( .A(n_286), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_291), .A2(n_414), .B(n_415), .C(n_422), .Y(n_413) );
O2A1O1Ixp33_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_298), .C(n_302), .Y(n_292) );
OAI211xp5_ASAP7_75t_SL g304 ( .A1(n_293), .A2(n_305), .B(n_312), .C(n_336), .Y(n_304) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_349), .C(n_393), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_306), .B(n_309), .Y(n_305) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_308), .Y(n_400) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g355 ( .A(n_311), .Y(n_355) );
NOR3xp33_ASAP7_75t_SL g312 ( .A(n_313), .B(n_325), .C(n_329), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B1(n_321), .B2(n_324), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g357 ( .A(n_317), .Y(n_357) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_317), .Y(n_424) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_SL g410 ( .A(n_323), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OR2x2_ASAP7_75t_L g360 ( .A(n_326), .B(n_346), .Y(n_360) );
OR2x2_ASAP7_75t_L g411 ( .A(n_326), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g409 ( .A(n_334), .Y(n_409) );
OR2x2_ASAP7_75t_L g425 ( .A(n_334), .B(n_364), .Y(n_425) );
OAI21xp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_340), .B(n_342), .Y(n_336) );
OAI31xp33_ASAP7_75t_L g350 ( .A1(n_337), .A2(n_351), .A3(n_352), .B(n_354), .Y(n_350) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_347), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g382 ( .A(n_347), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND4xp25_ASAP7_75t_SL g349 ( .A(n_350), .B(n_358), .C(n_369), .D(n_374), .Y(n_349) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_357), .Y(n_392) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_382), .B2(n_384), .C(n_386), .Y(n_374) );
NAND2xp33_ASAP7_75t_SL g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g419 ( .A(n_378), .Y(n_419) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI21xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_388), .B(n_390), .Y(n_386) );
INVx1_ASAP7_75t_L g414 ( .A(n_388), .Y(n_414) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_394), .B(n_413), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B1(n_397), .B2(n_399), .C(n_403), .Y(n_394) );
AND2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_408), .B(n_411), .Y(n_403) );
INVxp33_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
CKINVDCx11_ASAP7_75t_R g426 ( .A(n_427), .Y(n_426) );
AND2x6_ASAP7_75t_SL g427 ( .A(n_428), .B(n_429), .Y(n_427) );
OR2x6_ASAP7_75t_SL g730 ( .A(n_428), .B(n_731), .Y(n_730) );
OR2x2_ASAP7_75t_L g738 ( .A(n_428), .B(n_429), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_428), .B(n_731), .Y(n_749) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_429), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_431), .B(n_432), .Y(n_430) );
INVx3_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_SL g434 ( .A(n_435), .B(n_624), .Y(n_434) );
NOR3xp33_ASAP7_75t_SL g435 ( .A(n_436), .B(n_533), .C(n_565), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_461), .B1(n_490), .B2(n_507), .C(n_518), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_447), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g496 ( .A(n_439), .B(n_448), .Y(n_496) );
INVx4_ASAP7_75t_L g524 ( .A(n_439), .Y(n_524) );
AND2x4_ASAP7_75t_SL g564 ( .A(n_439), .B(n_498), .Y(n_564) );
BUFx2_ASAP7_75t_L g574 ( .A(n_439), .Y(n_574) );
NOR2x1_ASAP7_75t_L g640 ( .A(n_439), .B(n_579), .Y(n_640) );
AND2x2_ASAP7_75t_L g649 ( .A(n_439), .B(n_577), .Y(n_649) );
OR2x2_ASAP7_75t_L g657 ( .A(n_439), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g683 ( .A(n_439), .B(n_522), .Y(n_683) );
AND2x4_ASAP7_75t_L g702 ( .A(n_439), .B(n_703), .Y(n_702) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_446), .Y(n_439) );
INVx2_ASAP7_75t_SL g615 ( .A(n_447), .Y(n_615) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_456), .Y(n_447) );
AND2x2_ASAP7_75t_L g522 ( .A(n_448), .B(n_499), .Y(n_522) );
INVx2_ASAP7_75t_L g549 ( .A(n_448), .Y(n_549) );
INVx2_ASAP7_75t_L g579 ( .A(n_448), .Y(n_579) );
AND2x2_ASAP7_75t_L g593 ( .A(n_448), .B(n_498), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_454), .Y(n_449) );
AND2x2_ASAP7_75t_L g523 ( .A(n_456), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g546 ( .A(n_456), .Y(n_546) );
BUFx3_ASAP7_75t_L g560 ( .A(n_456), .Y(n_560) );
AND2x2_ASAP7_75t_L g589 ( .A(n_456), .B(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AND2x4_ASAP7_75t_L g494 ( .A(n_457), .B(n_458), .Y(n_494) );
INVx1_ASAP7_75t_L g595 ( .A(n_461), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_472), .Y(n_461) );
OR2x2_ASAP7_75t_L g706 ( .A(n_462), .B(n_507), .Y(n_706) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g562 ( .A(n_463), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_463), .B(n_472), .Y(n_623) );
OR2x2_ASAP7_75t_L g721 ( .A(n_463), .B(n_643), .Y(n_721) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g532 ( .A(n_464), .B(n_508), .Y(n_532) );
OR2x2_ASAP7_75t_SL g542 ( .A(n_464), .B(n_543), .Y(n_542) );
INVx4_ASAP7_75t_L g553 ( .A(n_464), .Y(n_553) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_464), .Y(n_604) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_464), .B(n_509), .Y(n_610) );
AND2x2_ASAP7_75t_L g635 ( .A(n_464), .B(n_474), .Y(n_635) );
OR2x2_ASAP7_75t_L g656 ( .A(n_464), .B(n_539), .Y(n_656) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g551 ( .A(n_472), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_472), .A2(n_645), .B(n_648), .C(n_650), .Y(n_644) );
AND2x2_ASAP7_75t_L g717 ( .A(n_472), .B(n_493), .Y(n_717) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
INVx1_ASAP7_75t_L g584 ( .A(n_473), .Y(n_584) );
AND2x2_ASAP7_75t_L g654 ( .A(n_473), .B(n_509), .Y(n_654) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
OR2x2_ASAP7_75t_L g543 ( .A(n_474), .B(n_509), .Y(n_543) );
INVx1_ASAP7_75t_L g559 ( .A(n_474), .Y(n_559) );
AND2x2_ASAP7_75t_L g571 ( .A(n_474), .B(n_481), .Y(n_571) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_474), .Y(n_677) );
NOR2x1_ASAP7_75t_SL g508 ( .A(n_481), .B(n_509), .Y(n_508) );
AO21x1_ASAP7_75t_SL g481 ( .A1(n_482), .A2(n_483), .B(n_489), .Y(n_481) );
AO21x2_ASAP7_75t_L g540 ( .A1(n_482), .A2(n_483), .B(n_489), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_488), .Y(n_483) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_495), .Y(n_491) );
OR2x2_ASAP7_75t_L g641 ( .A(n_492), .B(n_576), .Y(n_641) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_493), .B(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g723 ( .A(n_493), .B(n_620), .Y(n_723) );
INVx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g568 ( .A(n_494), .B(n_549), .Y(n_568) );
AND2x2_ASAP7_75t_L g664 ( .A(n_494), .B(n_577), .Y(n_664) );
INVx1_ASAP7_75t_L g581 ( .A(n_495), .Y(n_581) );
AND2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
INVx1_ASAP7_75t_L g631 ( .A(n_496), .Y(n_631) );
INVx2_ASAP7_75t_L g598 ( .A(n_497), .Y(n_598) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g548 ( .A(n_498), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g578 ( .A(n_498), .Y(n_578) );
INVx1_ASAP7_75t_L g703 ( .A(n_498), .Y(n_703) );
INVx3_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_499), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
OR2x2_ASAP7_75t_L g674 ( .A(n_507), .B(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_SL g529 ( .A(n_509), .Y(n_529) );
OR2x2_ASAP7_75t_L g552 ( .A(n_509), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g563 ( .A(n_509), .B(n_539), .Y(n_563) );
AND2x2_ASAP7_75t_L g637 ( .A(n_509), .B(n_553), .Y(n_637) );
BUFx2_ASAP7_75t_L g720 ( .A(n_509), .Y(n_720) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_517), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_525), .B(n_530), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
AND2x2_ASAP7_75t_L g672 ( .A(n_521), .B(n_594), .Y(n_672) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g531 ( .A(n_522), .B(n_524), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_523), .B(n_593), .Y(n_694) );
INVx1_ASAP7_75t_L g724 ( .A(n_523), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g620 ( .A(n_524), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_524), .B(n_660), .Y(n_697) );
INVxp67_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_529), .Y(n_526) );
AND2x4_ASAP7_75t_SL g561 ( .A(n_527), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_527), .B(n_555), .Y(n_708) );
INVx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_528), .B(n_610), .Y(n_666) );
AND2x2_ASAP7_75t_L g684 ( .A(n_528), .B(n_637), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_529), .B(n_571), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_529), .A2(n_575), .B(n_617), .C(n_622), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_529), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_531), .A2(n_604), .B1(n_712), .B2(n_718), .C(n_722), .Y(n_711) );
INVx1_ASAP7_75t_SL g699 ( .A(n_532), .Y(n_699) );
OAI221xp5_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_544), .B1(n_550), .B2(n_554), .C(n_776), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g609 ( .A(n_538), .Y(n_609) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g583 ( .A(n_539), .B(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g614 ( .A(n_539), .B(n_559), .Y(n_614) );
INVx2_ASAP7_75t_L g647 ( .A(n_539), .Y(n_647) );
INVx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI32xp33_ASAP7_75t_L g698 ( .A1(n_542), .A2(n_589), .A3(n_620), .B1(n_699), .B2(n_700), .Y(n_698) );
OR2x2_ASAP7_75t_L g669 ( .A(n_543), .B(n_656), .Y(n_669) );
INVx1_ASAP7_75t_L g679 ( .A(n_544), .Y(n_679) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_547), .Y(n_544) );
INVx2_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
AND2x2_ASAP7_75t_L g665 ( .A(n_545), .B(n_640), .Y(n_665) );
OR2x2_ASAP7_75t_L g696 ( .A(n_545), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_546), .B(n_601), .Y(n_600) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx1_ASAP7_75t_L g590 ( .A(n_549), .Y(n_590) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx2_ASAP7_75t_SL g555 ( .A(n_552), .Y(n_555) );
OR2x2_ASAP7_75t_L g642 ( .A(n_552), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_553), .B(n_571), .Y(n_570) );
NOR2xp67_ASAP7_75t_L g676 ( .A(n_553), .B(n_677), .Y(n_676) );
BUFx2_ASAP7_75t_L g689 ( .A(n_553), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_556), .B(n_561), .C(n_564), .Y(n_554) );
AND2x2_ASAP7_75t_L g704 ( .A(n_556), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_560), .Y(n_557) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g630 ( .A(n_560), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_560), .B(n_564), .Y(n_651) );
AND2x2_ASAP7_75t_L g682 ( .A(n_560), .B(n_683), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_562), .A2(n_693), .B(n_695), .C(n_698), .Y(n_692) );
AOI222xp33_ASAP7_75t_L g566 ( .A1(n_563), .A2(n_567), .B1(n_569), .B2(n_572), .C1(n_580), .C2(n_582), .Y(n_566) );
AND2x2_ASAP7_75t_L g634 ( .A(n_563), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g567 ( .A(n_564), .B(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g588 ( .A(n_564), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g565 ( .A(n_566), .B(n_585), .C(n_606), .D(n_616), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_568), .B(n_574), .Y(n_628) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g636 ( .A(n_571), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g643 ( .A(n_571), .Y(n_643) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
A2O1A1Ixp33_ASAP7_75t_L g606 ( .A1(n_573), .A2(n_607), .B(n_611), .C(n_615), .Y(n_606) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_574), .B(n_589), .Y(n_710) );
OR2x2_ASAP7_75t_L g714 ( .A(n_574), .B(n_600), .Y(n_714) );
INVx1_ASAP7_75t_L g687 ( .A(n_575), .Y(n_687) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_SL g621 ( .A(n_578), .Y(n_621) );
INVx1_ASAP7_75t_L g601 ( .A(n_579), .Y(n_601) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_581), .B(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g605 ( .A(n_583), .Y(n_605) );
AOI322xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_588), .A3(n_589), .B1(n_591), .B2(n_595), .C1(n_596), .C2(n_602), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
O2A1O1Ixp33_ASAP7_75t_SL g667 ( .A1(n_588), .A2(n_668), .B(n_669), .C(n_670), .Y(n_667) );
INVx1_ASAP7_75t_L g690 ( .A(n_589), .Y(n_690) );
NOR2xp67_ASAP7_75t_L g591 ( .A(n_592), .B(n_594), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g648 ( .A(n_594), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_600), .Y(n_670) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
INVx3_ASAP7_75t_L g613 ( .A(n_610), .Y(n_613) );
OR2x2_ASAP7_75t_L g681 ( .A(n_610), .B(n_643), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_610), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
INVx1_ASAP7_75t_SL g713 ( .A(n_614), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_615), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_SL g718 ( .A(n_623), .B(n_719), .C(n_721), .Y(n_718) );
NOR3xp33_ASAP7_75t_SL g624 ( .A(n_625), .B(n_662), .C(n_691), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_626), .B(n_644), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B(n_632), .C(n_638), .Y(n_626) );
OAI31xp33_ASAP7_75t_L g671 ( .A1(n_627), .A2(n_649), .A3(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx2_ASAP7_75t_L g686 ( .A(n_634), .Y(n_686) );
INVx1_ASAP7_75t_L g661 ( .A(n_636), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_641), .B(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OR2x2_ASAP7_75t_L g688 ( .A(n_646), .B(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_L g727 ( .A(n_647), .Y(n_727) );
OAI22xp33_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B1(n_657), .B2(n_661), .Y(n_650) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_656), .Y(n_668) );
OR2x2_ASAP7_75t_L g719 ( .A(n_656), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_671), .C(n_678), .Y(n_662) );
O2A1O1Ixp33_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B(n_666), .C(n_667), .Y(n_663) );
INVx2_ASAP7_75t_L g700 ( .A(n_664), .Y(n_700) );
INVx1_ASAP7_75t_SL g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_680), .B1(n_682), .B2(n_684), .C(n_685), .Y(n_678) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_687), .B1(n_688), .B2(n_690), .Y(n_685) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_701), .C(n_711), .Y(n_691) );
INVxp33_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g695 ( .A(n_696), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_702), .A2(n_704), .B1(n_707), .B2(n_709), .Y(n_701) );
INVx2_ASAP7_75t_L g715 ( .A(n_702), .Y(n_715) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_SL g722 ( .A1(n_721), .A2(n_723), .B1(n_724), .B2(n_725), .Y(n_722) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx4f_ASAP7_75t_SL g736 ( .A(n_728), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
CKINVDCx11_ASAP7_75t_R g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
AND2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_748), .Y(n_741) );
INVxp67_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_744), .B(n_747), .Y(n_743) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_SL g765 ( .A(n_745), .B(n_747), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_745), .A2(n_770), .B(n_773), .Y(n_769) );
INVx1_ASAP7_75t_SL g755 ( .A(n_748), .Y(n_755) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
BUFx3_ASAP7_75t_L g760 ( .A(n_749), .Y(n_760) );
BUFx2_ASAP7_75t_L g774 ( .A(n_749), .Y(n_774) );
INVxp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_754), .B(n_756), .Y(n_751) );
INVx1_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_SL g756 ( .A(n_757), .B(n_761), .Y(n_756) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
BUFx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx11_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx8_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
endmodule