module real_aes_7834_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g186 ( .A1(n_0), .A2(n_187), .B(n_188), .C(n_192), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_1), .B(n_181), .Y(n_194) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_3), .B(n_166), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_4), .A2(n_175), .B(n_481), .Y(n_480) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_5), .A2(n_155), .B(n_172), .C(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_6), .A2(n_175), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_7), .B(n_181), .Y(n_487) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_8), .A2(n_147), .B(n_269), .Y(n_268) );
AND2x6_ASAP7_75t_L g172 ( .A(n_9), .B(n_173), .Y(n_172) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_10), .A2(n_155), .B(n_172), .C(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g578 ( .A(n_11), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_40), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_12), .B(n_40), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_13), .B(n_191), .Y(n_527) );
INVx1_ASAP7_75t_L g152 ( .A(n_14), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_15), .B(n_166), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_16), .A2(n_167), .B(n_536), .C(n_538), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_17), .B(n_181), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_18), .B(n_209), .Y(n_501) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_19), .A2(n_155), .B(n_201), .C(n_208), .Y(n_200) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_20), .A2(n_190), .B(n_243), .C(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_21), .B(n_191), .Y(n_509) );
AOI222xp33_ASAP7_75t_L g456 ( .A1(n_22), .A2(n_457), .B1(n_726), .B2(n_727), .C1(n_736), .C2(n_740), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_23), .B(n_191), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g505 ( .A(n_24), .Y(n_505) );
INVx1_ASAP7_75t_L g475 ( .A(n_25), .Y(n_475) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_26), .A2(n_155), .B(n_208), .C(n_272), .Y(n_271) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_27), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_28), .Y(n_523) );
INVx1_ASAP7_75t_L g499 ( .A(n_29), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_30), .A2(n_175), .B(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_31), .B(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g157 ( .A(n_32), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_33), .A2(n_170), .B(n_224), .C(n_225), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_34), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_35), .A2(n_190), .B(n_484), .C(n_486), .Y(n_483) );
INVxp67_ASAP7_75t_L g500 ( .A(n_36), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_37), .B(n_274), .Y(n_273) );
CKINVDCx14_ASAP7_75t_R g482 ( .A(n_38), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g473 ( .A1(n_39), .A2(n_155), .B(n_208), .C(n_474), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_41), .A2(n_192), .B(n_576), .C(n_577), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_42), .B(n_199), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g246 ( .A(n_43), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_44), .B(n_166), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_45), .B(n_175), .Y(n_270) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_46), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_47), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_48), .A2(n_170), .B(n_224), .C(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g189 ( .A(n_49), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g133 ( .A1(n_50), .A2(n_67), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_50), .Y(n_135) );
INVx1_ASAP7_75t_L g253 ( .A(n_51), .Y(n_253) );
INVx1_ASAP7_75t_L g543 ( .A(n_52), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_53), .B(n_175), .Y(n_250) );
OAI22xp5_ASAP7_75t_SL g137 ( .A1(n_54), .A2(n_72), .B1(n_138), .B2(n_139), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_54), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_55), .Y(n_213) );
CKINVDCx14_ASAP7_75t_R g574 ( .A(n_56), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_57), .A2(n_105), .B1(n_118), .B2(n_743), .Y(n_104) );
INVx1_ASAP7_75t_L g173 ( .A(n_58), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_59), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_60), .B(n_181), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_61), .A2(n_162), .B(n_207), .C(n_264), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g732 ( .A1(n_62), .A2(n_71), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_62), .Y(n_733) );
INVx1_ASAP7_75t_L g151 ( .A(n_63), .Y(n_151) );
INVx1_ASAP7_75t_SL g485 ( .A(n_64), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_65), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_66), .B(n_166), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_67), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_67), .B(n_181), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_68), .B(n_167), .Y(n_240) );
INVx1_ASAP7_75t_L g508 ( .A(n_69), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_70), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_71), .Y(n_734) );
INVx1_ASAP7_75t_L g139 ( .A(n_72), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_73), .B(n_203), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_74), .A2(n_155), .B(n_160), .C(n_170), .Y(n_154) );
CKINVDCx16_ASAP7_75t_R g262 ( .A(n_75), .Y(n_262) );
INVx1_ASAP7_75t_L g117 ( .A(n_76), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_77), .A2(n_175), .B(n_573), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_78), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_79), .A2(n_175), .B(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_80), .A2(n_199), .B(n_495), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g472 ( .A(n_81), .Y(n_472) );
INVx1_ASAP7_75t_L g534 ( .A(n_82), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_83), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_83), .Y(n_730) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_84), .B(n_205), .Y(n_204) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_85), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_86), .A2(n_175), .B(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g537 ( .A(n_87), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_88), .A2(n_728), .B1(n_729), .B2(n_735), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_88), .Y(n_728) );
INVx2_ASAP7_75t_L g149 ( .A(n_89), .Y(n_149) );
INVx1_ASAP7_75t_L g526 ( .A(n_90), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_91), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_92), .B(n_191), .Y(n_241) );
INVx2_ASAP7_75t_L g114 ( .A(n_93), .Y(n_114) );
OR2x2_ASAP7_75t_L g128 ( .A(n_93), .B(n_129), .Y(n_128) );
OR2x2_ASAP7_75t_L g461 ( .A(n_93), .B(n_130), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_94), .A2(n_155), .B(n_170), .C(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_95), .B(n_175), .Y(n_222) );
INVx1_ASAP7_75t_L g226 ( .A(n_96), .Y(n_226) );
INVxp67_ASAP7_75t_L g265 ( .A(n_97), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_98), .B(n_147), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_99), .B(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g161 ( .A(n_100), .Y(n_161) );
INVx1_ASAP7_75t_L g236 ( .A(n_101), .Y(n_236) );
INVx2_ASAP7_75t_L g546 ( .A(n_102), .Y(n_546) );
AND2x2_ASAP7_75t_L g255 ( .A(n_103), .B(n_211), .Y(n_255) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g743 ( .A(n_107), .Y(n_743) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .C(n_115), .Y(n_112) );
AND2x2_ASAP7_75t_L g130 ( .A(n_113), .B(n_131), .Y(n_130) );
OR2x2_ASAP7_75t_L g725 ( .A(n_114), .B(n_130), .Y(n_725) );
NOR2x2_ASAP7_75t_L g742 ( .A(n_114), .B(n_129), .Y(n_742) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_124), .B(n_455), .Y(n_118) );
BUFx2_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
NAND3xp33_ASAP7_75t_L g455 ( .A(n_120), .B(n_452), .C(n_456), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_132), .B(n_452), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_SL g127 ( .A(n_128), .Y(n_127) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_128), .Y(n_454) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AOI22xp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_136), .B1(n_450), .B2(n_451), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_133), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_136), .Y(n_451) );
XNOR2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_140), .Y(n_136) );
INVx1_ASAP7_75t_L g458 ( .A(n_140), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g736 ( .A1(n_140), .A2(n_463), .B1(n_737), .B2(n_738), .Y(n_736) );
OR3x1_ASAP7_75t_L g140 ( .A(n_141), .B(n_358), .C(n_407), .Y(n_140) );
NAND5xp2_ASAP7_75t_L g141 ( .A(n_142), .B(n_292), .C(n_321), .D(n_329), .E(n_344), .Y(n_141) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_215), .B(n_231), .C(n_276), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_195), .Y(n_143) );
AND2x2_ASAP7_75t_L g287 ( .A(n_144), .B(n_284), .Y(n_287) );
AND2x2_ASAP7_75t_L g320 ( .A(n_144), .B(n_196), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_144), .B(n_219), .Y(n_413) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_180), .Y(n_144) );
INVx2_ASAP7_75t_L g218 ( .A(n_145), .Y(n_218) );
BUFx2_ASAP7_75t_L g387 ( .A(n_145), .Y(n_387) );
AO21x2_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_153), .B(n_178), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_146), .B(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g181 ( .A(n_146), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_146), .B(n_230), .Y(n_229) );
AO21x2_ASAP7_75t_L g234 ( .A1(n_146), .A2(n_235), .B(n_245), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_146), .B(n_478), .Y(n_477) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_146), .A2(n_504), .B(n_511), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_146), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_147), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_147), .A2(n_270), .B(n_271), .Y(n_269) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g247 ( .A(n_148), .Y(n_247) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
AND2x2_ASAP7_75t_SL g211 ( .A(n_149), .B(n_150), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_174), .Y(n_153) );
INVx5_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
BUFx3_ASAP7_75t_L g193 ( .A(n_156), .Y(n_193) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g177 ( .A(n_157), .Y(n_177) );
INVx1_ASAP7_75t_L g244 ( .A(n_157), .Y(n_244) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_159), .Y(n_164) );
INVx3_ASAP7_75t_L g167 ( .A(n_159), .Y(n_167) );
AND2x2_ASAP7_75t_L g176 ( .A(n_159), .B(n_177), .Y(n_176) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVx1_ASAP7_75t_L g274 ( .A(n_159), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_165), .C(n_168), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp33_ASAP7_75t_L g498 ( .A1(n_163), .A2(n_166), .B1(n_499), .B2(n_500), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_163), .B(n_537), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_163), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
INVx2_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_166), .B(n_265), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g474 ( .A1(n_166), .A2(n_206), .B(n_475), .C(n_476), .Y(n_474) );
INVx5_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_167), .B(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx3_ASAP7_75t_L g486 ( .A(n_169), .Y(n_486) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g183 ( .A1(n_171), .A2(n_184), .B(n_185), .C(n_186), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_171), .A2(n_185), .B(n_262), .C(n_263), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g481 ( .A1(n_171), .A2(n_185), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g495 ( .A1(n_171), .A2(n_185), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_171), .A2(n_185), .B(n_534), .C(n_535), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_SL g542 ( .A1(n_171), .A2(n_185), .B(n_543), .C(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_SL g573 ( .A1(n_171), .A2(n_185), .B(n_574), .C(n_575), .Y(n_573) );
INVx4_ASAP7_75t_SL g171 ( .A(n_172), .Y(n_171) );
AND2x4_ASAP7_75t_L g175 ( .A(n_172), .B(n_176), .Y(n_175) );
BUFx3_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_172), .B(n_176), .Y(n_237) );
BUFx2_ASAP7_75t_L g199 ( .A(n_175), .Y(n_199) );
INVx1_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
AND2x2_ASAP7_75t_L g195 ( .A(n_180), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g285 ( .A(n_180), .Y(n_285) );
AND2x2_ASAP7_75t_L g371 ( .A(n_180), .B(n_284), .Y(n_371) );
AND2x2_ASAP7_75t_L g426 ( .A(n_180), .B(n_218), .Y(n_426) );
OA21x2_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_194), .Y(n_180) );
INVx2_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_190), .B(n_485), .Y(n_484) );
INVx4_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g576 ( .A(n_191), .Y(n_576) );
INVx2_ASAP7_75t_L g510 ( .A(n_192), .Y(n_510) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_193), .Y(n_228) );
INVx1_ASAP7_75t_L g538 ( .A(n_193), .Y(n_538) );
INVx1_ASAP7_75t_L g343 ( .A(n_195), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_195), .B(n_219), .Y(n_390) );
INVx5_ASAP7_75t_L g284 ( .A(n_196), .Y(n_284) );
AND2x4_ASAP7_75t_L g305 ( .A(n_196), .B(n_285), .Y(n_305) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_196), .Y(n_327) );
AND2x2_ASAP7_75t_L g402 ( .A(n_196), .B(n_387), .Y(n_402) );
AND2x2_ASAP7_75t_L g405 ( .A(n_196), .B(n_220), .Y(n_405) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_212), .Y(n_196) );
AOI21xp5_ASAP7_75t_SL g197 ( .A1(n_198), .A2(n_200), .B(n_209), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B(n_206), .Y(n_201) );
INVx2_ASAP7_75t_L g205 ( .A(n_203), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_205), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g252 ( .A1(n_205), .A2(n_228), .B(n_253), .C(n_254), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_205), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
O2A1O1Ixp5_ASAP7_75t_L g525 ( .A1(n_205), .A2(n_510), .B(n_526), .C(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_207), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_210), .B(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g214 ( .A(n_211), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_211), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_211), .A2(n_250), .B(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g471 ( .A1(n_211), .A2(n_237), .B(n_472), .C(n_473), .Y(n_471) );
OA21x2_ASAP7_75t_L g571 ( .A1(n_211), .A2(n_572), .B(n_579), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_214), .A2(n_522), .B(n_528), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_215), .B(n_285), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_215), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_219), .Y(n_216) );
AND2x2_ASAP7_75t_L g310 ( .A(n_217), .B(n_285), .Y(n_310) );
AND2x2_ASAP7_75t_L g328 ( .A(n_217), .B(n_220), .Y(n_328) );
INVx1_ASAP7_75t_L g348 ( .A(n_217), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_217), .B(n_284), .Y(n_393) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_217), .Y(n_435) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_218), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_219), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_219), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_219), .A2(n_280), .B(n_341), .C(n_343), .Y(n_340) );
AND2x2_ASAP7_75t_L g347 ( .A(n_219), .B(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g356 ( .A(n_219), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g360 ( .A(n_219), .B(n_284), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_219), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g375 ( .A(n_219), .B(n_285), .Y(n_375) );
AND2x2_ASAP7_75t_L g425 ( .A(n_219), .B(n_426), .Y(n_425) );
INVx5_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx2_ASAP7_75t_L g289 ( .A(n_220), .Y(n_289) );
AND2x2_ASAP7_75t_L g330 ( .A(n_220), .B(n_283), .Y(n_330) );
AND2x2_ASAP7_75t_L g342 ( .A(n_220), .B(n_317), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_220), .B(n_371), .Y(n_389) );
OR2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_229), .Y(n_220) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_256), .Y(n_231) );
INVx1_ASAP7_75t_L g278 ( .A(n_232), .Y(n_278) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_248), .Y(n_232) );
OR2x2_ASAP7_75t_L g280 ( .A(n_233), .B(n_248), .Y(n_280) );
NAND3xp33_ASAP7_75t_L g286 ( .A(n_233), .B(n_287), .C(n_288), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_233), .B(n_258), .Y(n_297) );
OR2x2_ASAP7_75t_L g312 ( .A(n_233), .B(n_300), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_233), .B(n_267), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_233), .B(n_449), .Y(n_448) );
INVx5_ASAP7_75t_SL g233 ( .A(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_234), .B(n_258), .Y(n_315) );
AND2x2_ASAP7_75t_L g354 ( .A(n_234), .B(n_268), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_234), .B(n_267), .Y(n_382) );
OR2x2_ASAP7_75t_L g385 ( .A(n_234), .B(n_267), .Y(n_385) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_238), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_237), .A2(n_505), .B(n_506), .Y(n_504) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_237), .A2(n_523), .B(n_524), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_241), .B(n_242), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_273), .B(n_275), .Y(n_272) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g493 ( .A(n_247), .Y(n_493) );
INVx5_ASAP7_75t_SL g300 ( .A(n_248), .Y(n_300) );
OR2x2_ASAP7_75t_L g306 ( .A(n_248), .B(n_257), .Y(n_306) );
AND2x2_ASAP7_75t_L g322 ( .A(n_248), .B(n_323), .Y(n_322) );
AOI321xp33_ASAP7_75t_L g329 ( .A1(n_248), .A2(n_330), .A3(n_331), .B1(n_332), .B2(n_338), .C(n_340), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_248), .B(n_256), .Y(n_339) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_248), .Y(n_352) );
OR2x2_ASAP7_75t_L g399 ( .A(n_248), .B(n_297), .Y(n_399) );
AND2x2_ASAP7_75t_L g421 ( .A(n_248), .B(n_318), .Y(n_421) );
AND2x2_ASAP7_75t_L g440 ( .A(n_248), .B(n_258), .Y(n_440) );
OR2x6_ASAP7_75t_L g248 ( .A(n_249), .B(n_255), .Y(n_248) );
INVx1_ASAP7_75t_SL g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_267), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_258), .B(n_267), .Y(n_281) );
AND2x2_ASAP7_75t_L g290 ( .A(n_258), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g317 ( .A(n_258), .Y(n_317) );
AND2x2_ASAP7_75t_L g323 ( .A(n_258), .B(n_318), .Y(n_323) );
INVxp67_ASAP7_75t_L g353 ( .A(n_258), .Y(n_353) );
OR2x2_ASAP7_75t_L g395 ( .A(n_258), .B(n_300), .Y(n_395) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_266), .Y(n_258) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_259), .A2(n_480), .B(n_487), .Y(n_479) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_259), .A2(n_532), .B(n_539), .Y(n_531) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_259), .A2(n_541), .B(n_547), .Y(n_540) );
OR2x2_ASAP7_75t_L g277 ( .A(n_267), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g291 ( .A(n_267), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_267), .B(n_280), .Y(n_324) );
AND2x2_ASAP7_75t_L g373 ( .A(n_267), .B(n_317), .Y(n_373) );
AND2x2_ASAP7_75t_L g411 ( .A(n_267), .B(n_300), .Y(n_411) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_268), .B(n_300), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .B(n_282), .C(n_286), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_277), .A2(n_279), .B1(n_404), .B2(n_406), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_279), .A2(n_302), .B1(n_357), .B2(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_SL g431 ( .A(n_280), .Y(n_431) );
INVx1_ASAP7_75t_SL g331 ( .A(n_281), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_283), .B(n_303), .Y(n_333) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_283), .A2(n_324), .B1(n_331), .B2(n_345), .C1(n_349), .C2(n_355), .Y(n_344) );
AND2x2_ASAP7_75t_L g434 ( .A(n_283), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g309 ( .A(n_284), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_284), .B(n_304), .Y(n_379) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_284), .Y(n_416) );
AND2x2_ASAP7_75t_L g419 ( .A(n_284), .B(n_328), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_284), .B(n_435), .Y(n_445) );
INVx1_ASAP7_75t_L g336 ( .A(n_285), .Y(n_336) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_285), .Y(n_364) );
O2A1O1Ixp33_ASAP7_75t_L g427 ( .A1(n_287), .A2(n_428), .B(n_429), .C(n_432), .Y(n_427) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g350 ( .A(n_289), .B(n_351), .C(n_354), .Y(n_350) );
OR2x2_ASAP7_75t_L g378 ( .A(n_289), .B(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_289), .B(n_305), .Y(n_406) );
OR2x2_ASAP7_75t_L g311 ( .A(n_291), .B(n_312), .Y(n_311) );
AOI211xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_295), .B(n_301), .C(n_313), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_294), .B(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g400 ( .A(n_295), .B(n_401), .Y(n_400) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_296), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g314 ( .A(n_299), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_300), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g368 ( .A(n_300), .B(n_318), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_300), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_300), .B(n_317), .Y(n_383) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_306), .B1(n_307), .B2(n_311), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_303), .B(n_375), .Y(n_374) );
BUFx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_305), .B(n_347), .Y(n_346) );
OAI221xp5_ASAP7_75t_SL g369 ( .A1(n_306), .A2(n_370), .B1(n_372), .B2(n_374), .C(n_376), .Y(n_369) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g424 ( .A(n_309), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g437 ( .A(n_309), .B(n_426), .Y(n_437) );
INVx1_ASAP7_75t_L g357 ( .A(n_310), .Y(n_357) );
INVx1_ASAP7_75t_L g428 ( .A(n_311), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_312), .A2(n_395), .B(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_316), .B(n_319), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
OAI21xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_324), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g361 ( .A(n_322), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_323), .A2(n_409), .B1(n_412), .B2(n_414), .C(n_417), .Y(n_408) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_331), .A2(n_421), .B1(n_422), .B2(n_424), .Y(n_420) );
NAND2xp5_ASAP7_75t_SL g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g397 ( .A(n_333), .Y(n_397) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NOR2xp67_ASAP7_75t_SL g335 ( .A(n_336), .B(n_337), .Y(n_335) );
AND2x2_ASAP7_75t_L g401 ( .A(n_337), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g366 ( .A(n_342), .Y(n_366) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_347), .B(n_371), .Y(n_423) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_353), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g439 ( .A(n_354), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g446 ( .A(n_354), .B(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI211xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_362), .C(n_396), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_369), .C(n_388), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g449 ( .A(n_373), .Y(n_449) );
AND2x2_ASAP7_75t_L g386 ( .A(n_375), .B(n_387), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B1(n_384), .B2(n_386), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
OR2x2_ASAP7_75t_L g394 ( .A(n_382), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g447 ( .A(n_383), .Y(n_447) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI31xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .A3(n_391), .B(n_394), .Y(n_388) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_398), .B(n_400), .C(n_403), .Y(n_396) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_405), .Y(n_404) );
NAND5xp2_ASAP7_75t_L g407 ( .A(n_408), .B(n_420), .C(n_427), .D(n_441), .E(n_444), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_419), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_444) );
INVx1_ASAP7_75t_SL g443 ( .A(n_421), .Y(n_443) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AOI21xp33_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_436), .B(n_438), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
OAI22xp5_ASAP7_75t_SL g457 ( .A1(n_458), .A2(n_459), .B1(n_462), .B2(n_725), .Y(n_457) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g737 ( .A(n_460), .Y(n_737) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR3x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_636), .C(n_683), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_582), .C(n_607), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_520), .B1(n_548), .B2(n_551), .C(n_559), .Y(n_465) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_488), .B(n_513), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_468), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_468), .B(n_564), .Y(n_680) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_479), .Y(n_468) );
AND2x2_ASAP7_75t_L g550 ( .A(n_469), .B(n_519), .Y(n_550) );
AND2x2_ASAP7_75t_L g600 ( .A(n_469), .B(n_518), .Y(n_600) );
AND2x2_ASAP7_75t_L g621 ( .A(n_469), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g626 ( .A(n_469), .B(n_593), .Y(n_626) );
OR2x2_ASAP7_75t_L g634 ( .A(n_469), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g706 ( .A(n_469), .B(n_502), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_469), .B(n_655), .Y(n_720) );
INVx3_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g565 ( .A(n_470), .B(n_479), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_470), .B(n_502), .Y(n_566) );
AND2x4_ASAP7_75t_L g588 ( .A(n_470), .B(n_519), .Y(n_588) );
AND2x2_ASAP7_75t_L g618 ( .A(n_470), .B(n_490), .Y(n_618) );
AND2x2_ASAP7_75t_L g627 ( .A(n_470), .B(n_617), .Y(n_627) );
AND2x2_ASAP7_75t_L g643 ( .A(n_470), .B(n_503), .Y(n_643) );
OR2x2_ASAP7_75t_L g652 ( .A(n_470), .B(n_635), .Y(n_652) );
AND2x2_ASAP7_75t_L g658 ( .A(n_470), .B(n_593), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_470), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g672 ( .A(n_470), .B(n_515), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_470), .B(n_561), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_470), .B(n_622), .Y(n_711) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_477), .Y(n_470) );
INVx2_ASAP7_75t_L g519 ( .A(n_479), .Y(n_519) );
AND2x2_ASAP7_75t_L g617 ( .A(n_479), .B(n_502), .Y(n_617) );
AND2x2_ASAP7_75t_L g622 ( .A(n_479), .B(n_503), .Y(n_622) );
INVx1_ASAP7_75t_L g678 ( .A(n_479), .Y(n_678) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g587 ( .A(n_489), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_502), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_490), .B(n_550), .Y(n_549) );
BUFx3_ASAP7_75t_L g564 ( .A(n_490), .Y(n_564) );
OR2x2_ASAP7_75t_L g635 ( .A(n_490), .B(n_502), .Y(n_635) );
OR2x2_ASAP7_75t_L g696 ( .A(n_490), .B(n_603), .Y(n_696) );
OA21x2_ASAP7_75t_L g490 ( .A1(n_491), .A2(n_494), .B(n_501), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_492), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g516 ( .A(n_494), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_501), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_502), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g655 ( .A(n_502), .B(n_515), .Y(n_655) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_514), .A2(n_700), .B1(n_704), .B2(n_707), .C(n_708), .Y(n_699) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_518), .Y(n_514) );
INVx1_ASAP7_75t_SL g562 ( .A(n_515), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_515), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g694 ( .A(n_515), .B(n_550), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_518), .B(n_564), .Y(n_686) );
AND2x2_ASAP7_75t_L g593 ( .A(n_519), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_SL g597 ( .A(n_520), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_520), .B(n_603), .Y(n_633) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g558 ( .A(n_521), .B(n_531), .Y(n_558) );
INVx4_ASAP7_75t_L g570 ( .A(n_521), .Y(n_570) );
BUFx3_ASAP7_75t_L g613 ( .A(n_521), .Y(n_613) );
AND3x2_ASAP7_75t_L g628 ( .A(n_521), .B(n_629), .C(n_630), .Y(n_628) );
AND2x2_ASAP7_75t_L g710 ( .A(n_530), .B(n_624), .Y(n_710) );
AND2x2_ASAP7_75t_L g718 ( .A(n_530), .B(n_603), .Y(n_718) );
INVx1_ASAP7_75t_SL g723 ( .A(n_530), .Y(n_723) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_540), .Y(n_530) );
INVx1_ASAP7_75t_SL g581 ( .A(n_531), .Y(n_581) );
AND2x2_ASAP7_75t_L g604 ( .A(n_531), .B(n_570), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_531), .B(n_554), .Y(n_606) );
HB1xp67_ASAP7_75t_L g646 ( .A(n_531), .Y(n_646) );
OR2x2_ASAP7_75t_L g651 ( .A(n_531), .B(n_570), .Y(n_651) );
INVx2_ASAP7_75t_L g556 ( .A(n_540), .Y(n_556) );
AND2x2_ASAP7_75t_L g591 ( .A(n_540), .B(n_571), .Y(n_591) );
OR2x2_ASAP7_75t_L g611 ( .A(n_540), .B(n_571), .Y(n_611) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_540), .Y(n_631) );
INVx1_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_549), .A2(n_590), .B(n_682), .Y(n_681) );
AOI322xp5_ASAP7_75t_L g717 ( .A1(n_551), .A2(n_561), .A3(n_588), .B1(n_718), .B2(n_719), .C1(n_721), .C2(n_724), .Y(n_717) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_553), .B(n_557), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_553), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_554), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g580 ( .A(n_555), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g648 ( .A(n_556), .B(n_570), .Y(n_648) );
AND2x2_ASAP7_75t_L g715 ( .A(n_556), .B(n_571), .Y(n_715) );
INVx1_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g656 ( .A(n_558), .B(n_610), .Y(n_656) );
AOI31xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_563), .A3(n_566), .B(n_567), .Y(n_559) );
AND2x2_ASAP7_75t_L g615 ( .A(n_561), .B(n_593), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_561), .B(n_585), .Y(n_697) );
AND2x2_ASAP7_75t_L g716 ( .A(n_561), .B(n_621), .Y(n_716) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_564), .B(n_593), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g639 ( .A(n_564), .B(n_622), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_564), .B(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_564), .B(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_565), .B(n_622), .Y(n_654) );
INVx1_ASAP7_75t_L g698 ( .A(n_565), .Y(n_698) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_580), .Y(n_568) );
INVxp67_ASAP7_75t_L g650 ( .A(n_569), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_570), .B(n_581), .Y(n_586) );
INVx1_ASAP7_75t_L g692 ( .A(n_570), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_570), .B(n_669), .Y(n_703) );
BUFx3_ASAP7_75t_L g603 ( .A(n_571), .Y(n_603) );
AND2x2_ASAP7_75t_L g629 ( .A(n_571), .B(n_581), .Y(n_629) );
INVx2_ASAP7_75t_L g669 ( .A(n_571), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_580), .B(n_702), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_587), .B(n_589), .C(n_598), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_584), .A2(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_585), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_585), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g665 ( .A(n_586), .B(n_611), .Y(n_665) );
INVx3_ASAP7_75t_L g596 ( .A(n_588), .Y(n_596) );
OAI22xp5_ASAP7_75t_SL g589 ( .A1(n_590), .A2(n_592), .B1(n_595), .B2(n_597), .Y(n_589) );
OAI21xp5_ASAP7_75t_SL g614 ( .A1(n_591), .A2(n_615), .B(n_616), .Y(n_614) );
AND2x2_ASAP7_75t_L g640 ( .A(n_591), .B(n_604), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_591), .B(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OR2x2_ASAP7_75t_L g595 ( .A(n_594), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g664 ( .A(n_594), .Y(n_664) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_595), .A2(n_609), .B(n_614), .Y(n_608) );
OAI22xp33_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_601), .B1(n_605), .B2(n_606), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_600), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
INVx1_ASAP7_75t_L g624 ( .A(n_603), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_603), .B(n_646), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_619), .C(n_632), .Y(n_607) );
OAI22xp5_ASAP7_75t_SL g674 ( .A1(n_609), .A2(n_675), .B1(n_679), .B2(n_680), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
OR2x2_ASAP7_75t_L g679 ( .A(n_611), .B(n_612), .Y(n_679) );
AND2x2_ASAP7_75t_L g687 ( .A(n_612), .B(n_668), .Y(n_687) );
CKINVDCx16_ASAP7_75t_R g612 ( .A(n_613), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_SL g695 ( .A1(n_613), .A2(n_696), .B(n_697), .C(n_698), .Y(n_695) );
OR2x2_ASAP7_75t_L g722 ( .A(n_613), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_625), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_621), .A2(n_658), .B(n_659), .C(n_662), .Y(n_657) );
OAI21xp33_ASAP7_75t_SL g625 ( .A1(n_626), .A2(n_627), .B(n_628), .Y(n_625) );
AND2x2_ASAP7_75t_L g690 ( .A(n_629), .B(n_648), .Y(n_690) );
INVxp67_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g668 ( .A(n_631), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g673 ( .A(n_633), .Y(n_673) );
NAND3xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_657), .C(n_670), .Y(n_636) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_641), .C(n_649), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
INVx1_ASAP7_75t_L g707 ( .A(n_644), .Y(n_707) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_L g667 ( .A(n_646), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_646), .B(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
A2O1A1Ixp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B(n_652), .C(n_653), .Y(n_649) );
INVx2_ASAP7_75t_SL g661 ( .A(n_651), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_652), .A2(n_663), .B1(n_665), .B2(n_666), .Y(n_662) );
OAI21xp33_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_673), .B(n_674), .C(n_681), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVxp33_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g724 ( .A(n_678), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g683 ( .A(n_684), .B(n_699), .C(n_712), .D(n_717), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_685), .A2(n_687), .B(n_688), .C(n_695), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_693), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g708 ( .A1(n_689), .A2(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_696), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_716), .Y(n_712) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g739 ( .A(n_725), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_727), .Y(n_726) );
CKINVDCx16_ASAP7_75t_R g735 ( .A(n_729), .Y(n_735) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_SL g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
endmodule