module fake_jpeg_10161_n_77 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_18),
.B1(n_33),
.B2(n_4),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_54),
.Y(n_63)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_0),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_58),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_45),
.Y(n_62)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_38),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_22),
.B1(n_5),
.B2(n_7),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_10),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_1),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_64),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_46),
.C(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_59),
.C(n_66),
.Y(n_71)
);

A2O1A1O1Ixp25_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_63),
.B(n_57),
.C(n_67),
.D(n_40),
.Y(n_72)
);

NOR3xp33_ASAP7_75t_SL g73 ( 
.A(n_72),
.B(n_39),
.C(n_36),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_73),
.A2(n_60),
.B1(n_13),
.B2(n_16),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_11),
.B(n_17),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_23),
.A3(n_25),
.B1(n_27),
.B2(n_28),
.C1(n_29),
.C2(n_31),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_34),
.Y(n_77)
);


endmodule