module fake_jpeg_4844_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_28;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx2_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx10_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_18),
.Y(n_27)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_10),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_20),
.Y(n_23)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_25),
.A2(n_10),
.B(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_8),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_21),
.B1(n_14),
.B2(n_11),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_33),
.C(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_10),
.B1(n_16),
.B2(n_13),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_35),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_22),
.B1(n_16),
.B2(n_12),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_37),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_46),
.B1(n_28),
.B2(n_40),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_34),
.B1(n_28),
.B2(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_41),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_43),
.C(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_46),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_51),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_50),
.C(n_6),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.C(n_6),
.Y(n_56)
);

BUFx24_ASAP7_75t_SL g57 ( 
.A(n_56),
.Y(n_57)
);


endmodule