module fake_aes_9523_n_902 (n_120, n_107, n_103, n_52, n_114, n_50, n_7, n_3, n_34, n_25, n_9, n_96, n_72, n_77, n_90, n_99, n_43, n_73, n_62, n_97, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_66, n_88, n_46, n_121, n_108, n_37, n_122, n_18, n_65, n_87, n_5, n_81, n_85, n_112, n_102, n_47, n_109, n_1, n_16, n_78, n_95, n_40, n_68, n_105, n_36, n_11, n_115, n_15, n_71, n_117, n_70, n_94, n_2, n_17, n_58, n_113, n_20, n_84, n_12, n_56, n_80, n_67, n_116, n_22, n_118, n_19, n_26, n_39, n_101, n_98, n_38, n_104, n_100, n_24, n_35, n_91, n_32, n_93, n_48, n_63, n_54, n_41, n_55, n_29, n_60, n_111, n_10, n_30, n_13, n_92, n_75, n_82, n_53, n_64, n_69, n_83, n_23, n_0, n_110, n_119, n_57, n_51, n_106, n_45, n_42, n_21, n_86, n_27, n_89, n_28, n_79, n_49, n_14, n_31, n_902, n_901);
input n_120;
input n_107;
input n_103;
input n_52;
input n_114;
input n_50;
input n_7;
input n_3;
input n_34;
input n_25;
input n_9;
input n_96;
input n_72;
input n_77;
input n_90;
input n_99;
input n_43;
input n_73;
input n_62;
input n_97;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_66;
input n_88;
input n_46;
input n_121;
input n_108;
input n_37;
input n_122;
input n_18;
input n_65;
input n_87;
input n_5;
input n_81;
input n_85;
input n_112;
input n_102;
input n_47;
input n_109;
input n_1;
input n_16;
input n_78;
input n_95;
input n_40;
input n_68;
input n_105;
input n_36;
input n_11;
input n_115;
input n_15;
input n_71;
input n_117;
input n_70;
input n_94;
input n_2;
input n_17;
input n_58;
input n_113;
input n_20;
input n_84;
input n_12;
input n_56;
input n_80;
input n_67;
input n_116;
input n_22;
input n_118;
input n_19;
input n_26;
input n_39;
input n_101;
input n_98;
input n_38;
input n_104;
input n_100;
input n_24;
input n_35;
input n_91;
input n_32;
input n_93;
input n_48;
input n_63;
input n_54;
input n_41;
input n_55;
input n_29;
input n_60;
input n_111;
input n_10;
input n_30;
input n_13;
input n_92;
input n_75;
input n_82;
input n_53;
input n_64;
input n_69;
input n_83;
input n_23;
input n_0;
input n_110;
input n_119;
input n_57;
input n_51;
input n_106;
input n_45;
input n_42;
input n_21;
input n_86;
input n_27;
input n_89;
input n_28;
input n_79;
input n_49;
input n_14;
input n_31;
output n_902;
output n_901;
wire n_890;
wire n_646;
wire n_107;
wire n_759;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_895;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_769;
wire n_169;
wire n_370;
wire n_439;
wire n_545;
wire n_384;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_831;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_394;
wire n_44;
wire n_189;
wire n_681;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_535;
wire n_689;
wire n_886;
wire n_595;
wire n_875;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_850;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_753;
wire n_859;
wire n_436;
wire n_438;
wire n_869;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_833;
wire n_405;
wire n_830;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_838;
wire n_569;
wire n_534;
wire n_707;
wire n_526;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_864;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_876;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_553;
wire n_555;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_880;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_836;
wire n_127;
wire n_312;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_887;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_806;
wire n_155;
wire n_162;
wire n_114;
wire n_772;
wire n_50;
wire n_789;
wire n_816;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_882;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_884;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_699;
wire n_857;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_883;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_868;
wire n_628;
wire n_425;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_332;
wire n_109;
wire n_198;
wire n_386;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_863;
wire n_671;
wire n_892;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_765;
wire n_829;
wire n_599;
wire n_715;
wire n_849;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_837;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_851;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_855;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_800;
wire n_491;
wire n_711;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_679;
wire n_522;
wire n_546;
wire n_615;
wire n_684;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_879;
wire n_888;
wire n_576;
wire n_275;
wire n_691;
wire n_622;
wire n_661;
wire n_493;
wire n_274;
wire n_235;
wire n_150;
wire n_690;
wire n_533;
wire n_38;
wire n_272;
wire n_686;
wire n_100;
wire n_299;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_844;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_878;
wire n_783;
wire n_812;
wire n_147;
wire n_185;
wire n_367;
wire n_795;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_873;
wire n_899;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_779;
wire n_212;
wire n_746;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_728;
wire n_435;
wire n_704;
wire n_583;
wire n_841;
wire n_64;
wire n_69;
wire n_248;
wire n_866;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_119;
wire n_667;
wire n_503;
wire n_856;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_163;
wire n_348;
wire n_762;
wire n_669;
wire n_685;
wire n_77;
wire n_90;
wire n_72;
wire n_594;
wire n_787;
wire n_214;
wire n_96;
wire n_770;
wire n_167;
wire n_861;
wire n_809;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_224;
wire n_161;
wire n_484;
wire n_165;
wire n_860;
wire n_413;
wire n_537;
wire n_710;
wire n_65;
wire n_560;
wire n_525;
wire n_5;
wire n_496;
wire n_393;
wire n_843;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_846;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_792;
wire n_277;
wire n_259;
wire n_885;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_827;
wire n_297;
wire n_276;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_815;
wire n_523;
wire n_854;
wire n_901;
wire n_528;
wire n_419;
wire n_252;
wire n_519;
wire n_168;
wire n_839;
wire n_271;
wire n_693;
wire n_785;
wire n_896;
wire n_739;
wire n_94;
wire n_194;
wire n_858;
wire n_758;
wire n_825;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_321;
wire n_284;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_597;
wire n_554;
wire n_741;
wire n_698;
wire n_257;
wire n_705;
wire n_828;
wire n_722;
wire n_203;
wire n_26;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_146;
wire n_337;
wire n_637;
wire n_32;
wire n_641;
wire n_726;
wire n_531;
wire n_872;
wire n_93;
wire n_539;
wire n_847;
wire n_406;
wire n_372;
wire n_842;
wire n_820;
wire n_713;
wire n_467;
wire n_702;
wire n_41;
wire n_760;
wire n_826;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_898;
wire n_647;
wire n_445;
wire n_500;
wire n_732;
wire n_845;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_834;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_835;
wire n_437;
wire n_871;
wire n_620;
wire n_89;
wire n_480;
wire n_130;
wire n_310;
wire n_341;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_136;
wire n_260;
wire n_891;
wire n_580;
wire n_610;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_142;
wire n_34;
wire n_853;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_781;
wire n_852;
wire n_376;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_88;
wire n_568;
wire n_46;
wire n_174;
wire n_717;
wire n_807;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_865;
wire n_672;
wire n_867;
wire n_466;
wire n_87;
wire n_207;
wire n_197;
wire n_81;
wire n_572;
wire n_541;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_416;
wire n_36;
wire n_870;
wire n_889;
wire n_432;
wire n_465;
wire n_414;
wire n_730;
wire n_680;
wire n_369;
wire n_469;
wire n_361;
wire n_767;
wire n_237;
wire n_881;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_803;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_804;
wire n_796;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_591;
wire n_391;
wire n_209;
wire n_241;
wire n_874;
wire n_84;
wire n_20;
wire n_782;
wire n_449;
wire n_832;
wire n_12;
wire n_56;
wire n_412;
wire n_455;
wire n_504;
wire n_618;
wire n_67;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_877;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_862;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_472;
wire n_490;
wire n_540;
wire n_840;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_893;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_894;
wire n_138;
wire n_60;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_745;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_505;
wire n_313;
wire n_358;
wire n_333;
wire n_627;
wire n_750;
wire n_706;
wire n_740;
wire n_589;
wire n_92;
wire n_175;
wire n_897;
wire n_128;
wire n_306;
wire n_415;
wire n_31;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_642;
wire n_675;
wire n_234;
wire n_607;
wire n_848;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_738;
wire n_27;
wire n_86;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_349;
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_81), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_77), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_9), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_17), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_71), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_62), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_15), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
NOR2xp67_ASAP7_75t_L g134 ( .A(n_98), .B(n_69), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_49), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_4), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_47), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_13), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_122), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_73), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_93), .Y(n_143) );
INVx2_ASAP7_75t_SL g144 ( .A(n_21), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_106), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_37), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_30), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_61), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_59), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_3), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_56), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_91), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_90), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_100), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_42), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_113), .Y(n_157) );
BUFx10_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_85), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_104), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_95), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_1), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_9), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_33), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_103), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_19), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_4), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_115), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_16), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_84), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_11), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_35), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_25), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_139), .Y(n_177) );
BUFx2_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_139), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_167), .B(n_0), .Y(n_180) );
INVx6_ASAP7_75t_L g181 ( .A(n_158), .Y(n_181) );
INVx5_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_144), .B(n_125), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_130), .Y(n_185) );
BUFx2_ASAP7_75t_L g186 ( .A(n_168), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_144), .B(n_0), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_124), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
OA21x2_ASAP7_75t_L g191 ( .A1(n_127), .A2(n_53), .B(n_120), .Y(n_191) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_131), .A2(n_52), .B(n_119), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_158), .B(n_1), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_170), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_123), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_129), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g198 ( .A(n_182), .B(n_123), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_190), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_177), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_186), .B(n_168), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_183), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_183), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_190), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
NAND2xp33_ASAP7_75t_SL g206 ( .A(n_193), .B(n_135), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_182), .B(n_128), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_195), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_177), .Y(n_209) );
AND2x2_ASAP7_75t_SL g210 ( .A(n_191), .B(n_142), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_195), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_177), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_177), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_182), .B(n_128), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_182), .B(n_149), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_180), .A2(n_148), .B1(n_135), .B2(n_126), .Y(n_216) );
OR2x2_ASAP7_75t_SL g217 ( .A(n_181), .B(n_140), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_190), .Y(n_218) );
AOI21x1_ASAP7_75t_L g219 ( .A1(n_175), .A2(n_154), .B(n_145), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_177), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_190), .Y(n_221) );
NAND2xp33_ASAP7_75t_L g222 ( .A(n_182), .B(n_137), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_182), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_182), .Y(n_225) );
INVx5_ASAP7_75t_L g226 ( .A(n_177), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_190), .Y(n_227) );
INVx3_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
OR2x2_ASAP7_75t_L g229 ( .A(n_178), .B(n_132), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_190), .Y(n_230) );
AND3x2_ASAP7_75t_L g231 ( .A(n_178), .B(n_172), .C(n_151), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_175), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_195), .B(n_149), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_181), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_176), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_208), .B(n_195), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_208), .B(n_181), .Y(n_238) );
NOR2xp33_ASAP7_75t_SL g239 ( .A(n_229), .B(n_148), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_229), .B(n_180), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_201), .B(n_181), .Y(n_241) );
INVxp67_ASAP7_75t_SL g242 ( .A(n_205), .Y(n_242) );
NAND2xp33_ASAP7_75t_L g243 ( .A(n_211), .B(n_193), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_201), .B(n_181), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_234), .B(n_186), .Y(n_246) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_202), .A2(n_197), .B(n_196), .C(n_188), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_205), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_205), .B(n_180), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_210), .B(n_189), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_228), .B(n_189), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_228), .B(n_189), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_232), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_228), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_216), .B(n_184), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_235), .B(n_184), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_206), .B(n_187), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_216), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_228), .B(n_187), .Y(n_260) );
NAND3xp33_ASAP7_75t_L g261 ( .A(n_231), .B(n_163), .C(n_164), .Y(n_261) );
NAND3xp33_ASAP7_75t_L g262 ( .A(n_210), .B(n_194), .C(n_192), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_225), .B(n_197), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_232), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_235), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_224), .B(n_197), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_233), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_233), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_202), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_225), .B(n_146), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_236), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_224), .B(n_185), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_203), .B(n_165), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_203), .B(n_165), .Y(n_274) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_222), .B(n_194), .C(n_192), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_223), .B(n_173), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_217), .B(n_188), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_198), .A2(n_173), .B1(n_170), .B2(n_150), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_223), .B(n_196), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_225), .B(n_147), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_225), .B(n_141), .Y(n_281) );
AND2x4_ASAP7_75t_SL g282 ( .A(n_217), .B(n_136), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_207), .B(n_155), .Y(n_283) );
AOI22xp5_ASAP7_75t_L g284 ( .A1(n_214), .A2(n_166), .B1(n_157), .B2(n_160), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_215), .B(n_143), .Y(n_285) );
NAND2xp33_ASAP7_75t_L g286 ( .A(n_236), .B(n_152), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_219), .B(n_191), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_219), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_226), .B(n_153), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_226), .B(n_169), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_226), .B(n_136), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g293 ( .A1(n_288), .A2(n_191), .B(n_192), .Y(n_293) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_256), .A2(n_161), .B1(n_156), .B2(n_159), .Y(n_294) );
INVx3_ASAP7_75t_L g295 ( .A(n_245), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_258), .B(n_171), .Y(n_296) );
O2A1O1Ixp5_ASAP7_75t_L g297 ( .A1(n_251), .A2(n_283), .B(n_270), .C(n_280), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_240), .B(n_162), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_257), .B(n_174), .Y(n_299) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_258), .B(n_136), .Y(n_300) );
NAND2xp5_ASAP7_75t_SL g301 ( .A(n_249), .B(n_134), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_249), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_245), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_251), .A2(n_192), .B(n_191), .Y(n_304) );
O2A1O1Ixp5_ASAP7_75t_L g305 ( .A1(n_283), .A2(n_212), .B(n_200), .C(n_209), .Y(n_305) );
O2A1O1Ixp33_ASAP7_75t_L g306 ( .A1(n_259), .A2(n_176), .B(n_191), .C(n_192), .Y(n_306) );
NOR2x1_ASAP7_75t_L g307 ( .A(n_261), .B(n_176), .Y(n_307) );
A2O1A1Ixp33_ASAP7_75t_L g308 ( .A1(n_262), .A2(n_179), .B(n_227), .C(n_199), .Y(n_308) );
BUFx2_ASAP7_75t_L g309 ( .A(n_258), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_257), .B(n_2), .Y(n_310) );
OAI21xp5_ASAP7_75t_L g311 ( .A1(n_287), .A2(n_213), .B(n_200), .Y(n_311) );
BUFx4f_ASAP7_75t_L g312 ( .A(n_282), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_237), .A2(n_213), .B(n_209), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_254), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_250), .B(n_5), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_249), .B(n_226), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_287), .A2(n_213), .B(n_200), .Y(n_318) );
AOI21x1_ASAP7_75t_L g319 ( .A1(n_270), .A2(n_209), .B(n_212), .Y(n_319) );
O2A1O1Ixp33_ASAP7_75t_L g320 ( .A1(n_247), .A2(n_212), .B(n_227), .C(n_221), .Y(n_320) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_275), .B(n_199), .Y(n_321) );
OAI321xp33_ASAP7_75t_L g322 ( .A1(n_241), .A2(n_179), .A3(n_221), .B1(n_218), .B2(n_204), .C(n_230), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_239), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g324 ( .A1(n_243), .A2(n_6), .B(n_7), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_249), .B(n_255), .Y(n_325) );
O2A1O1Ixp5_ASAP7_75t_L g326 ( .A1(n_280), .A2(n_230), .B(n_218), .C(n_204), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_260), .B(n_6), .Y(n_327) );
BUFx8_ASAP7_75t_L g328 ( .A(n_277), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_282), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_254), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_246), .B(n_7), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_252), .A2(n_220), .B(n_226), .Y(n_332) );
AOI21xp5_ASAP7_75t_L g333 ( .A1(n_253), .A2(n_220), .B(n_226), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_246), .B(n_8), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_264), .Y(n_335) );
NAND2xp5_ASAP7_75t_SL g336 ( .A(n_264), .B(n_179), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_267), .B(n_179), .Y(n_337) );
CKINVDCx11_ASAP7_75t_R g338 ( .A(n_267), .Y(n_338) );
NAND3xp33_ASAP7_75t_L g339 ( .A(n_243), .B(n_179), .C(n_220), .Y(n_339) );
INVx2_ASAP7_75t_SL g340 ( .A(n_312), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_309), .B(n_244), .Y(n_341) );
OAI21xp5_ASAP7_75t_L g342 ( .A1(n_304), .A2(n_242), .B(n_263), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_297), .A2(n_263), .B(n_266), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_312), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_308), .A2(n_247), .B(n_276), .Y(n_345) );
O2A1O1Ixp5_ASAP7_75t_L g346 ( .A1(n_301), .A2(n_290), .B(n_238), .C(n_274), .Y(n_346) );
AOI21xp5_ASAP7_75t_SL g347 ( .A1(n_306), .A2(n_279), .B(n_272), .Y(n_347) );
OAI21xp5_ASAP7_75t_L g348 ( .A1(n_321), .A2(n_273), .B(n_268), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_293), .A2(n_285), .B(n_281), .Y(n_351) );
AOI21xp5_ASAP7_75t_L g352 ( .A1(n_311), .A2(n_286), .B(n_290), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_318), .A2(n_286), .B(n_271), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_325), .A2(n_313), .B(n_292), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
INVx5_ASAP7_75t_L g356 ( .A(n_302), .Y(n_356) );
OAI21xp5_ASAP7_75t_L g357 ( .A1(n_327), .A2(n_271), .B(n_268), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_302), .B(n_284), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_334), .B(n_278), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_302), .B(n_265), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_320), .A2(n_289), .B(n_291), .Y(n_363) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_325), .A2(n_220), .B(n_179), .Y(n_364) );
AND3x4_ASAP7_75t_L g365 ( .A(n_307), .B(n_8), .C(n_10), .Y(n_365) );
HAxp5_ASAP7_75t_L g366 ( .A(n_328), .B(n_10), .CON(n_366), .SN(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_300), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_292), .A2(n_220), .B(n_60), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_330), .A2(n_58), .B(n_118), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_330), .A2(n_57), .B(n_117), .Y(n_370) );
OAI21x1_ASAP7_75t_SL g371 ( .A1(n_310), .A2(n_12), .B(n_13), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_319), .A2(n_63), .B(n_116), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_349), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_359), .Y(n_376) );
OR2x6_ASAP7_75t_L g377 ( .A(n_347), .B(n_302), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_359), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_347), .A2(n_301), .B(n_305), .Y(n_379) );
BUFx3_ASAP7_75t_L g380 ( .A(n_356), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_372), .A2(n_326), .B(n_333), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_372), .A2(n_332), .B(n_337), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_356), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_351), .A2(n_337), .B(n_336), .Y(n_384) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g386 ( .A(n_356), .B(n_316), .Y(n_386) );
OA21x2_ASAP7_75t_L g387 ( .A1(n_345), .A2(n_322), .B(n_339), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_373), .B(n_334), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_373), .Y(n_389) );
OAI21x1_ASAP7_75t_L g390 ( .A1(n_353), .A2(n_336), .B(n_316), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_331), .B(n_300), .Y(n_391) );
OAI21x1_ASAP7_75t_L g392 ( .A1(n_348), .A2(n_317), .B(n_295), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_369), .A2(n_295), .B(n_303), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_367), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_358), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_356), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_343), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_363), .A2(n_324), .B(n_296), .Y(n_398) );
OAI21x1_ASAP7_75t_L g399 ( .A1(n_352), .A2(n_299), .B(n_296), .Y(n_399) );
AO31x2_ASAP7_75t_L g400 ( .A1(n_361), .A2(n_298), .A3(n_15), .B(n_16), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_376), .Y(n_403) );
INVx3_ASAP7_75t_L g404 ( .A(n_380), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_378), .Y(n_405) );
BUFx2_ASAP7_75t_L g406 ( .A(n_374), .Y(n_406) );
OAI21x1_ASAP7_75t_L g407 ( .A1(n_393), .A2(n_368), .B(n_342), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_378), .B(n_366), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_389), .Y(n_410) );
AOI21x1_ASAP7_75t_L g411 ( .A1(n_377), .A2(n_360), .B(n_364), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_395), .A2(n_323), .B1(n_366), .B2(n_355), .C(n_294), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_377), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_391), .A2(n_346), .B(n_357), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_389), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_389), .Y(n_416) );
INVxp67_ASAP7_75t_L g417 ( .A(n_389), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_375), .Y(n_418) );
AOI21x1_ASAP7_75t_L g419 ( .A1(n_377), .A2(n_360), .B(n_370), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_375), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_375), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g422 ( .A1(n_399), .A2(n_397), .B(n_391), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
OR2x6_ASAP7_75t_L g424 ( .A(n_377), .B(n_362), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_394), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_385), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_380), .B(n_340), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_380), .Y(n_428) );
AOI21x1_ASAP7_75t_L g429 ( .A1(n_377), .A2(n_371), .B(n_341), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_394), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_392), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_380), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_395), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_392), .Y(n_435) );
BUFx2_ASAP7_75t_L g436 ( .A(n_406), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_425), .B(n_400), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_416), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_408), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_410), .B(n_396), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_409), .A2(n_365), .B1(n_388), .B2(n_338), .Y(n_442) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_409), .A2(n_383), .B1(n_385), .B2(n_396), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_410), .B(n_401), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_413), .B(n_377), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_413), .A2(n_365), .B1(n_388), .B2(n_398), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_415), .B(n_401), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_415), .B(n_401), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_417), .B(n_401), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_408), .B(n_400), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_417), .B(n_396), .Y(n_451) );
INVx2_ASAP7_75t_R g452 ( .A(n_418), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_406), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_425), .B(n_400), .Y(n_454) );
INVx4_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
NAND2x1_ASAP7_75t_L g456 ( .A(n_424), .B(n_418), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_426), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_423), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_423), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_430), .B(n_400), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_420), .B(n_430), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_402), .B(n_400), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
NOR2x1p5_ASAP7_75t_L g464 ( .A(n_404), .B(n_396), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_402), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_428), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_403), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_403), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_420), .B(n_388), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_421), .B(n_400), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_428), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_404), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_421), .B(n_400), .Y(n_474) );
BUFx2_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
BUFx3_ASAP7_75t_L g476 ( .A(n_404), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_421), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_433), .B(n_392), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_405), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_405), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_434), .B(n_400), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_434), .B(n_399), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_433), .B(n_391), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_427), .B(n_383), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_432), .B(n_399), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_432), .B(n_398), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_422), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_422), .A2(n_379), .B(n_393), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_471), .B(n_431), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_471), .B(n_431), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_465), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_474), .B(n_435), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_465), .Y(n_495) );
OAI21xp5_ASAP7_75t_SL g496 ( .A1(n_443), .A2(n_427), .B(n_432), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_467), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_474), .B(n_435), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_446), .A2(n_427), .B1(n_398), .B2(n_424), .Y(n_499) );
INVxp67_ASAP7_75t_SL g500 ( .A(n_439), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_477), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_481), .B(n_435), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_436), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_467), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_469), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_481), .B(n_482), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_470), .B(n_432), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_469), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_479), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_482), .B(n_414), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_479), .Y(n_511) );
AOI211x1_ASAP7_75t_L g512 ( .A1(n_437), .A2(n_429), .B(n_412), .C(n_411), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_470), .B(n_427), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_461), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_461), .Y(n_515) );
BUFx3_ASAP7_75t_L g516 ( .A(n_436), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_438), .B(n_424), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_477), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_438), .B(n_424), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_458), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_449), .B(n_414), .Y(n_521) );
BUFx2_ASAP7_75t_L g522 ( .A(n_453), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_442), .A2(n_398), .B1(n_414), .B2(n_385), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_449), .B(n_414), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_480), .B(n_398), .Y(n_525) );
BUFx2_ASAP7_75t_L g526 ( .A(n_453), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_455), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_475), .A2(n_414), .B1(n_350), .B2(n_387), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_451), .B(n_429), .Y(n_529) );
INVx3_ASAP7_75t_L g530 ( .A(n_455), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_441), .B(n_14), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_441), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_477), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_451), .B(n_411), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_444), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_444), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_447), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_447), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_437), .B(n_412), .C(n_387), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_448), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_458), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_459), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_453), .A2(n_344), .B1(n_386), .B2(n_387), .Y(n_543) );
AND2x4_ASAP7_75t_L g544 ( .A(n_445), .B(n_419), .Y(n_544) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_438), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_453), .A2(n_386), .B1(n_344), .B2(n_362), .Y(n_546) );
BUFx2_ASAP7_75t_L g547 ( .A(n_440), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_448), .B(n_379), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_484), .Y(n_549) );
AND2x4_ASAP7_75t_L g550 ( .A(n_445), .B(n_419), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_459), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_486), .B(n_379), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_463), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_486), .B(n_407), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_440), .B(n_407), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_440), .B(n_407), .Y(n_556) );
AND2x4_ASAP7_75t_L g557 ( .A(n_445), .B(n_390), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_463), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_483), .B(n_390), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_460), .B(n_14), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_483), .B(n_390), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_462), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_484), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_445), .B(n_382), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_484), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_483), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_483), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_464), .A2(n_386), .B1(n_387), .B2(n_19), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_462), .Y(n_569) );
INVxp67_ASAP7_75t_L g570 ( .A(n_468), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_488), .B(n_387), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_455), .B(n_386), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_514), .B(n_460), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_493), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_506), .B(n_450), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_506), .B(n_478), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_493), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_549), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_514), .B(n_454), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_495), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_522), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_500), .B(n_450), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_495), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_522), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_502), .B(n_478), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_497), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_502), .B(n_478), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_563), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_532), .B(n_466), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_515), .B(n_466), .Y(n_591) );
BUFx3_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_529), .B(n_478), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_535), .B(n_472), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_547), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_529), .B(n_491), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_491), .B(n_488), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_497), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_492), .B(n_487), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_492), .B(n_494), .Y(n_600) );
AND2x4_ASAP7_75t_SL g601 ( .A(n_527), .B(n_455), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_526), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_512), .A2(n_457), .B1(n_454), .B2(n_487), .C(n_475), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_504), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_494), .B(n_452), .Y(n_605) );
BUFx2_ASAP7_75t_SL g606 ( .A(n_527), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_498), .B(n_452), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_527), .B(n_489), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_498), .B(n_452), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_547), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_504), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_515), .B(n_472), .Y(n_612) );
BUFx2_ASAP7_75t_SL g613 ( .A(n_530), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_536), .B(n_476), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_537), .B(n_464), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_505), .Y(n_616) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_530), .B(n_456), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_538), .B(n_456), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_505), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_508), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_508), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_540), .B(n_485), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_562), .B(n_473), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_563), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_513), .B(n_476), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_570), .B(n_476), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_507), .B(n_473), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_503), .B(n_489), .Y(n_628) );
HB1xp67_ASAP7_75t_SL g629 ( .A(n_516), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_562), .B(n_489), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_530), .Y(n_631) );
NOR2x1p5_ASAP7_75t_L g632 ( .A(n_516), .B(n_489), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_560), .B(n_489), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_523), .A2(n_393), .B(n_382), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_566), .B(n_489), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_510), .B(n_490), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_509), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_509), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_511), .B(n_490), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_569), .B(n_490), .Y(n_640) );
INVxp33_ASAP7_75t_L g641 ( .A(n_496), .Y(n_641) );
AND2x2_ASAP7_75t_L g642 ( .A(n_569), .B(n_490), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_545), .B(n_17), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_517), .B(n_18), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_521), .B(n_18), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_566), .B(n_382), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_511), .B(n_20), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_565), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_572), .A2(n_384), .B(n_381), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_520), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_510), .B(n_384), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_520), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_565), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_541), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_501), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_521), .B(n_20), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_567), .B(n_381), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_541), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_501), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_518), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_552), .B(n_384), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_524), .B(n_21), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_524), .B(n_22), .Y(n_663) );
AND2x2_ASAP7_75t_L g664 ( .A(n_552), .B(n_381), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_567), .B(n_22), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_542), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_542), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_534), .B(n_23), .Y(n_668) );
AND2x4_ASAP7_75t_SL g669 ( .A(n_600), .B(n_553), .Y(n_669) );
OAI21xp5_ASAP7_75t_L g670 ( .A1(n_641), .A2(n_539), .B(n_568), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_574), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_577), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_580), .Y(n_673) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_595), .Y(n_674) );
AND2x4_ASAP7_75t_L g675 ( .A(n_601), .B(n_544), .Y(n_675) );
INVx3_ASAP7_75t_L g676 ( .A(n_601), .Y(n_676) );
OR2x2_ASAP7_75t_L g677 ( .A(n_575), .B(n_517), .Y(n_677) );
AND2x4_ASAP7_75t_L g678 ( .A(n_592), .B(n_544), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_583), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_600), .B(n_559), .Y(n_680) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_631), .B(n_544), .Y(n_681) );
OAI21xp33_ASAP7_75t_SL g682 ( .A1(n_632), .A2(n_543), .B(n_499), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_596), .B(n_519), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_596), .B(n_559), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_576), .B(n_561), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_587), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_598), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_636), .B(n_525), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_604), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_636), .B(n_551), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_576), .B(n_561), .Y(n_691) );
INVxp33_ASAP7_75t_L g692 ( .A(n_629), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_611), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_585), .B(n_557), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_582), .B(n_519), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_595), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_616), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_655), .Y(n_698) );
NOR2x1_ASAP7_75t_L g699 ( .A(n_606), .B(n_546), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_592), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_619), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_599), .B(n_534), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_597), .B(n_551), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_585), .B(n_557), .Y(n_704) );
NOR2xp67_ASAP7_75t_SL g705 ( .A(n_613), .B(n_531), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_588), .B(n_557), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_620), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_637), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_655), .Y(n_710) );
OR2x2_ASAP7_75t_L g711 ( .A(n_599), .B(n_548), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_597), .B(n_558), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_638), .Y(n_713) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_610), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_573), .B(n_558), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_622), .B(n_579), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_610), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_650), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_660), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_652), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_660), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_654), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_658), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_666), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_581), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_581), .B(n_548), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_667), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_588), .B(n_593), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_593), .B(n_564), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_623), .Y(n_730) );
OR2x6_ASAP7_75t_L g731 ( .A(n_617), .B(n_550), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_590), .Y(n_732) );
OR2x2_ASAP7_75t_L g733 ( .A(n_602), .B(n_554), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_641), .A2(n_528), .B1(n_518), .B2(n_533), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_625), .B(n_564), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_594), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_615), .Y(n_737) );
INVx4_ASAP7_75t_L g738 ( .A(n_617), .Y(n_738) );
NOR4xp75_ASAP7_75t_L g739 ( .A(n_656), .B(n_554), .C(n_556), .D(n_555), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_627), .B(n_564), .Y(n_740) );
AND2x4_ASAP7_75t_SL g741 ( .A(n_614), .B(n_533), .Y(n_741) );
OR2x2_ASAP7_75t_L g742 ( .A(n_602), .B(n_556), .Y(n_742) );
OR2x2_ASAP7_75t_L g743 ( .A(n_630), .B(n_555), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_584), .B(n_571), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_591), .Y(n_745) );
AND2x2_ASAP7_75t_L g746 ( .A(n_626), .B(n_550), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_628), .B(n_550), .Y(n_747) );
OAI222xp33_ASAP7_75t_L g748 ( .A1(n_584), .A2(n_571), .B1(n_27), .B2(n_28), .C1(n_29), .C2(n_31), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_605), .B(n_26), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_605), .B(n_32), .Y(n_750) );
OR2x2_ASAP7_75t_L g751 ( .A(n_651), .B(n_34), .Y(n_751) );
NOR2xp67_ASAP7_75t_L g752 ( .A(n_631), .B(n_36), .Y(n_752) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_607), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_645), .A2(n_38), .B1(n_39), .B2(n_40), .Y(n_754) );
NOR2x1p5_ASAP7_75t_L g755 ( .A(n_643), .B(n_41), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_669), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_692), .B(n_662), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_703), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_703), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_682), .A2(n_603), .B1(n_663), .B2(n_651), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_712), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_741), .Y(n_762) );
OAI31xp33_ASAP7_75t_L g763 ( .A1(n_755), .A2(n_644), .A3(n_668), .B(n_618), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g764 ( .A1(n_738), .A2(n_668), .B1(n_633), .B2(n_647), .Y(n_764) );
INVxp67_ASAP7_75t_L g765 ( .A(n_696), .Y(n_765) );
AND2x2_ASAP7_75t_SL g766 ( .A(n_738), .B(n_608), .Y(n_766) );
INVx2_ASAP7_75t_L g767 ( .A(n_698), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_688), .B(n_690), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_688), .B(n_639), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_712), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_671), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_672), .Y(n_772) );
AND2x4_ASAP7_75t_L g773 ( .A(n_681), .B(n_608), .Y(n_773) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_674), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_737), .B(n_612), .Y(n_775) );
AOI321xp33_ASAP7_75t_L g776 ( .A1(n_734), .A2(n_664), .A3(n_665), .B1(n_661), .B2(n_607), .C(n_609), .Y(n_776) );
AOI32xp33_ASAP7_75t_L g777 ( .A1(n_699), .A2(n_609), .A3(n_608), .B1(n_661), .B2(n_640), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_673), .Y(n_778) );
OAI21xp33_ASAP7_75t_L g779 ( .A1(n_682), .A2(n_642), .B(n_664), .Y(n_779) );
AND2x2_ASAP7_75t_L g780 ( .A(n_685), .B(n_635), .Y(n_780) );
NAND4xp75_ASAP7_75t_L g781 ( .A(n_670), .B(n_634), .C(n_649), .D(n_653), .Y(n_781) );
NAND2xp5_ASAP7_75t_SL g782 ( .A(n_676), .B(n_635), .Y(n_782) );
XOR2x2_ASAP7_75t_L g783 ( .A(n_739), .B(n_635), .Y(n_783) );
O2A1O1Ixp33_ASAP7_75t_L g784 ( .A1(n_670), .A2(n_659), .B(n_586), .C(n_653), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_734), .A2(n_646), .B1(n_657), .B2(n_648), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_710), .Y(n_786) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_676), .A2(n_659), .B1(n_578), .B2(n_648), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_679), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_686), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_687), .Y(n_790) );
HB1xp67_ASAP7_75t_L g791 ( .A(n_717), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_689), .Y(n_792) );
OAI22xp33_ASAP7_75t_SL g793 ( .A1(n_731), .A2(n_624), .B1(n_589), .B2(n_586), .Y(n_793) );
HB1xp67_ASAP7_75t_L g794 ( .A(n_714), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_674), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_719), .Y(n_796) );
OR2x2_ASAP7_75t_L g797 ( .A(n_690), .B(n_624), .Y(n_797) );
INVx2_ASAP7_75t_SL g798 ( .A(n_700), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_693), .Y(n_799) );
NAND2x1_ASAP7_75t_L g800 ( .A(n_731), .B(n_589), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_721), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_697), .Y(n_802) );
NOR3xp33_ASAP7_75t_L g803 ( .A(n_748), .B(n_578), .C(n_657), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_705), .A2(n_646), .B1(n_657), .B2(n_45), .Y(n_804) );
AND2x2_ASAP7_75t_L g805 ( .A(n_691), .B(n_646), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_701), .Y(n_806) );
OR2x2_ASAP7_75t_L g807 ( .A(n_702), .B(n_43), .Y(n_807) );
NOR2xp67_ASAP7_75t_SL g808 ( .A(n_751), .B(n_44), .Y(n_808) );
INVx2_ASAP7_75t_L g809 ( .A(n_742), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_743), .Y(n_810) );
XOR2x2_ASAP7_75t_L g811 ( .A(n_752), .B(n_46), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_707), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_708), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_709), .Y(n_814) );
AOI21xp5_ASAP7_75t_L g815 ( .A1(n_800), .A2(n_731), .B(n_681), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g816 ( .A1(n_762), .A2(n_675), .B1(n_753), .B2(n_711), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_760), .B(n_730), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g818 ( .A1(n_762), .A2(n_675), .B1(n_716), .B2(n_683), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_758), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_779), .A2(n_736), .B1(n_732), .B2(n_745), .Y(n_820) );
OAI221xp5_ASAP7_75t_L g821 ( .A1(n_777), .A2(n_725), .B1(n_715), .B2(n_733), .C(n_754), .Y(n_821) );
NOR2x1_ASAP7_75t_L g822 ( .A(n_781), .B(n_752), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_803), .A2(n_746), .B1(n_678), .B2(n_747), .Y(n_823) );
O2A1O1Ixp33_ASAP7_75t_L g824 ( .A1(n_795), .A2(n_748), .B(n_715), .C(n_749), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_759), .Y(n_825) );
INVx1_ASAP7_75t_SL g826 ( .A(n_794), .Y(n_826) );
INVx1_ASAP7_75t_L g827 ( .A(n_761), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g828 ( .A(n_776), .B(n_754), .C(n_750), .Y(n_828) );
AOI21xp33_ASAP7_75t_SL g829 ( .A1(n_766), .A2(n_678), .B(n_726), .Y(n_829) );
INVx1_ASAP7_75t_SL g830 ( .A(n_798), .Y(n_830) );
OAI222xp33_ASAP7_75t_L g831 ( .A1(n_785), .A2(n_744), .B1(n_677), .B2(n_695), .C1(n_729), .C2(n_706), .Y(n_831) );
XOR2x2_ASAP7_75t_L g832 ( .A(n_811), .B(n_728), .Y(n_832) );
O2A1O1Ixp33_ASAP7_75t_L g833 ( .A1(n_795), .A2(n_720), .B(n_718), .C(n_727), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_791), .Y(n_834) );
XOR2x2_ASAP7_75t_L g835 ( .A(n_757), .B(n_680), .Y(n_835) );
INVx2_ASAP7_75t_SL g836 ( .A(n_756), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_770), .Y(n_837) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_803), .A2(n_694), .B1(n_704), .B2(n_684), .Y(n_838) );
OAI321xp33_ASAP7_75t_L g839 ( .A1(n_776), .A2(n_724), .A3(n_723), .B1(n_722), .B2(n_713), .C(n_735), .Y(n_839) );
OAI22xp33_ASAP7_75t_SL g840 ( .A1(n_774), .A2(n_740), .B1(n_50), .B2(n_51), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_768), .B(n_48), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_771), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_765), .B(n_54), .Y(n_843) );
OAI21xp33_ASAP7_75t_L g844 ( .A1(n_769), .A2(n_55), .B(n_64), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_772), .Y(n_845) );
NAND2x1_ASAP7_75t_L g846 ( .A(n_773), .B(n_65), .Y(n_846) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_783), .A2(n_66), .B1(n_67), .B2(n_68), .Y(n_847) );
AOI222xp33_ASAP7_75t_L g848 ( .A1(n_774), .A2(n_70), .B1(n_72), .B2(n_75), .C1(n_76), .C2(n_78), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_838), .A2(n_764), .B1(n_782), .B2(n_775), .Y(n_849) );
O2A1O1Ixp5_ASAP7_75t_L g850 ( .A1(n_817), .A2(n_787), .B(n_769), .C(n_812), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_819), .B(n_778), .Y(n_851) );
OAI21xp33_ASAP7_75t_L g852 ( .A1(n_823), .A2(n_793), .B(n_765), .Y(n_852) );
NAND4xp25_ASAP7_75t_L g853 ( .A(n_824), .B(n_763), .C(n_804), .D(n_784), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_826), .Y(n_854) );
NAND4xp25_ASAP7_75t_L g855 ( .A(n_822), .B(n_763), .C(n_784), .D(n_807), .Y(n_855) );
INVx2_ASAP7_75t_SL g856 ( .A(n_830), .Y(n_856) );
AOI21xp5_ASAP7_75t_L g857 ( .A1(n_839), .A2(n_791), .B(n_773), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_826), .Y(n_858) );
AOI22x1_ASAP7_75t_L g859 ( .A1(n_815), .A2(n_809), .B1(n_810), .B2(n_797), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_829), .B(n_796), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_842), .Y(n_861) );
NAND2xp5_ASAP7_75t_SL g862 ( .A(n_820), .B(n_840), .Y(n_862) );
OAI221xp5_ASAP7_75t_L g863 ( .A1(n_821), .A2(n_814), .B1(n_813), .B2(n_788), .C(n_806), .Y(n_863) );
OAI31xp33_ASAP7_75t_L g864 ( .A1(n_828), .A2(n_792), .A3(n_802), .B(n_799), .Y(n_864) );
AOI211xp5_ASAP7_75t_L g865 ( .A1(n_828), .A2(n_808), .B(n_789), .C(n_790), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_818), .A2(n_801), .B(n_786), .Y(n_866) );
AOI221xp5_ASAP7_75t_L g867 ( .A1(n_831), .A2(n_767), .B1(n_805), .B2(n_780), .C(n_86), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g868 ( .A1(n_864), .A2(n_816), .B1(n_833), .B2(n_836), .C(n_827), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g869 ( .A(n_856), .B(n_825), .Y(n_869) );
NAND2xp5_ASAP7_75t_SL g870 ( .A(n_859), .B(n_834), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_854), .B(n_837), .Y(n_871) );
NAND3xp33_ASAP7_75t_L g872 ( .A(n_865), .B(n_850), .C(n_858), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_851), .Y(n_873) );
INVx1_ASAP7_75t_L g874 ( .A(n_851), .Y(n_874) );
NAND2xp5_ASAP7_75t_SL g875 ( .A(n_867), .B(n_847), .Y(n_875) );
AOI222xp33_ASAP7_75t_L g876 ( .A1(n_862), .A2(n_832), .B1(n_835), .B2(n_845), .C1(n_841), .C2(n_843), .Y(n_876) );
AOI21xp5_ASAP7_75t_L g877 ( .A1(n_860), .A2(n_846), .B(n_848), .Y(n_877) );
NOR3xp33_ASAP7_75t_L g878 ( .A(n_872), .B(n_853), .C(n_855), .Y(n_878) );
NAND5xp2_ASAP7_75t_L g879 ( .A(n_876), .B(n_857), .C(n_863), .D(n_852), .E(n_849), .Y(n_879) );
INVxp67_ASAP7_75t_L g880 ( .A(n_869), .Y(n_880) );
NAND4xp25_ASAP7_75t_L g881 ( .A(n_877), .B(n_866), .C(n_844), .D(n_861), .Y(n_881) );
NAND3xp33_ASAP7_75t_SL g882 ( .A(n_868), .B(n_80), .C(n_82), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_873), .B(n_83), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_878), .B(n_874), .Y(n_884) );
NAND3xp33_ASAP7_75t_L g885 ( .A(n_880), .B(n_870), .C(n_875), .Y(n_885) );
NAND4xp25_ASAP7_75t_L g886 ( .A(n_879), .B(n_871), .C(n_89), .D(n_92), .Y(n_886) );
NOR3xp33_ASAP7_75t_L g887 ( .A(n_882), .B(n_87), .C(n_94), .Y(n_887) );
NAND4xp75_ASAP7_75t_L g888 ( .A(n_884), .B(n_883), .C(n_881), .D(n_99), .Y(n_888) );
INVx1_ASAP7_75t_SL g889 ( .A(n_885), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_886), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_889), .B(n_887), .Y(n_891) );
INVx1_ASAP7_75t_L g892 ( .A(n_890), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_892), .Y(n_893) );
AO21x1_ASAP7_75t_L g894 ( .A1(n_891), .A2(n_888), .B(n_97), .Y(n_894) );
XNOR2xp5_ASAP7_75t_SL g895 ( .A(n_893), .B(n_891), .Y(n_895) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_894), .A2(n_96), .B(n_101), .Y(n_896) );
AOI21xp5_ASAP7_75t_L g897 ( .A1(n_896), .A2(n_102), .B(n_107), .Y(n_897) );
AOI21x1_ASAP7_75t_L g898 ( .A1(n_897), .A2(n_895), .B(n_111), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_898), .A2(n_109), .B(n_112), .Y(n_899) );
INVx1_ASAP7_75t_L g900 ( .A(n_899), .Y(n_900) );
UNKNOWN g901 ( );
OAI21xp33_ASAP7_75t_L g902 ( .A1(n_901), .A2(n_114), .B(n_121), .Y(n_902) );
endmodule