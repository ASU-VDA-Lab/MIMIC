module fake_netlist_6_2494_n_110 (n_16, n_1, n_9, n_8, n_18, n_10, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_7, n_2, n_5, n_19, n_110);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_7;
input n_2;
input n_5;
input n_19;

output n_110;

wire n_52;
wire n_91;
wire n_46;
wire n_21;
wire n_88;
wire n_98;
wire n_39;
wire n_63;
wire n_73;
wire n_22;
wire n_68;
wire n_28;
wire n_50;
wire n_49;
wire n_83;
wire n_101;
wire n_77;
wire n_106;
wire n_92;
wire n_42;
wire n_96;
wire n_90;
wire n_24;
wire n_105;
wire n_54;
wire n_102;
wire n_87;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_100;
wire n_23;
wire n_20;
wire n_47;
wire n_62;
wire n_29;
wire n_75;
wire n_109;
wire n_45;
wire n_34;
wire n_70;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_27;
wire n_38;
wire n_61;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_26;
wire n_55;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_64;
wire n_48;
wire n_65;
wire n_25;
wire n_40;
wire n_93;
wire n_80;
wire n_41;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_72;
wire n_89;
wire n_103;
wire n_60;
wire n_35;
wire n_69;
wire n_30;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_48),
.B1(n_34),
.B2(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_31),
.Y(n_56)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_24),
.B1(n_33),
.B2(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_37),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_47),
.Y(n_60)
);

CKINVDCx11_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_38),
.B1(n_39),
.B2(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_45),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_40),
.Y(n_65)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_48),
.B(n_54),
.C(n_46),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_57),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_57),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_35),
.B(n_30),
.C(n_29),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_62),
.Y(n_71)
);

OAI21x1_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_60),
.B(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

OAI21x1_ASAP7_75t_SL g74 ( 
.A1(n_66),
.A2(n_60),
.B(n_30),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_68),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_69),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_74),
.A2(n_62),
.B(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_77),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_78),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_56),
.Y(n_88)
);

AOI222xp33_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_31),
.B1(n_61),
.B2(n_58),
.C1(n_57),
.C2(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_85),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_83),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_83),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_93),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_86),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_82),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_87),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_97),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_101),
.A2(n_98),
.A3(n_99),
.B1(n_100),
.B2(n_89),
.C1(n_4),
.C2(n_7),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_87),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_103),
.B(n_87),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_105),
.C(n_104),
.Y(n_107)
);

OAI322xp33_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_106),
.A3(n_6),
.B1(n_81),
.B2(n_70),
.C1(n_18),
.C2(n_11),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_6),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_109),
.Y(n_110)
);


endmodule