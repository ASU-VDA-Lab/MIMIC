module fake_jpeg_28278_n_223 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_223);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_223;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_42),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_32),
.Y(n_58)
);

AND2x2_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_20),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_23),
.B1(n_31),
.B2(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_58),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_19),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_34),
.A2(n_28),
.B1(n_22),
.B2(n_19),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_61),
.B1(n_30),
.B2(n_18),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_21),
.B(n_32),
.C(n_29),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_60),
.A2(n_63),
.B(n_19),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_28),
.B1(n_29),
.B2(n_24),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g63 ( 
.A(n_33),
.B(n_26),
.CON(n_63),
.SN(n_63)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_38),
.B1(n_37),
.B2(n_34),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_65),
.A2(n_48),
.B1(n_46),
.B2(n_55),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_76),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_38),
.B1(n_27),
.B2(n_19),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_44),
.B1(n_47),
.B2(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_83),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_54),
.Y(n_105)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_79),
.Y(n_94)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_80),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_35),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_68),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_106),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_39),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_44),
.C(n_56),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_98),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_99),
.B(n_77),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_107),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_52),
.B1(n_57),
.B2(n_55),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_102),
.A2(n_105),
.B1(n_50),
.B2(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_54),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_74),
.A2(n_56),
.B1(n_50),
.B2(n_46),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_107),
.A2(n_65),
.B1(n_46),
.B2(n_48),
.Y(n_119)
);

BUFx24_ASAP7_75t_SL g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_121),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_125),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_100),
.B1(n_97),
.B2(n_81),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_64),
.B(n_60),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_128),
.B(n_88),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_50),
.B1(n_65),
.B2(n_80),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_117),
.A2(n_123),
.B1(n_98),
.B2(n_86),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_120),
.B1(n_126),
.B2(n_96),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_65),
.B1(n_70),
.B2(n_73),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_78),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_122),
.B(n_101),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_18),
.B1(n_39),
.B2(n_42),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_81),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_124),
.B(n_42),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_82),
.B(n_72),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g127 ( 
.A1(n_101),
.A2(n_82),
.B(n_72),
.C(n_35),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_16),
.B(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_139),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_118),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_93),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_135),
.B(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_149),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_122),
.B1(n_126),
.B2(n_125),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_138),
.B1(n_145),
.B2(n_117),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_101),
.B1(n_88),
.B2(n_97),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_143),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_104),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_114),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_146),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_25),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_163),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_116),
.C(n_112),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_154),
.C(n_162),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_116),
.C(n_126),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_146),
.A2(n_123),
.B1(n_128),
.B2(n_116),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_100),
.B1(n_72),
.B2(n_81),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_160),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_144),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_152),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_72),
.C(n_108),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_14),
.Y(n_165)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_171),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_141),
.A3(n_137),
.B1(n_135),
.B2(n_145),
.C1(n_136),
.C2(n_149),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_169),
.B(n_172),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_167),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_177),
.C(n_164),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_175),
.B(n_1),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_134),
.C(n_108),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_25),
.B1(n_14),
.B2(n_12),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_182),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_155),
.B(n_166),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_184),
.A2(n_171),
.B(n_176),
.Y(n_199)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_189),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_164),
.C(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_191),
.Y(n_196)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_16),
.C(n_2),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_178),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_172),
.B(n_178),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_194),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_197),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_193),
.B1(n_173),
.B2(n_188),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_202),
.A3(n_185),
.B1(n_184),
.B2(n_182),
.C1(n_176),
.C2(n_179),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_200),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_192),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_186),
.C(n_189),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

O2A1O1Ixp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_180),
.B(n_16),
.C(n_4),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_16),
.C(n_3),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_1),
.B(n_4),
.Y(n_214)
);

AOI221xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_204),
.B1(n_201),
.B2(n_202),
.C(n_209),
.Y(n_210)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_210),
.A2(n_213),
.B(n_214),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_196),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_207),
.B(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_211),
.A2(n_6),
.B(n_7),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_217),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_216),
.C(n_8),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g221 ( 
.A(n_220),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_219),
.C(n_6),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_10),
.Y(n_223)
);


endmodule