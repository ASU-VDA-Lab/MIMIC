module fake_ariane_2993_n_1428 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_372, n_377, n_15, n_23, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_357, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_359, n_155, n_127, n_1428);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_359;
input n_155;
input n_127;

output n_1428;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_520;
wire n_870;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_261),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_169),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_271),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_276),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_75),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_56),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_27),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_96),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_250),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_155),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_41),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_179),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_46),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_42),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_222),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_368),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_293),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_159),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_246),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_26),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_100),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_259),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_163),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_187),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_108),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_134),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_60),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_83),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_270),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_226),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_348),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_269),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_341),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_135),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_150),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_316),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_212),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_205),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_272),
.Y(n_421)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_52),
.B(n_171),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_60),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_166),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_24),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_14),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_195),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_310),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_20),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_40),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_115),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_170),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_153),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_257),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_370),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_311),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_216),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_277),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_9),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_308),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_149),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_130),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_176),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_214),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_114),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_238),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_227),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_274),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_138),
.Y(n_451)
);

BUFx5_ASAP7_75t_L g452 ( 
.A(n_93),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_55),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_26),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_113),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_373),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_128),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_157),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_192),
.Y(n_459)
);

CKINVDCx14_ASAP7_75t_R g460 ( 
.A(n_283),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_137),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_175),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_89),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_129),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_320),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_262),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_142),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_210),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_13),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_80),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_224),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_297),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_312),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_352),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_353),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_14),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_204),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_42),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_339),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_19),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_304),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_67),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_35),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_229),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_190),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_321),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_267),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_206),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_295),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_333),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_172),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_337),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_305),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_56),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_288),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_263),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_349),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_248),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_38),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_5),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_1),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_313),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_240),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_2),
.Y(n_504)
);

INVx2_ASAP7_75t_SL g505 ( 
.A(n_141),
.Y(n_505)
);

BUFx8_ASAP7_75t_SL g506 ( 
.A(n_95),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_69),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_29),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_239),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_196),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_53),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_291),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_17),
.B(n_44),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_54),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_275),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_25),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_37),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_110),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_328),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_292),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_282),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_294),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_203),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_290),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_285),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_256),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_343),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_98),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_139),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_254),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_178),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_231),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_234),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_3),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_245),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_217),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_88),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_64),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_64),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_174),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_165),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_243),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_350),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_110),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_19),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_152),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_318),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_322),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_252),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_247),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_258),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_249),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_29),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_286),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_364),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_335),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_72),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_363),
.Y(n_558)
);

INVxp33_ASAP7_75t_SL g559 ( 
.A(n_177),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_452),
.B(n_0),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_383),
.B(n_0),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_452),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_428),
.B(n_1),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_511),
.B(n_2),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_428),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_407),
.B(n_3),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_452),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_414),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_414),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_469),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_423),
.B(n_4),
.Y(n_571)
);

CKINVDCx6p67_ASAP7_75t_R g572 ( 
.A(n_384),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_414),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_406),
.B(n_4),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_539),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_414),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_475),
.B(n_5),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_442),
.B(n_6),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_452),
.Y(n_579)
);

NAND2x1_ASAP7_75t_L g580 ( 
.A(n_488),
.B(n_6),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_452),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_454),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_452),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_411),
.Y(n_584)
);

NOR2x1_ASAP7_75t_L g585 ( 
.A(n_411),
.B(n_127),
.Y(n_585)
);

XNOR2x2_ASAP7_75t_L g586 ( 
.A(n_386),
.B(n_513),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_387),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_491),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_384),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_460),
.B(n_7),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_388),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_391),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_393),
.Y(n_593)
);

OA21x2_ASAP7_75t_L g594 ( 
.A1(n_381),
.A2(n_7),
.B(n_8),
.Y(n_594)
);

BUFx8_ASAP7_75t_L g595 ( 
.A(n_380),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_449),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

OA21x2_ASAP7_75t_L g598 ( 
.A1(n_382),
.A2(n_8),
.B(n_9),
.Y(n_598)
);

BUFx8_ASAP7_75t_L g599 ( 
.A(n_505),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_394),
.Y(n_600)
);

BUFx12f_ASAP7_75t_L g601 ( 
.A(n_412),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_449),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_401),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_390),
.B(n_10),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_554),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_395),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_489),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_10),
.Y(n_608)
);

BUFx12f_ASAP7_75t_L g609 ( 
.A(n_412),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_399),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_402),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_490),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_405),
.Y(n_615)
);

XNOR2x2_ASAP7_75t_L g616 ( 
.A(n_409),
.B(n_11),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_506),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_466),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_466),
.Y(n_619)
);

OAI21x1_ASAP7_75t_L g620 ( 
.A1(n_398),
.A2(n_132),
.B(n_131),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_499),
.B(n_432),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_466),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_447),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_389),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_470),
.B(n_11),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_466),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_416),
.Y(n_629)
);

BUFx2_ASAP7_75t_L g630 ( 
.A(n_441),
.Y(n_630)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_441),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_417),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_418),
.B(n_12),
.Y(n_633)
);

AND2x6_ASAP7_75t_L g634 ( 
.A(n_486),
.B(n_133),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_419),
.Y(n_635)
);

INVx5_ASAP7_75t_L g636 ( 
.A(n_486),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_517),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_476),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_486),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_465),
.A2(n_140),
.B(n_136),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_478),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_455),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_522),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_611),
.B(n_555),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_590),
.B(n_559),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_617),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_608),
.B(n_444),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_576),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_568),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_568),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_611),
.Y(n_652)
);

INVx8_ASAP7_75t_L g653 ( 
.A(n_634),
.Y(n_653)
);

CKINVDCx16_ASAP7_75t_R g654 ( 
.A(n_617),
.Y(n_654)
);

INVx8_ASAP7_75t_L g655 ( 
.A(n_634),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_576),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

CKINVDCx6p67_ASAP7_75t_R g658 ( 
.A(n_572),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_573),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_579),
.Y(n_660)
);

NAND3xp33_ASAP7_75t_L g661 ( 
.A(n_643),
.B(n_637),
.C(n_561),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_573),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_573),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_583),
.A2(n_421),
.B(n_420),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_625),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_566),
.B(n_444),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_614),
.B(n_461),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_587),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_596),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_596),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_596),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_602),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_591),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_566),
.B(n_422),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_628),
.Y(n_675)
);

NOR2x1p5_ASAP7_75t_L g676 ( 
.A(n_614),
.B(n_455),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_602),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_628),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_571),
.B(n_468),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_592),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_643),
.A2(n_517),
.B1(n_385),
.B2(n_424),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_571),
.A2(n_577),
.B1(n_570),
.B2(n_630),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_593),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_607),
.B(n_461),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_564),
.B(n_547),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_607),
.B(n_595),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_561),
.B(n_558),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_626),
.B(n_563),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_613),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_613),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_626),
.B(n_379),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_668),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_687),
.A2(n_586),
.B1(n_578),
.B2(n_574),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_667),
.B(n_589),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_673),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_649),
.B(n_595),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_653),
.B(n_604),
.Y(n_697)
);

INVxp67_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_649),
.B(n_599),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_645),
.B(n_652),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_653),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_656),
.B(n_599),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_666),
.A2(n_560),
.B(n_633),
.C(n_604),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_656),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_L g705 ( 
.A1(n_661),
.A2(n_578),
.B1(n_631),
.B2(n_637),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_676),
.B(n_622),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_654),
.B(n_575),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_680),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_675),
.B(n_584),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_675),
.B(n_584),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_677),
.Y(n_711)
);

NAND2xp33_ASAP7_75t_L g712 ( 
.A(n_653),
.B(n_633),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_683),
.Y(n_713)
);

NOR2xp67_ASAP7_75t_L g714 ( 
.A(n_657),
.B(n_569),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_650),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_650),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_684),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_651),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_660),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_678),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_678),
.B(n_588),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_664),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_682),
.B(n_601),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_646),
.B(n_609),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_679),
.B(n_597),
.Y(n_726)
);

NAND3xp33_ASAP7_75t_L g727 ( 
.A(n_687),
.B(n_560),
.C(n_594),
.Y(n_727)
);

AND2x6_ASAP7_75t_L g728 ( 
.A(n_653),
.B(n_585),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_686),
.B(n_622),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_666),
.A2(n_631),
.B1(n_396),
.B2(n_403),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_646),
.B(n_621),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_R g732 ( 
.A(n_658),
.B(n_625),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_691),
.B(n_648),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_681),
.B(n_580),
.C(n_501),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_677),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_685),
.B(n_648),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_665),
.B(n_575),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_688),
.B(n_605),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_688),
.B(n_408),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_677),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_674),
.B(n_605),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_674),
.B(n_565),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_655),
.B(n_562),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_659),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_655),
.B(n_606),
.Y(n_745)
);

NOR3xp33_ASAP7_75t_L g746 ( 
.A(n_690),
.B(n_514),
.C(n_500),
.Y(n_746)
);

BUFx8_ASAP7_75t_L g747 ( 
.A(n_662),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_663),
.B(n_582),
.Y(n_748)
);

BUFx5_ASAP7_75t_L g749 ( 
.A(n_655),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_663),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_655),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_689),
.B(n_427),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_669),
.B(n_606),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_669),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_727),
.A2(n_640),
.B(n_620),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_700),
.B(n_610),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_701),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_SL g758 ( 
.A(n_698),
.B(n_392),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_717),
.B(n_610),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_703),
.B(n_615),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_743),
.A2(n_567),
.B(n_562),
.Y(n_761)
);

OAI21xp33_ASAP7_75t_L g762 ( 
.A1(n_694),
.A2(n_433),
.B(n_431),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_732),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_743),
.A2(n_581),
.B(n_567),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_697),
.A2(n_581),
.B(n_657),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_725),
.B(n_404),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_701),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_712),
.A2(n_657),
.B(n_598),
.Y(n_768)
);

AOI21x1_ASAP7_75t_L g769 ( 
.A1(n_723),
.A2(n_745),
.B(n_727),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_720),
.A2(n_598),
.B(n_594),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_696),
.B(n_413),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_748),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_733),
.A2(n_693),
.B1(n_705),
.B2(n_742),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_706),
.B(n_582),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_724),
.B(n_440),
.Y(n_775)
);

INVxp67_ASAP7_75t_L g776 ( 
.A(n_707),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_704),
.A2(n_710),
.B(n_709),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_705),
.A2(n_477),
.B1(n_532),
.B2(n_484),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_736),
.B(n_719),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_721),
.A2(n_598),
.B(n_594),
.Y(n_780)
);

OAI21x1_ASAP7_75t_SL g781 ( 
.A1(n_699),
.A2(n_616),
.B(n_537),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_751),
.A2(n_671),
.B(n_670),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_737),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_739),
.B(n_551),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_738),
.B(n_629),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_702),
.B(n_552),
.Y(n_786)
);

O2A1O1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_692),
.A2(n_534),
.B(n_553),
.C(n_538),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_695),
.A2(n_600),
.B(n_624),
.C(n_603),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_708),
.A2(n_430),
.B(n_426),
.Y(n_789)
);

NOR2xp67_ASAP7_75t_L g790 ( 
.A(n_741),
.B(n_629),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_751),
.A2(n_672),
.B(n_671),
.Y(n_791)
);

AND2x2_ASAP7_75t_SL g792 ( 
.A(n_730),
.B(n_734),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_731),
.A2(n_713),
.B(n_752),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_730),
.A2(n_435),
.B1(n_438),
.B2(n_434),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_729),
.B(n_453),
.Y(n_795)
);

NOR3xp33_ASAP7_75t_L g796 ( 
.A(n_746),
.B(n_480),
.C(n_463),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_726),
.B(n_632),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_753),
.Y(n_798)
);

O2A1O1Ixp5_ASAP7_75t_L g799 ( 
.A1(n_750),
.A2(n_445),
.B(n_456),
.C(n_450),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_747),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_714),
.A2(n_458),
.B(n_457),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_744),
.B(n_482),
.Y(n_802)
);

INVx4_ASAP7_75t_L g803 ( 
.A(n_711),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_747),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_711),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_728),
.Y(n_806)
);

INVx1_ASAP7_75t_SL g807 ( 
.A(n_715),
.Y(n_807)
);

OAI321xp33_ASAP7_75t_L g808 ( 
.A1(n_716),
.A2(n_642),
.A3(n_641),
.B1(n_638),
.B2(n_612),
.C(n_635),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_718),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_722),
.A2(n_464),
.B(n_462),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_754),
.B(n_504),
.C(n_483),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_728),
.B(n_429),
.Y(n_812)
);

OAI21xp33_ASAP7_75t_L g813 ( 
.A1(n_735),
.A2(n_508),
.B(n_507),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_735),
.A2(n_495),
.B(n_492),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_740),
.B(n_516),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_749),
.A2(n_498),
.B(n_497),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_740),
.A2(n_509),
.B(n_503),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_740),
.A2(n_493),
.B1(n_502),
.B2(n_446),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_749),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_749),
.B(n_518),
.Y(n_820)
);

AO32x1_ASAP7_75t_L g821 ( 
.A1(n_749),
.A2(n_524),
.A3(n_526),
.B1(n_521),
.B2(n_520),
.Y(n_821)
);

NOR2x1_ASAP7_75t_L g822 ( 
.A(n_725),
.B(n_529),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_707),
.B(n_530),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_700),
.B(n_528),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_703),
.A2(n_536),
.B(n_540),
.C(n_535),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_743),
.A2(n_546),
.B(n_543),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_725),
.B(n_544),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_700),
.B(n_545),
.Y(n_828)
);

O2A1O1Ixp5_ASAP7_75t_L g829 ( 
.A1(n_703),
.A2(n_549),
.B(n_550),
.C(n_548),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_743),
.A2(n_556),
.B(n_569),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_700),
.B(n_557),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_737),
.B(n_15),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_703),
.A2(n_400),
.B1(n_410),
.B2(n_397),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_743),
.A2(n_636),
.B(n_425),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_725),
.B(n_415),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_704),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_700),
.B(n_436),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_737),
.Y(n_838)
);

NOR3xp33_ASAP7_75t_L g839 ( 
.A(n_705),
.B(n_439),
.C(n_437),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_748),
.Y(n_840)
);

BUFx8_ASAP7_75t_L g841 ( 
.A(n_737),
.Y(n_841)
);

A2O1A1Ixp33_ASAP7_75t_L g842 ( 
.A1(n_703),
.A2(n_448),
.B(n_451),
.C(n_443),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_700),
.B(n_459),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_743),
.A2(n_636),
.B(n_467),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_700),
.B(n_471),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_743),
.A2(n_473),
.B(n_472),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_743),
.A2(n_479),
.B(n_474),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_706),
.B(n_634),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_743),
.A2(n_485),
.B(n_481),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_725),
.B(n_487),
.Y(n_850)
);

NOR2xp67_ASAP7_75t_L g851 ( 
.A(n_725),
.B(n_496),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_701),
.Y(n_852)
);

AOI21x1_ASAP7_75t_SL g853 ( 
.A1(n_824),
.A2(n_16),
.B(n_17),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_760),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_773),
.A2(n_512),
.B1(n_515),
.B2(n_510),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_798),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_777),
.A2(n_523),
.B(n_519),
.Y(n_857)
);

CKINVDCx8_ASAP7_75t_R g858 ( 
.A(n_800),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_770),
.A2(n_769),
.B(n_755),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_765),
.A2(n_531),
.B(n_527),
.Y(n_860)
);

OAI21x1_ASAP7_75t_L g861 ( 
.A1(n_768),
.A2(n_780),
.B(n_819),
.Y(n_861)
);

AO31x2_ASAP7_75t_L g862 ( 
.A1(n_825),
.A2(n_634),
.A3(n_618),
.B(n_619),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_761),
.A2(n_525),
.B(n_522),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_828),
.A2(n_541),
.B1(n_542),
.B2(n_533),
.Y(n_864)
);

BUFx2_ASAP7_75t_L g865 ( 
.A(n_776),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_779),
.A2(n_816),
.B(n_834),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_797),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_766),
.B(n_18),
.Y(n_868)
);

OAI21x1_ASAP7_75t_L g869 ( 
.A1(n_764),
.A2(n_525),
.B(n_522),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_756),
.B(n_20),
.Y(n_870)
);

INVx2_ASAP7_75t_SL g871 ( 
.A(n_841),
.Y(n_871)
);

OAI21x1_ASAP7_75t_L g872 ( 
.A1(n_830),
.A2(n_525),
.B(n_522),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_783),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_842),
.A2(n_618),
.A3(n_619),
.B(n_613),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_835),
.B(n_21),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_785),
.Y(n_876)
);

NOR2x1_ASAP7_75t_L g877 ( 
.A(n_806),
.B(n_689),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_850),
.B(n_22),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_844),
.A2(n_689),
.B(n_618),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_782),
.A2(n_144),
.B(n_143),
.Y(n_880)
);

AOI211x1_ASAP7_75t_L g881 ( 
.A1(n_793),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_839),
.A2(n_623),
.B1(n_627),
.B2(n_619),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_829),
.A2(n_146),
.B(n_145),
.Y(n_883)
);

AOI21x1_ASAP7_75t_SL g884 ( 
.A1(n_831),
.A2(n_23),
.B(n_25),
.Y(n_884)
);

OAI21x1_ASAP7_75t_L g885 ( 
.A1(n_791),
.A2(n_148),
.B(n_147),
.Y(n_885)
);

AOI221x1_ASAP7_75t_L g886 ( 
.A1(n_833),
.A2(n_639),
.B1(n_644),
.B2(n_627),
.C(n_623),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_772),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_804),
.B(n_27),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_826),
.A2(n_154),
.B(n_151),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_836),
.A2(n_31),
.B1(n_28),
.B2(n_30),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_820),
.A2(n_158),
.B(n_156),
.Y(n_891)
);

AOI221x1_ASAP7_75t_L g892 ( 
.A1(n_789),
.A2(n_644),
.B1(n_639),
.B2(n_627),
.C(n_31),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_822),
.B(n_28),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_838),
.B(n_30),
.Y(n_894)
);

AOI21xp33_ASAP7_75t_L g895 ( 
.A1(n_778),
.A2(n_32),
.B(n_33),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_837),
.A2(n_161),
.B(n_160),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_823),
.B(n_32),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_767),
.B(n_33),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_848),
.B(n_34),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_774),
.B(n_34),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_843),
.B(n_36),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_801),
.A2(n_164),
.B(n_162),
.Y(n_902)
);

INVxp67_ASAP7_75t_L g903 ( 
.A(n_758),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_759),
.B(n_38),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_851),
.B(n_39),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_792),
.B(n_39),
.Y(n_906)
);

AND3x1_ASAP7_75t_SL g907 ( 
.A(n_840),
.B(n_40),
.C(n_41),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_SL g908 ( 
.A(n_757),
.B(n_43),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_794),
.B(n_43),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_841),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_799),
.A2(n_168),
.B(n_167),
.Y(n_911)
);

AND3x4_ASAP7_75t_L g912 ( 
.A(n_796),
.B(n_848),
.C(n_790),
.Y(n_912)
);

OAI21xp33_ASAP7_75t_L g913 ( 
.A1(n_762),
.A2(n_44),
.B(n_45),
.Y(n_913)
);

AO31x2_ASAP7_75t_L g914 ( 
.A1(n_810),
.A2(n_47),
.A3(n_45),
.B(n_46),
.Y(n_914)
);

NOR2xp67_ASAP7_75t_L g915 ( 
.A(n_775),
.B(n_173),
.Y(n_915)
);

AOI21xp33_ASAP7_75t_L g916 ( 
.A1(n_784),
.A2(n_47),
.B(n_48),
.Y(n_916)
);

AND3x4_ASAP7_75t_L g917 ( 
.A(n_763),
.B(n_48),
.C(n_49),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_823),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_809),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_845),
.A2(n_181),
.B(n_180),
.Y(n_920)
);

OAI21x1_ASAP7_75t_L g921 ( 
.A1(n_814),
.A2(n_183),
.B(n_182),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_802),
.B(n_812),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_807),
.B(n_50),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_767),
.B(n_51),
.Y(n_924)
);

NOR4xp25_ASAP7_75t_L g925 ( 
.A(n_787),
.B(n_54),
.C(n_52),
.D(n_53),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_817),
.A2(n_185),
.B(n_184),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_846),
.A2(n_188),
.B(n_186),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_847),
.A2(n_191),
.B(n_189),
.Y(n_928)
);

AOI221xp5_ASAP7_75t_SL g929 ( 
.A1(n_813),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.C(n_59),
.Y(n_929)
);

OA22x2_ASAP7_75t_L g930 ( 
.A1(n_781),
.A2(n_59),
.B1(n_57),
.B2(n_58),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_849),
.A2(n_194),
.B(n_193),
.Y(n_931)
);

OAI21x1_ASAP7_75t_SL g932 ( 
.A1(n_852),
.A2(n_61),
.B(n_62),
.Y(n_932)
);

OR2x6_ASAP7_75t_L g933 ( 
.A(n_832),
.B(n_61),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_757),
.B(n_62),
.Y(n_934)
);

NOR2x1_ASAP7_75t_SL g935 ( 
.A(n_852),
.B(n_757),
.Y(n_935)
);

AOI211x1_ASAP7_75t_L g936 ( 
.A1(n_811),
.A2(n_66),
.B(n_63),
.C(n_65),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_771),
.B(n_67),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_815),
.B(n_68),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_795),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_818),
.B(n_788),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_786),
.B(n_70),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_808),
.A2(n_74),
.B(n_71),
.C(n_73),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_803),
.A2(n_198),
.B(n_197),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_803),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_944)
);

O2A1O1Ixp5_ASAP7_75t_L g945 ( 
.A1(n_821),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_821),
.A2(n_200),
.B(n_199),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_805),
.A2(n_202),
.B(n_201),
.Y(n_947)
);

NAND2x1p5_ASAP7_75t_L g948 ( 
.A(n_800),
.B(n_77),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_78),
.Y(n_949)
);

NOR2xp67_ASAP7_75t_SL g950 ( 
.A(n_757),
.B(n_79),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_770),
.A2(n_208),
.B(n_207),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_800),
.B(n_79),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_768),
.A2(n_211),
.B(n_209),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_829),
.A2(n_215),
.B(n_213),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_770),
.A2(n_219),
.B(n_218),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_SL g956 ( 
.A1(n_767),
.A2(n_221),
.B(n_220),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_827),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_957)
);

OAI21x1_ASAP7_75t_L g958 ( 
.A1(n_770),
.A2(n_225),
.B(n_223),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_800),
.B(n_81),
.Y(n_959)
);

AO31x2_ASAP7_75t_L g960 ( 
.A1(n_825),
.A2(n_82),
.A3(n_83),
.B(n_84),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_777),
.A2(n_230),
.B(n_228),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_760),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_770),
.A2(n_233),
.B(n_232),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_770),
.A2(n_236),
.B(n_235),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_783),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_777),
.A2(n_241),
.B(n_237),
.Y(n_966)
);

INVx4_ASAP7_75t_L g967 ( 
.A(n_757),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_776),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_767),
.B(n_84),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_777),
.A2(n_244),
.B(n_242),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_783),
.B(n_85),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_773),
.B(n_85),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_773),
.B(n_86),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_829),
.A2(n_255),
.B(n_253),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_757),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_773),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_976)
);

AO31x2_ASAP7_75t_L g977 ( 
.A1(n_825),
.A2(n_87),
.A3(n_89),
.B(n_90),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_777),
.A2(n_264),
.B(n_260),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_777),
.A2(n_266),
.B(n_265),
.Y(n_979)
);

BUFx2_ASAP7_75t_L g980 ( 
.A(n_776),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_773),
.B(n_90),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_777),
.A2(n_273),
.B(n_268),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_800),
.B(n_91),
.Y(n_983)
);

INVxp67_ASAP7_75t_SL g984 ( 
.A(n_757),
.Y(n_984)
);

INVx3_ASAP7_75t_SL g985 ( 
.A(n_763),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_800),
.B(n_92),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_777),
.A2(n_279),
.B(n_278),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_827),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_899),
.B(n_94),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_873),
.Y(n_990)
);

AND2x4_ASAP7_75t_L g991 ( 
.A(n_899),
.B(n_96),
.Y(n_991)
);

OAI21xp5_ASAP7_75t_L g992 ( 
.A1(n_866),
.A2(n_901),
.B(n_859),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_875),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_993)
);

AO31x2_ASAP7_75t_L g994 ( 
.A1(n_886),
.A2(n_332),
.A3(n_377),
.B(n_376),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_985),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_SL g996 ( 
.A1(n_878),
.A2(n_100),
.B(n_101),
.C(n_102),
.Y(n_996)
);

CKINVDCx6p67_ASAP7_75t_R g997 ( 
.A(n_918),
.Y(n_997)
);

INVxp67_ASAP7_75t_L g998 ( 
.A(n_965),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_858),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_870),
.A2(n_101),
.B(n_102),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_887),
.Y(n_1001)
);

OAI21x1_ASAP7_75t_SL g1002 ( 
.A1(n_972),
.A2(n_103),
.B(n_104),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_856),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_856),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_919),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_919),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_865),
.B(n_968),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_980),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_904),
.A2(n_105),
.B(n_106),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_967),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_891),
.A2(n_922),
.B(n_883),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_863),
.A2(n_334),
.B(n_375),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_867),
.B(n_107),
.Y(n_1013)
);

OR2x6_ASAP7_75t_L g1014 ( 
.A(n_871),
.B(n_107),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_868),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_SL g1016 ( 
.A1(n_908),
.A2(n_109),
.B(n_111),
.C(n_112),
.Y(n_1016)
);

INVx6_ASAP7_75t_L g1017 ( 
.A(n_952),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_981),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_910),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_952),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_895),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_867),
.B(n_876),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_971),
.B(n_115),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_876),
.Y(n_1024)
);

OR2x2_ASAP7_75t_SL g1025 ( 
.A(n_897),
.B(n_116),
.Y(n_1025)
);

INVxp33_ASAP7_75t_L g1026 ( 
.A(n_894),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_906),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_R g1028 ( 
.A(n_893),
.B(n_280),
.Y(n_1028)
);

OA21x2_ASAP7_75t_L g1029 ( 
.A1(n_869),
.A2(n_338),
.B(n_374),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_937),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_957),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_903),
.B(n_119),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_912),
.A2(n_909),
.B1(n_933),
.B2(n_938),
.Y(n_1033)
);

OAI21x1_ASAP7_75t_L g1034 ( 
.A1(n_951),
.A2(n_340),
.B(n_372),
.Y(n_1034)
);

NOR3xp33_ASAP7_75t_SL g1035 ( 
.A(n_890),
.B(n_120),
.C(n_121),
.Y(n_1035)
);

NOR2xp67_ASAP7_75t_SL g1036 ( 
.A(n_956),
.B(n_120),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_SL g1037 ( 
.A1(n_917),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_975),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_959),
.B(n_122),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_959),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_955),
.A2(n_342),
.B(n_371),
.Y(n_1041)
);

CKINVDCx11_ASAP7_75t_R g1042 ( 
.A(n_983),
.Y(n_1042)
);

AO32x2_ASAP7_75t_L g1043 ( 
.A1(n_976),
.A2(n_123),
.A3(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_1043)
);

AOI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_933),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_954),
.A2(n_281),
.B(n_284),
.Y(n_1045)
);

OAI21x1_ASAP7_75t_L g1046 ( 
.A1(n_958),
.A2(n_287),
.B(n_289),
.Y(n_1046)
);

CKINVDCx11_ASAP7_75t_R g1047 ( 
.A(n_986),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_854),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_962),
.Y(n_1049)
);

AO32x2_ASAP7_75t_L g1050 ( 
.A1(n_944),
.A2(n_296),
.A3(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_963),
.A2(n_301),
.B(n_302),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_986),
.B(n_303),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_855),
.A2(n_306),
.B1(n_307),
.B2(n_309),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_964),
.A2(n_314),
.B(n_315),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_923),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_940),
.B(n_319),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_888),
.B(n_323),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_900),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_941),
.B(n_324),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_892),
.A2(n_325),
.A3(n_326),
.B(n_327),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_974),
.A2(n_329),
.B(n_330),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_916),
.B(n_331),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_934),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_950),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_888),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_935),
.Y(n_1066)
);

OR2x6_ASAP7_75t_L g1067 ( 
.A(n_948),
.B(n_346),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_857),
.A2(n_347),
.B(n_351),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_913),
.A2(n_354),
.B(n_355),
.C(n_356),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_975),
.B(n_357),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_893),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_984),
.B(n_359),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_930),
.B(n_378),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_864),
.B(n_360),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_953),
.A2(n_361),
.B(n_362),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_915),
.B(n_942),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_939),
.B(n_365),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_946),
.A2(n_366),
.B(n_367),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_SL g1079 ( 
.A1(n_928),
.A2(n_889),
.B(n_932),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_905),
.Y(n_1080)
);

INVx3_ASAP7_75t_SL g1081 ( 
.A(n_898),
.Y(n_1081)
);

OR2x2_ASAP7_75t_L g1082 ( 
.A(n_924),
.B(n_369),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_960),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_872),
.A2(n_880),
.B(n_885),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_SL g1085 ( 
.A1(n_969),
.A2(n_988),
.B(n_927),
.C(n_931),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_896),
.A2(n_920),
.B(n_945),
.C(n_947),
.Y(n_1086)
);

OA21x2_ASAP7_75t_L g1087 ( 
.A1(n_902),
.A2(n_879),
.B(n_911),
.Y(n_1087)
);

INVxp67_ASAP7_75t_L g1088 ( 
.A(n_877),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_925),
.A2(n_860),
.B(n_987),
.C(n_982),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_977),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_882),
.B(n_943),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_929),
.A2(n_907),
.B1(n_978),
.B2(n_970),
.C(n_961),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_977),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_921),
.B(n_926),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_914),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_881),
.B(n_936),
.Y(n_1096)
);

AND2x6_ASAP7_75t_L g1097 ( 
.A(n_853),
.B(n_884),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_966),
.B(n_979),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_914),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_874),
.Y(n_1100)
);

INVx1_ASAP7_75t_SL g1101 ( 
.A(n_874),
.Y(n_1101)
);

OAI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_862),
.A2(n_878),
.B1(n_875),
.B2(n_773),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_862),
.A2(n_878),
.B1(n_875),
.B2(n_773),
.Y(n_1103)
);

AOI221x1_ASAP7_75t_L g1104 ( 
.A1(n_862),
.A2(n_946),
.B1(n_972),
.B2(n_973),
.C(n_949),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_873),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_868),
.A2(n_878),
.B(n_875),
.C(n_827),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_865),
.B(n_766),
.Y(n_1107)
);

OA21x2_ASAP7_75t_L g1108 ( 
.A1(n_861),
.A2(n_859),
.B(n_886),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_967),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_865),
.B(n_783),
.Y(n_1110)
);

AOI211xp5_ASAP7_75t_L g1111 ( 
.A1(n_868),
.A2(n_827),
.B(n_766),
.C(n_705),
.Y(n_1111)
);

BUFx2_ASAP7_75t_SL g1112 ( 
.A(n_967),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_887),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_873),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_1083),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1011),
.A2(n_1111),
.B(n_1106),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1110),
.B(n_1007),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1090),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1005),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_1071),
.B(n_1040),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_990),
.B(n_1105),
.Y(n_1121)
);

OAI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1028),
.A2(n_1044),
.B1(n_1033),
.B2(n_1057),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1114),
.B(n_1020),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1008),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1006),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1070),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1001),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1022),
.B(n_1024),
.Y(n_1128)
);

INVx5_ASAP7_75t_L g1129 ( 
.A(n_1057),
.Y(n_1129)
);

INVxp67_ASAP7_75t_L g1130 ( 
.A(n_1107),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_1065),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1113),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1004),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1003),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_999),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_989),
.B(n_991),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1048),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_989),
.B(n_991),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1049),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_997),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_1017),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_998),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1013),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1018),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1039),
.B(n_1023),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1093),
.Y(n_1146)
);

OR2x6_ASAP7_75t_L g1147 ( 
.A(n_1052),
.B(n_1112),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_995),
.Y(n_1148)
);

BUFx8_ASAP7_75t_SL g1149 ( 
.A(n_1014),
.Y(n_1149)
);

INVx8_ASAP7_75t_L g1150 ( 
.A(n_1052),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1030),
.A2(n_1058),
.B1(n_1035),
.B2(n_1000),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_1042),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1056),
.B(n_1055),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1064),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1063),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_1037),
.Y(n_1156)
);

BUFx2_ASAP7_75t_L g1157 ( 
.A(n_1019),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1099),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1095),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1026),
.B(n_1032),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_1109),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1109),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_1102),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1014),
.B(n_1081),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1103),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1002),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1066),
.B(n_1010),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1076),
.B(n_1080),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1047),
.Y(n_1169)
);

AO22x2_ASAP7_75t_L g1170 ( 
.A1(n_1104),
.A2(n_1079),
.B1(n_1101),
.B2(n_1100),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1002),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1104),
.A2(n_1061),
.B(n_1045),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1096),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_996),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_992),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1009),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_993),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1088),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1082),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1043),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1043),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1067),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1015),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1038),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_1091),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1067),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1025),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1027),
.Y(n_1188)
);

INVxp67_ASAP7_75t_L g1189 ( 
.A(n_1112),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1073),
.B(n_1021),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1091),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_1072),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1031),
.B(n_1050),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1077),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1097),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1050),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1059),
.B(n_1074),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1050),
.B(n_1062),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1108),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1036),
.A2(n_1053),
.B1(n_1078),
.B2(n_1092),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1094),
.Y(n_1201)
);

CKINVDCx14_ASAP7_75t_R g1202 ( 
.A(n_1036),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1085),
.B(n_1089),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1087),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1060),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1060),
.B(n_1069),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1117),
.B(n_1145),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1134),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1128),
.B(n_1197),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1121),
.B(n_1060),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1168),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1128),
.B(n_1098),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1130),
.B(n_994),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1137),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1148),
.Y(n_1215)
);

INVx3_ASAP7_75t_SL g1216 ( 
.A(n_1140),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1201),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1139),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1129),
.B(n_1012),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1135),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_SL g1221 ( 
.A1(n_1190),
.A2(n_1068),
.B1(n_1029),
.B2(n_1075),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1197),
.B(n_1086),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1129),
.B(n_1051),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1138),
.B(n_994),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1136),
.B(n_1029),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1127),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_L g1227 ( 
.A(n_1129),
.B(n_1016),
.Y(n_1227)
);

AND2x2_ASAP7_75t_L g1228 ( 
.A(n_1136),
.B(n_1034),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1160),
.B(n_1041),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1156),
.B(n_1046),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1163),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1187),
.B(n_1054),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1132),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1153),
.B(n_1116),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1116),
.B(n_1087),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1119),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1125),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1133),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1124),
.B(n_1084),
.Y(n_1239)
);

INVxp67_ASAP7_75t_L g1240 ( 
.A(n_1168),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1122),
.A2(n_1084),
.B1(n_1193),
.B2(n_1198),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1144),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1142),
.B(n_1123),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1142),
.B(n_1186),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1201),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1131),
.B(n_1120),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1147),
.B(n_1126),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1163),
.B(n_1165),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1118),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1165),
.B(n_1194),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1140),
.Y(n_1251)
);

INVxp67_ASAP7_75t_SL g1252 ( 
.A(n_1118),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1154),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1158),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1152),
.Y(n_1255)
);

NOR2xp67_ASAP7_75t_SL g1256 ( 
.A(n_1169),
.B(n_1182),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1141),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1179),
.Y(n_1258)
);

INVxp67_ASAP7_75t_SL g1259 ( 
.A(n_1196),
.Y(n_1259)
);

NOR2x1_ASAP7_75t_R g1260 ( 
.A(n_1182),
.B(n_1164),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1150),
.B(n_1178),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1196),
.A2(n_1202),
.B1(n_1183),
.B2(n_1122),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1157),
.B(n_1184),
.Y(n_1263)
);

NOR2xp33_ASAP7_75t_L g1264 ( 
.A(n_1126),
.B(n_1202),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1150),
.B(n_1143),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1155),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1151),
.B(n_1161),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1151),
.B(n_1173),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1150),
.B(n_1185),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1176),
.A2(n_1188),
.B1(n_1177),
.B2(n_1200),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1195),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1175),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1146),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1167),
.B(n_1191),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1166),
.Y(n_1275)
);

INVxp67_ASAP7_75t_SL g1276 ( 
.A(n_1231),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1249),
.B(n_1180),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1213),
.B(n_1181),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1253),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1249),
.Y(n_1280)
);

INVxp67_ASAP7_75t_SL g1281 ( 
.A(n_1231),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1241),
.B(n_1170),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1254),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1248),
.B(n_1252),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1236),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1237),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1241),
.B(n_1170),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1238),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1239),
.B(n_1170),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1252),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1209),
.B(n_1189),
.Y(n_1291)
);

BUFx2_ASAP7_75t_L g1292 ( 
.A(n_1272),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1209),
.B(n_1192),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1226),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1259),
.B(n_1199),
.Y(n_1295)
);

HB1xp67_ASAP7_75t_L g1296 ( 
.A(n_1217),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1233),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1217),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1234),
.B(n_1162),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1272),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1242),
.Y(n_1301)
);

OR2x6_ASAP7_75t_SL g1302 ( 
.A(n_1262),
.B(n_1203),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1245),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1224),
.B(n_1205),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1212),
.B(n_1204),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1212),
.B(n_1268),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1247),
.B(n_1115),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1243),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1211),
.B(n_1240),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1208),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1271),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1207),
.B(n_1115),
.Y(n_1312)
);

NOR2x1_ASAP7_75t_L g1313 ( 
.A(n_1250),
.B(n_1174),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1214),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_1220),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1218),
.Y(n_1316)
);

OR2x2_ASAP7_75t_L g1317 ( 
.A(n_1250),
.B(n_1159),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1266),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1306),
.B(n_1275),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1306),
.B(n_1235),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1315),
.B(n_1216),
.Y(n_1321)
);

AND2x4_ASAP7_75t_L g1322 ( 
.A(n_1307),
.B(n_1271),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1289),
.B(n_1235),
.Y(n_1323)
);

INVxp67_ASAP7_75t_L g1324 ( 
.A(n_1280),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1296),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1298),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1303),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1289),
.B(n_1229),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1307),
.B(n_1225),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1278),
.B(n_1210),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1279),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1291),
.B(n_1240),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1307),
.B(n_1273),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1278),
.B(n_1267),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1283),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1305),
.B(n_1270),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1290),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1315),
.Y(n_1338)
);

NOR2xp67_ASAP7_75t_L g1339 ( 
.A(n_1284),
.B(n_1215),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1305),
.B(n_1270),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1285),
.Y(n_1341)
);

OR2x2_ASAP7_75t_L g1342 ( 
.A(n_1284),
.B(n_1262),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_SL g1343 ( 
.A(n_1317),
.B(n_1269),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1290),
.B(n_1274),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1312),
.B(n_1232),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1286),
.Y(n_1346)
);

NAND2xp33_ASAP7_75t_L g1347 ( 
.A(n_1313),
.B(n_1222),
.Y(n_1347)
);

INVxp67_ASAP7_75t_SL g1348 ( 
.A(n_1276),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1334),
.B(n_1308),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1338),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1334),
.B(n_1317),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1331),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1330),
.B(n_1292),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1335),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1341),
.Y(n_1355)
);

NOR2x1_ASAP7_75t_L g1356 ( 
.A(n_1321),
.B(n_1220),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1346),
.Y(n_1357)
);

NAND3xp33_ASAP7_75t_L g1358 ( 
.A(n_1347),
.B(n_1222),
.C(n_1309),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1332),
.B(n_1312),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1324),
.B(n_1311),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1320),
.B(n_1295),
.Y(n_1361)
);

OAI21xp33_ASAP7_75t_L g1362 ( 
.A1(n_1336),
.A2(n_1287),
.B(n_1282),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1345),
.B(n_1292),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1345),
.B(n_1300),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1336),
.B(n_1281),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1325),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1340),
.B(n_1320),
.Y(n_1367)
);

INVx3_ASAP7_75t_L g1368 ( 
.A(n_1322),
.Y(n_1368)
);

NOR2x1_ASAP7_75t_L g1369 ( 
.A(n_1347),
.B(n_1311),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1326),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1327),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1328),
.B(n_1300),
.Y(n_1372)
);

INVxp67_ASAP7_75t_SL g1373 ( 
.A(n_1348),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1352),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1358),
.A2(n_1287),
.B1(n_1282),
.B2(n_1230),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1373),
.B(n_1340),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1373),
.B(n_1365),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1354),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1367),
.A2(n_1302),
.B1(n_1342),
.B2(n_1339),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1369),
.B(n_1343),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1355),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1357),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1366),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1361),
.B(n_1319),
.Y(n_1384)
);

AOI322xp5_ASAP7_75t_L g1385 ( 
.A1(n_1362),
.A2(n_1330),
.A3(n_1323),
.B1(n_1328),
.B2(n_1319),
.C1(n_1293),
.C2(n_1206),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1361),
.B(n_1337),
.Y(n_1386)
);

AOI322xp5_ASAP7_75t_L g1387 ( 
.A1(n_1359),
.A2(n_1323),
.A3(n_1304),
.B1(n_1302),
.B2(n_1349),
.C1(n_1221),
.C2(n_1360),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1360),
.B(n_1344),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1351),
.B(n_1342),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1370),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1371),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1374),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1376),
.B(n_1363),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1388),
.B(n_1216),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1387),
.B(n_1364),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1389),
.B(n_1353),
.Y(n_1396)
);

OAI31xp33_ASAP7_75t_L g1397 ( 
.A1(n_1379),
.A2(n_1310),
.A3(n_1314),
.B(n_1316),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1380),
.A2(n_1356),
.B(n_1350),
.Y(n_1398)
);

INVxp67_ASAP7_75t_L g1399 ( 
.A(n_1383),
.Y(n_1399)
);

OAI21xp33_ASAP7_75t_L g1400 ( 
.A1(n_1395),
.A2(n_1377),
.B(n_1380),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1397),
.A2(n_1375),
.B(n_1390),
.Y(n_1401)
);

AOI211xp5_ASAP7_75t_L g1402 ( 
.A1(n_1398),
.A2(n_1256),
.B(n_1375),
.C(n_1260),
.Y(n_1402)
);

AOI221xp5_ASAP7_75t_L g1403 ( 
.A1(n_1392),
.A2(n_1391),
.B1(n_1378),
.B2(n_1381),
.C(n_1382),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1394),
.A2(n_1329),
.B1(n_1333),
.B2(n_1264),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1401),
.B(n_1396),
.Y(n_1405)
);

XNOR2xp5_ASAP7_75t_L g1406 ( 
.A(n_1402),
.B(n_1255),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1403),
.B(n_1399),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1400),
.A2(n_1393),
.B(n_1350),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1404),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_L g1410 ( 
.A(n_1400),
.B(n_1257),
.C(n_1264),
.Y(n_1410)
);

NOR4xp25_ASAP7_75t_L g1411 ( 
.A(n_1407),
.B(n_1244),
.C(n_1263),
.D(n_1246),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1410),
.A2(n_1409),
.B1(n_1405),
.B2(n_1406),
.Y(n_1412)
);

OAI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1408),
.A2(n_1385),
.B1(n_1221),
.B2(n_1227),
.C(n_1172),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1412),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_SL g1415 ( 
.A(n_1411),
.B(n_1251),
.Y(n_1415)
);

AND3x4_ASAP7_75t_L g1416 ( 
.A(n_1415),
.B(n_1149),
.C(n_1413),
.Y(n_1416)
);

NAND5xp2_ASAP7_75t_L g1417 ( 
.A(n_1416),
.B(n_1414),
.C(n_1149),
.D(n_1171),
.E(n_1372),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1417),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1417),
.A2(n_1223),
.B1(n_1288),
.B2(n_1294),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1419),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1418),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1421),
.A2(n_1386),
.B(n_1384),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1420),
.A2(n_1277),
.B1(n_1299),
.B2(n_1265),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1423),
.A2(n_1422),
.B1(n_1258),
.B2(n_1228),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1423),
.A2(n_1223),
.B1(n_1258),
.B2(n_1219),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1424),
.A2(n_1261),
.B(n_1368),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1426),
.B(n_1425),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1427),
.A2(n_1297),
.B1(n_1301),
.B2(n_1318),
.Y(n_1428)
);


endmodule