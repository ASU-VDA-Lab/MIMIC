module fake_netlist_5_1967_n_821 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_821);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_821;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_804;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_750;
wire n_472;
wire n_742;
wire n_669;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_727;
wire n_311;
wire n_813;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

BUFx3_ASAP7_75t_L g158 ( 
.A(n_35),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_29),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_57),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_115),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_19),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_62),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_119),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_31),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_131),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_152),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_154),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_6),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_140),
.Y(n_179)
);

NOR2xp67_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_40),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_84),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_60),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_16),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_153),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_85),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_11),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_4),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_96),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_25),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_102),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_41),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_47),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_92),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_2),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_4),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_134),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_82),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_97),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_32),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_88),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_108),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_112),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_147),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_7),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_16),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_126),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_20),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_50),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_24),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_151),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_117),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_178),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_165),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

BUFx8_ASAP7_75t_SL g228 ( 
.A(n_166),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_190),
.B(n_0),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

OAI21x1_ASAP7_75t_L g232 ( 
.A1(n_172),
.A2(n_1),
.B(n_2),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_166),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_158),
.B(n_21),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_1),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_3),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_199),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g239 ( 
.A(n_158),
.B(n_22),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_3),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_168),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_209),
.B(n_23),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g250 ( 
.A(n_168),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_251)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_159),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_5),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_160),
.Y(n_256)
);

INVxp33_ASAP7_75t_SL g257 ( 
.A(n_162),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_8),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_164),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_219),
.Y(n_261)
);

BUFx8_ASAP7_75t_SL g262 ( 
.A(n_175),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_179),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_171),
.B(n_9),
.Y(n_264)
);

BUFx8_ASAP7_75t_SL g265 ( 
.A(n_179),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_185),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_186),
.B(n_10),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_228),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_233),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_262),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_265),
.Y(n_276)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_252),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_234),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_250),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_204),
.B1(n_197),
.B2(n_191),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_250),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_257),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_244),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_223),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_223),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_R g290 ( 
.A(n_227),
.B(n_167),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_227),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_224),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_R g293 ( 
.A(n_224),
.B(n_169),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_246),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_266),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_267),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_247),
.B(n_173),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_267),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_261),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_198),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_237),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_R g303 ( 
.A(n_237),
.B(n_176),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_SL g304 ( 
.A(n_254),
.B(n_219),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_239),
.B(n_202),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_245),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_256),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_256),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_235),
.B(n_205),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_256),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_239),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_230),
.B(n_207),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_240),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_R g317 ( 
.A(n_260),
.B(n_177),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

OR2x6_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_251),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g320 ( 
.A(n_282),
.B(n_268),
.C(n_264),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_289),
.B(n_260),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_258),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_305),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_269),
.B(n_181),
.Y(n_324)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_254),
.C(n_249),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_239),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_258),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_249),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_315),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_314),
.B(n_249),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_236),
.C(n_229),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_316),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_273),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_284),
.B(n_180),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_318),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_284),
.B(n_255),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_275),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_255),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_255),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_308),
.B(n_248),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_306),
.B(n_219),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_255),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_270),
.Y(n_344)
);

NAND3xp33_ASAP7_75t_L g345 ( 
.A(n_302),
.B(n_229),
.C(n_236),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_296),
.Y(n_346)
);

NAND3xp33_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_241),
.C(n_226),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_271),
.B(n_241),
.C(n_231),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_278),
.Y(n_351)
);

OR2x2_ASAP7_75t_SL g352 ( 
.A(n_303),
.B(n_211),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_312),
.B(n_304),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_297),
.B(n_248),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_301),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_278),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_317),
.B(n_242),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_303),
.A2(n_232),
.B1(n_225),
.B2(n_243),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_290),
.B(n_242),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_295),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_290),
.B(n_242),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_299),
.B(n_219),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_307),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_291),
.B(n_215),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_285),
.B(n_242),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_287),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_293),
.B(n_242),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_281),
.B(n_225),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_279),
.Y(n_371)
);

A2O1A1Ixp33_ASAP7_75t_L g372 ( 
.A1(n_277),
.A2(n_232),
.B(n_243),
.C(n_238),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_272),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_277),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_283),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_292),
.B(n_255),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_274),
.B(n_184),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_276),
.B(n_188),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_313),
.B(n_216),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_313),
.B(n_217),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g382 ( 
.A(n_289),
.B(n_189),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_280),
.B(n_193),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_305),
.Y(n_384)
);

OAI221xp5_ASAP7_75t_L g385 ( 
.A1(n_328),
.A2(n_331),
.B1(n_330),
.B2(n_325),
.C(n_320),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_366),
.B(n_194),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_336),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_328),
.B(n_195),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_330),
.B(n_196),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_364),
.A2(n_210),
.B1(n_222),
.B2(n_221),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_201),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_338),
.Y(n_393)
);

NAND2x1p5_ASAP7_75t_L g394 ( 
.A(n_337),
.B(n_238),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_332),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_348),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_327),
.A2(n_208),
.B(n_206),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_358),
.B(n_203),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_321),
.B(n_212),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_R g401 ( 
.A(n_373),
.B(n_27),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_358),
.B(n_343),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_382),
.B(n_12),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_345),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_323),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_13),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_354),
.B(n_14),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_15),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g410 ( 
.A(n_354),
.B(n_15),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_367),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_340),
.B(n_28),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_333),
.B(n_30),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_365),
.B(n_17),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_349),
.B(n_340),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_342),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_384),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

AOI22xp33_ASAP7_75t_L g423 ( 
.A1(n_341),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_341),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g425 ( 
.A1(n_322),
.A2(n_18),
.B1(n_34),
.B2(n_36),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_351),
.Y(n_426)
);

NAND3xp33_ASAP7_75t_SL g427 ( 
.A(n_363),
.B(n_37),
.C(n_38),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_355),
.B(n_39),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_359),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_347),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_374),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_367),
.B(n_42),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_356),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_360),
.B(n_43),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_44),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_357),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_334),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_376),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_334),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_363),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_368),
.Y(n_443)
);

AND2x6_ASAP7_75t_L g444 ( 
.A(n_353),
.B(n_45),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_377),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_372),
.B(n_46),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_372),
.B(n_370),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

AOI21x1_ASAP7_75t_L g451 ( 
.A1(n_380),
.A2(n_48),
.B(n_49),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_378),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

NOR3xp33_ASAP7_75t_SL g455 ( 
.A(n_370),
.B(n_361),
.C(n_379),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_412),
.B(n_375),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_402),
.A2(n_319),
.B(n_324),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_402),
.A2(n_319),
.B(n_52),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

O2A1O1Ixp33_ASAP7_75t_L g460 ( 
.A1(n_385),
.A2(n_319),
.B(n_53),
.C(n_54),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_408),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_396),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_430),
.B(n_51),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_415),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_55),
.Y(n_465)
);

O2A1O1Ixp33_ASAP7_75t_L g466 ( 
.A1(n_385),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_466)
);

BUFx3_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_404),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_449),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_69),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g471 ( 
.A(n_432),
.B(n_442),
.Y(n_471)
);

AOI21xp5_ASAP7_75t_L g472 ( 
.A1(n_437),
.A2(n_70),
.B(n_71),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_416),
.A2(n_454),
.B1(n_446),
.B2(n_452),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_72),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_453),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_475)
);

AND2x4_ASAP7_75t_SL g476 ( 
.A(n_450),
.B(n_76),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_415),
.Y(n_478)
);

O2A1O1Ixp33_ASAP7_75t_L g479 ( 
.A1(n_449),
.A2(n_77),
.B(n_80),
.C(n_81),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_437),
.A2(n_392),
.B(n_390),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_392),
.A2(n_83),
.B(n_86),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_406),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_SL g483 ( 
.A(n_432),
.B(n_87),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_419),
.A2(n_157),
.B(n_90),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_443),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_89),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_441),
.B(n_91),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_389),
.B(n_94),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_397),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_390),
.A2(n_98),
.B(n_99),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_397),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_431),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_407),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_386),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_435),
.A2(n_100),
.B(n_103),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_389),
.B(n_104),
.Y(n_498)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_414),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_109),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

A2O1A1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_414),
.A2(n_110),
.B(n_114),
.C(n_116),
.Y(n_503)
);

O2A1O1Ixp33_ASAP7_75t_L g504 ( 
.A1(n_399),
.A2(n_118),
.B(n_120),
.C(n_121),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_399),
.A2(n_122),
.B(n_123),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_388),
.B(n_125),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_455),
.B(n_391),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_440),
.B(n_127),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_387),
.B(n_128),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_435),
.A2(n_129),
.B(n_132),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_418),
.B(n_133),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_464),
.Y(n_513)
);

INVx6_ASAP7_75t_SL g514 ( 
.A(n_461),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_486),
.Y(n_515)
);

OAI22xp33_ASAP7_75t_L g516 ( 
.A1(n_495),
.A2(n_432),
.B1(n_448),
.B2(n_424),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_484),
.A2(n_436),
.B(n_448),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_462),
.Y(n_518)
);

OA21x2_ASAP7_75t_L g519 ( 
.A1(n_480),
.A2(n_436),
.B(n_428),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_482),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_497),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_464),
.B(n_419),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_490),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_493),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_393),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_464),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_478),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_496),
.Y(n_529)
);

INVx6_ASAP7_75t_SL g530 ( 
.A(n_461),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_467),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_478),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_451),
.B(n_434),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_478),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_388),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_501),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_388),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_459),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_506),
.A2(n_422),
.B(n_426),
.Y(n_540)
);

AO21x2_ASAP7_75t_L g541 ( 
.A1(n_458),
.A2(n_398),
.B(n_427),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_482),
.Y(n_542)
);

BUFx4f_ASAP7_75t_SL g543 ( 
.A(n_507),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_505),
.A2(n_433),
.B(n_398),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_459),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_474),
.A2(n_420),
.B(n_413),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_485),
.Y(n_547)
);

BUFx2_ASAP7_75t_SL g548 ( 
.A(n_471),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_492),
.B(n_400),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_508),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_502),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_463),
.A2(n_421),
.B(n_425),
.Y(n_552)
);

AO21x2_ASAP7_75t_L g553 ( 
.A1(n_488),
.A2(n_401),
.B(n_409),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_473),
.B(n_457),
.Y(n_554)
);

BUFx12f_ASAP7_75t_L g555 ( 
.A(n_470),
.Y(n_555)
);

CKINVDCx6p67_ASAP7_75t_R g556 ( 
.A(n_498),
.Y(n_556)
);

OAI21x1_ASAP7_75t_L g557 ( 
.A1(n_472),
.A2(n_491),
.B(n_481),
.Y(n_557)
);

INVx2_ASAP7_75t_R g558 ( 
.A(n_466),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_465),
.Y(n_559)
);

BUFx2_ASAP7_75t_SL g560 ( 
.A(n_509),
.Y(n_560)
);

OAI21x1_ASAP7_75t_L g561 ( 
.A1(n_540),
.A2(n_511),
.B(n_479),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_542),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_529),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_SL g564 ( 
.A1(n_543),
.A2(n_468),
.B1(n_487),
.B2(n_500),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_540),
.A2(n_504),
.B(n_510),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_518),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_521),
.Y(n_567)
);

OAI21x1_ASAP7_75t_L g568 ( 
.A1(n_533),
.A2(n_460),
.B(n_469),
.Y(n_568)
);

AOI21x1_ASAP7_75t_L g569 ( 
.A1(n_517),
.A2(n_483),
.B(n_469),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_554),
.A2(n_432),
.B1(n_512),
.B2(n_423),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_529),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_525),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_535),
.B(n_476),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

INVx2_ASAP7_75t_SL g575 ( 
.A(n_531),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_552),
.A2(n_559),
.B(n_516),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_537),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_547),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_524),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_409),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_527),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_536),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_520),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_551),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_546),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_545),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_545),
.Y(n_590)
);

OAI21xp33_ASAP7_75t_SL g591 ( 
.A1(n_559),
.A2(n_503),
.B(n_499),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_550),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_519),
.A2(n_517),
.B(n_557),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_546),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_515),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_513),
.B(n_409),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_532),
.Y(n_598)
);

INVx8_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_SL g600 ( 
.A1(n_536),
.A2(n_444),
.B1(n_393),
.B2(n_429),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_533),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_545),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_557),
.A2(n_393),
.B(n_475),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_545),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_578),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_581),
.B(n_515),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_578),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_R g608 ( 
.A(n_583),
.B(n_549),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_584),
.B(n_556),
.Y(n_609)
);

NAND2x1_ASAP7_75t_L g610 ( 
.A(n_602),
.B(n_513),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_573),
.B(n_532),
.Y(n_611)
);

CKINVDCx16_ASAP7_75t_R g612 ( 
.A(n_596),
.Y(n_612)
);

INVx6_ASAP7_75t_SL g613 ( 
.A(n_580),
.Y(n_613)
);

INVx3_ASAP7_75t_SL g614 ( 
.A(n_583),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_566),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_562),
.B(n_556),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_585),
.Y(n_617)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_576),
.A2(n_593),
.B(n_570),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_586),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_599),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_567),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_L g622 ( 
.A1(n_564),
.A2(n_538),
.B(n_544),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_585),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_580),
.B(n_555),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_R g626 ( 
.A(n_596),
.B(n_555),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_513),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_580),
.B(n_528),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_592),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_599),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_R g631 ( 
.A(n_575),
.B(n_527),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_587),
.Y(n_632)
);

O2A1O1Ixp33_ASAP7_75t_L g633 ( 
.A1(n_591),
.A2(n_538),
.B(n_553),
.C(n_541),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_R g634 ( 
.A(n_597),
.B(n_598),
.Y(n_634)
);

NAND3xp33_ASAP7_75t_SL g635 ( 
.A(n_600),
.B(n_538),
.C(n_523),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_575),
.B(n_528),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_597),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_599),
.A2(n_560),
.B1(n_444),
.B2(n_541),
.Y(n_638)
);

INVx4_ASAP7_75t_L g639 ( 
.A(n_599),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_577),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_577),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_563),
.B(n_528),
.Y(n_643)
);

NAND2xp33_ASAP7_75t_R g644 ( 
.A(n_589),
.B(n_522),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_582),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_579),
.A2(n_444),
.B1(n_553),
.B2(n_548),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_563),
.B(n_527),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_571),
.B(n_586),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_594),
.A2(n_572),
.B(n_553),
.C(n_541),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_571),
.B(n_534),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_572),
.A2(n_444),
.B1(n_534),
.B2(n_527),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_R g652 ( 
.A(n_589),
.B(n_522),
.Y(n_652)
);

BUFx10_ASAP7_75t_L g653 ( 
.A(n_582),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_582),
.B(n_534),
.Y(n_654)
);

NOR3xp33_ASAP7_75t_SL g655 ( 
.A(n_590),
.B(n_514),
.C(n_530),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_574),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_574),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_631),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_624),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_632),
.B(n_601),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_640),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_642),
.B(n_650),
.Y(n_662)
);

AOI21xp33_ASAP7_75t_L g663 ( 
.A1(n_622),
.A2(n_633),
.B(n_649),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_615),
.B(n_601),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_611),
.A2(n_558),
.B1(n_530),
.B2(n_514),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_621),
.B(n_595),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_629),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_657),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_623),
.B(n_582),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_608),
.A2(n_634),
.B1(n_612),
.B2(n_616),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_656),
.B(n_588),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_605),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_607),
.B(n_588),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_619),
.B(n_595),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_617),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_606),
.Y(n_676)
);

AO22x1_ASAP7_75t_L g677 ( 
.A1(n_620),
.A2(n_630),
.B1(n_609),
.B2(n_636),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_648),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_647),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_641),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_643),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_637),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_646),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_654),
.Y(n_684)
);

INVxp67_ASAP7_75t_L g685 ( 
.A(n_627),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_653),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_628),
.B(n_527),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_646),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

NAND2x1_ASAP7_75t_L g690 ( 
.A(n_639),
.B(n_522),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_611),
.B(n_530),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_638),
.B(n_651),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_645),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_620),
.B(n_590),
.Y(n_694)
);

AOI211xp5_ASAP7_75t_SL g695 ( 
.A1(n_635),
.A2(n_604),
.B(n_602),
.C(n_558),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_653),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_651),
.B(n_568),
.Y(n_697)
);

AND2x4_ASAP7_75t_SL g698 ( 
.A(n_639),
.B(n_604),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_610),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_662),
.B(n_568),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_662),
.B(n_569),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_659),
.B(n_569),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_659),
.B(n_565),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_661),
.B(n_565),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_667),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_675),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_661),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_666),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_666),
.B(n_603),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_664),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_664),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_660),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_683),
.B(n_688),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_670),
.A2(n_676),
.B1(n_689),
.B2(n_692),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_660),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_689),
.B(n_625),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_668),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_668),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_697),
.B(n_603),
.Y(n_719)
);

AOI221xp5_ASAP7_75t_L g720 ( 
.A1(n_663),
.A2(n_655),
.B1(n_626),
.B2(n_534),
.C(n_614),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_671),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_681),
.B(n_630),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_667),
.B(n_561),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_679),
.B(n_678),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_671),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_672),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_685),
.B(n_561),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_672),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_665),
.B(n_652),
.C(n_644),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_706),
.B(n_677),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_684),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_716),
.B(n_693),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_727),
.B(n_697),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_707),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_707),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_718),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_700),
.B(n_719),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_716),
.B(n_677),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_705),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_726),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_724),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_700),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_708),
.B(n_680),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_713),
.B(n_692),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_717),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_719),
.B(n_695),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_717),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_714),
.A2(n_682),
.B1(n_613),
.B2(n_691),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_701),
.B(n_673),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_728),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_741),
.B(n_701),
.Y(n_751)
);

OA222x2_ASAP7_75t_L g752 ( 
.A1(n_738),
.A2(n_725),
.B1(n_721),
.B2(n_715),
.C1(n_712),
.C2(n_710),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_745),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_735),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_732),
.B(n_713),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_737),
.B(n_711),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_745),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_749),
.B(n_702),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_730),
.B(n_729),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_740),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_SL g761 ( 
.A(n_746),
.B(n_684),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_750),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_734),
.Y(n_763)
);

NAND4xp75_ASAP7_75t_SL g764 ( 
.A(n_746),
.B(n_732),
.C(n_703),
.D(n_704),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_739),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_754),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_759),
.B(n_744),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_755),
.Y(n_768)
);

INVxp33_ASAP7_75t_L g769 ( 
.A(n_761),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_759),
.A2(n_714),
.B(n_748),
.Y(n_770)
);

NAND4xp25_ASAP7_75t_L g771 ( 
.A(n_761),
.B(n_748),
.C(n_720),
.D(n_722),
.Y(n_771)
);

BUFx3_ASAP7_75t_L g772 ( 
.A(n_766),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_767),
.B(n_759),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_768),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_770),
.B(n_762),
.Y(n_775)
);

OAI221xp5_ASAP7_75t_L g776 ( 
.A1(n_771),
.A2(n_765),
.B1(n_751),
.B2(n_760),
.C(n_682),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_769),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_772),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_775),
.B(n_758),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_777),
.B(n_752),
.Y(n_780)
);

NOR3x1_ASAP7_75t_L g781 ( 
.A(n_776),
.B(n_658),
.C(n_758),
.Y(n_781)
);

OAI31xp33_ASAP7_75t_L g782 ( 
.A1(n_780),
.A2(n_775),
.A3(n_773),
.B(n_774),
.Y(n_782)
);

AOI221x1_ASAP7_75t_SL g783 ( 
.A1(n_778),
.A2(n_763),
.B1(n_736),
.B2(n_757),
.C(n_753),
.Y(n_783)
);

NAND4xp25_ASAP7_75t_SL g784 ( 
.A(n_779),
.B(n_733),
.C(n_764),
.D(n_756),
.Y(n_784)
);

AOI221xp5_ASAP7_75t_L g785 ( 
.A1(n_782),
.A2(n_781),
.B1(n_747),
.B2(n_742),
.C(n_669),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_783),
.A2(n_658),
.B(n_696),
.C(n_731),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_784),
.A2(n_731),
.B1(n_694),
.B2(n_749),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_SL g788 ( 
.A1(n_782),
.A2(n_686),
.B(n_699),
.C(n_514),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_786),
.Y(n_789)
);

NOR2x1_ASAP7_75t_L g790 ( 
.A(n_788),
.B(n_534),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_787),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_785),
.A2(n_694),
.B1(n_703),
.B2(n_704),
.Y(n_792)
);

OAI211xp5_ASAP7_75t_SL g793 ( 
.A1(n_788),
.A2(n_687),
.B(n_743),
.C(n_699),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_787),
.B(n_737),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_791),
.B(n_747),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_789),
.B(n_135),
.Y(n_796)
);

NOR2x1_ASAP7_75t_L g797 ( 
.A(n_790),
.B(n_686),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_794),
.Y(n_798)
);

OR2x2_ASAP7_75t_L g799 ( 
.A(n_792),
.B(n_793),
.Y(n_799)
);

NAND4xp75_ASAP7_75t_L g800 ( 
.A(n_790),
.B(n_702),
.C(n_734),
.D(n_519),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_791),
.B(n_694),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_796),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_798),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_801),
.Y(n_804)
);

NOR2x1_ASAP7_75t_L g805 ( 
.A(n_797),
.B(n_690),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_795),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_SL g807 ( 
.A(n_802),
.B(n_799),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_803),
.A2(n_800),
.B1(n_698),
.B2(n_690),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_806),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_804),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_809),
.A2(n_805),
.B1(n_613),
.B2(n_698),
.Y(n_811)
);

AO22x2_ASAP7_75t_L g812 ( 
.A1(n_810),
.A2(n_674),
.B1(n_673),
.B2(n_709),
.Y(n_812)
);

BUFx2_ASAP7_75t_L g813 ( 
.A(n_807),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_808),
.B(n_709),
.Y(n_814)
);

OAI22x1_ASAP7_75t_L g815 ( 
.A1(n_813),
.A2(n_523),
.B1(n_519),
.B2(n_674),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_811),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_816),
.A2(n_814),
.B(n_812),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_817),
.Y(n_818)
);

AOI222xp33_ASAP7_75t_L g819 ( 
.A1(n_818),
.A2(n_815),
.B1(n_544),
.B2(n_139),
.C1(n_142),
.C2(n_145),
.Y(n_819)
);

OR2x6_ASAP7_75t_L g820 ( 
.A(n_819),
.B(n_429),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_820),
.A2(n_136),
.B1(n_138),
.B2(n_146),
.Y(n_821)
);


endmodule