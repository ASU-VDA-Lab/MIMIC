module fake_aes_3253_n_562 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_562);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_562;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_0), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_9), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_29), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_76), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_47), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_72), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_16), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_3), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_22), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_21), .Y(n_88) );
CKINVDCx16_ASAP7_75t_R g89 ( .A(n_62), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_40), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_34), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_51), .Y(n_92) );
OR2x2_ASAP7_75t_L g93 ( .A(n_66), .B(n_13), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_58), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_0), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_8), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_19), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_30), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_3), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_73), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_54), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_60), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_17), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_37), .Y(n_105) );
INVx3_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_45), .Y(n_107) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_78), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_27), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_1), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_31), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_11), .Y(n_118) );
CKINVDCx16_ASAP7_75t_R g119 ( .A(n_50), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_36), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_101), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
AND2x4_ASAP7_75t_L g124 ( .A(n_106), .B(n_1), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_81), .A2(n_41), .B(n_75), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_106), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_104), .B(n_2), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_104), .B(n_2), .Y(n_128) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_93), .B(n_39), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
INVx2_ASAP7_75t_SL g131 ( .A(n_88), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_94), .A2(n_43), .B(n_74), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_101), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_94), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
BUFx2_ASAP7_75t_L g136 ( .A(n_83), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_95), .B(n_4), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_79), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_97), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_79), .B(n_4), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_80), .B(n_5), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_124), .Y(n_143) );
INVx1_ASAP7_75t_SL g144 ( .A(n_136), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_130), .B(n_98), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_136), .B(n_138), .Y(n_146) );
INVx2_ASAP7_75t_SL g147 ( .A(n_124), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_136), .B(n_89), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_130), .B(n_98), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_142), .B(n_112), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_142), .B(n_89), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_122), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_124), .B(n_102), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_124), .B(n_80), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_122), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_137), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_121), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_141), .B(n_86), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_138), .B(n_99), .Y(n_164) );
AND2x6_ASAP7_75t_L g165 ( .A(n_141), .B(n_102), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_121), .B(n_120), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_134), .B(n_116), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_127), .B(n_95), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_151), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_152), .B(n_127), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_168), .A2(n_137), .B1(n_129), .B2(n_128), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_162), .Y(n_172) );
INVx2_ASAP7_75t_SL g173 ( .A(n_151), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_144), .B(n_128), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
BUFx4f_ASAP7_75t_L g176 ( .A(n_157), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g177 ( .A1(n_147), .A2(n_132), .B(n_125), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_143), .B(n_129), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_146), .B(n_134), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_144), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_146), .B(n_135), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_162), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_158), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_164), .B(n_135), .Y(n_184) );
INVx5_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
INVx2_ASAP7_75t_SL g186 ( .A(n_158), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_164), .B(n_139), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_157), .Y(n_190) );
INVx2_ASAP7_75t_SL g191 ( .A(n_157), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_163), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_148), .B(n_139), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_148), .B(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_143), .B(n_129), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_147), .Y(n_197) );
INVx5_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
NAND3xp33_ASAP7_75t_SL g199 ( .A(n_160), .B(n_117), .C(n_115), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_147), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
OR2x6_ASAP7_75t_L g202 ( .A(n_150), .B(n_129), .Y(n_202) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_180), .A2(n_168), .B1(n_150), .B2(n_85), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_178), .A2(n_163), .B(n_149), .Y(n_204) );
AOI221xp5_ASAP7_75t_L g205 ( .A1(n_184), .A2(n_153), .B1(n_166), .B2(n_141), .C(n_140), .Y(n_205) );
INVx4_ASAP7_75t_L g206 ( .A(n_176), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_180), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_197), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_171), .A2(n_165), .B1(n_157), .B2(n_141), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_178), .A2(n_167), .B(n_145), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_176), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_174), .B(n_193), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_170), .A2(n_167), .B(n_149), .C(n_145), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_197), .Y(n_215) );
BUFx12f_ASAP7_75t_L g216 ( .A(n_202), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_187), .B(n_157), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_179), .B(n_157), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_181), .B(n_195), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_202), .A2(n_165), .B1(n_131), .B2(n_140), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_200), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_202), .A2(n_126), .B1(n_107), .B2(n_119), .Y(n_223) );
BUFx4_ASAP7_75t_SL g224 ( .A(n_202), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_199), .B(n_165), .Y(n_226) );
AOI22xp5_ASAP7_75t_L g227 ( .A1(n_186), .A2(n_165), .B1(n_126), .B2(n_131), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_194), .B(n_165), .Y(n_228) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_177), .A2(n_109), .B(n_113), .Y(n_229) );
BUFx3_ASAP7_75t_L g230 ( .A(n_185), .Y(n_230) );
INVx4_ASAP7_75t_L g231 ( .A(n_176), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_194), .B(n_165), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_185), .B(n_99), .Y(n_233) );
INVx2_ASAP7_75t_SL g234 ( .A(n_186), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_182), .A2(n_131), .B(n_93), .C(n_109), .Y(n_235) );
OAI21x1_ASAP7_75t_SL g236 ( .A1(n_190), .A2(n_125), .B(n_132), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_203), .A2(n_194), .B1(n_165), .B2(n_192), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_213), .B(n_201), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_207), .B(n_183), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_209), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_207), .Y(n_242) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_236), .A2(n_196), .B(n_103), .Y(n_243) );
BUFx2_ASAP7_75t_L g244 ( .A(n_216), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_213), .B(n_188), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_203), .B(n_189), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_236), .A2(n_196), .B(n_132), .Y(n_247) );
OA21x2_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_103), .B(n_105), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_204), .A2(n_125), .B(n_132), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_224), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_208), .Y(n_251) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_223), .A2(n_165), .B1(n_169), .B2(n_175), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_216), .B(n_169), .Y(n_253) );
INVx1_ASAP7_75t_SL g254 ( .A(n_223), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_208), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_217), .A2(n_125), .B(n_132), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_215), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_215), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_222), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_217), .A2(n_125), .B(n_200), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_235), .A2(n_100), .B(n_86), .C(n_114), .Y(n_261) );
NAND4xp25_ASAP7_75t_SL g262 ( .A(n_210), .B(n_96), .C(n_111), .D(n_114), .Y(n_262) );
OAI222xp33_ASAP7_75t_L g263 ( .A1(n_210), .A2(n_119), .B1(n_107), .B2(n_96), .C1(n_111), .C2(n_118), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g264 ( .A(n_206), .B(n_185), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_214), .A2(n_173), .B(n_191), .Y(n_265) );
AOI211xp5_ASAP7_75t_SL g266 ( .A1(n_263), .A2(n_226), .B(n_220), .C(n_227), .Y(n_266) );
AOI221xp5_ASAP7_75t_L g267 ( .A1(n_246), .A2(n_205), .B1(n_221), .B2(n_118), .C(n_218), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_254), .B(n_242), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_245), .B(n_219), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_240), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_265), .A2(n_229), .B(n_222), .Y(n_271) );
OR2x6_ASAP7_75t_L g272 ( .A(n_250), .B(n_206), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_265), .A2(n_229), .B(n_233), .Y(n_273) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_254), .A2(n_234), .B1(n_228), .B2(n_175), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_262), .A2(n_234), .B1(n_175), .B2(n_232), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_242), .B(n_229), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_240), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_262), .A2(n_227), .B1(n_173), .B2(n_190), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_251), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_241), .B(n_217), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_241), .Y(n_281) );
AO21x2_ASAP7_75t_L g282 ( .A1(n_247), .A2(n_105), .B(n_113), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_245), .B(n_225), .Y(n_283) );
OAI322xp33_ASAP7_75t_L g284 ( .A1(n_261), .A2(n_116), .A3(n_108), .B1(n_133), .B2(n_123), .C1(n_84), .C2(n_90), .Y(n_284) );
OAI221xp5_ASAP7_75t_L g285 ( .A1(n_237), .A2(n_191), .B1(n_206), .B2(n_231), .C(n_175), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_239), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_238), .B(n_225), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_238), .B(n_225), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_239), .B(n_198), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_281), .B(n_255), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_279), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_271), .A2(n_259), .B(n_251), .Y(n_293) );
BUFx2_ASAP7_75t_L g294 ( .A(n_276), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_281), .Y(n_295) );
BUFx12f_ASAP7_75t_L g296 ( .A(n_272), .Y(n_296) );
NOR2x1_ASAP7_75t_L g297 ( .A(n_276), .B(n_243), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_270), .B(n_255), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_286), .A2(n_252), .B1(n_250), .B2(n_244), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_282), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_268), .B(n_257), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_257), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_280), .Y(n_305) );
INVx2_ASAP7_75t_SL g306 ( .A(n_288), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_282), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_288), .B(n_258), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_282), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_283), .B(n_258), .Y(n_310) );
AND2x4_ASAP7_75t_L g311 ( .A(n_273), .B(n_251), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_287), .B(n_259), .Y(n_312) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_294), .B(n_259), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_295), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_308), .B(n_243), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_302), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_299), .B(n_244), .Y(n_319) );
INVx1_ASAP7_75t_SL g320 ( .A(n_291), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_308), .B(n_243), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_307), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_302), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_291), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_302), .Y(n_326) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_267), .B1(n_275), .B2(n_266), .C(n_272), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_309), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_303), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_309), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_308), .B(n_243), .Y(n_333) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_292), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_304), .B(n_248), .Y(n_335) );
NOR3xp33_ASAP7_75t_L g336 ( .A(n_299), .B(n_284), .C(n_92), .Y(n_336) );
OA21x2_ASAP7_75t_L g337 ( .A1(n_293), .A2(n_247), .B(n_260), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_294), .B(n_248), .Y(n_338) );
NAND4xp25_ASAP7_75t_SL g339 ( .A(n_300), .B(n_278), .C(n_272), .D(n_285), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_329), .B(n_304), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_320), .B(n_296), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_319), .B(n_305), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_325), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_330), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_331), .B(n_301), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_313), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_332), .B(n_305), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_318), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_314), .B(n_301), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_315), .B(n_304), .Y(n_352) );
NAND2x1_ASAP7_75t_L g353 ( .A(n_325), .B(n_297), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_339), .A2(n_327), .B1(n_296), .B2(n_336), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_314), .B(n_306), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_317), .B(n_306), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_317), .B(n_306), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_321), .B(n_310), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_316), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_322), .B(n_311), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_320), .B(n_298), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_316), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_321), .B(n_297), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_333), .B(n_311), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_310), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_339), .B(n_296), .Y(n_369) );
OR2x6_ASAP7_75t_L g370 ( .A(n_338), .B(n_272), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_340), .B(n_310), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_312), .Y(n_372) );
OR2x2_ASAP7_75t_L g373 ( .A(n_338), .B(n_290), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_318), .Y(n_374) );
INVxp67_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_335), .B(n_311), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_322), .B(n_312), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_323), .B(n_298), .Y(n_378) );
OAI33xp33_ASAP7_75t_L g379 ( .A1(n_323), .A2(n_290), .A3(n_123), .B1(n_133), .B2(n_269), .B3(n_289), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_328), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_328), .Y(n_381) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_330), .B(n_88), .C(n_91), .D(n_87), .Y(n_382) );
NAND4xp25_ASAP7_75t_L g383 ( .A(n_330), .B(n_91), .C(n_298), .D(n_253), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_318), .B(n_312), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_383), .A2(n_293), .B(n_326), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_348), .B(n_324), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_355), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_359), .B(n_324), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_372), .B(n_324), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_375), .B(n_326), .Y(n_390) );
NOR2x1_ASAP7_75t_R g391 ( .A(n_345), .B(n_231), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_370), .B(n_326), .Y(n_392) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_370), .B(n_311), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_360), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_363), .Y(n_395) );
NAND2xp67_ASAP7_75t_L g396 ( .A(n_377), .B(n_123), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_375), .B(n_311), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_380), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_381), .B(n_337), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_366), .B(n_337), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_357), .B(n_337), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_378), .B(n_337), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_358), .B(n_101), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
OR2x6_ASAP7_75t_L g405 ( .A(n_362), .B(n_248), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_368), .B(n_5), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_345), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_342), .B(n_248), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_376), .B(n_101), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_376), .B(n_7), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_364), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_367), .B(n_7), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_344), .B(n_8), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_371), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_347), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_367), .B(n_9), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_365), .B(n_10), .Y(n_417) );
NAND2x1p5_ASAP7_75t_L g418 ( .A(n_343), .B(n_231), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_352), .B(n_133), .Y(n_419) );
OAI21xp33_ASAP7_75t_SL g420 ( .A1(n_343), .A2(n_274), .B(n_260), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_362), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_344), .B(n_10), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_365), .B(n_12), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_369), .B(n_12), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_351), .B(n_13), .Y(n_425) );
NOR2x1p5_ASAP7_75t_SL g426 ( .A(n_346), .B(n_155), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_349), .Y(n_427) );
OR2x2_ASAP7_75t_L g428 ( .A(n_373), .B(n_14), .Y(n_428) );
INVxp67_ASAP7_75t_L g429 ( .A(n_370), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
NOR3xp33_ASAP7_75t_L g431 ( .A(n_382), .B(n_82), .C(n_110), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_356), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_346), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_374), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_361), .B(n_15), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_374), .B(n_15), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_424), .A2(n_369), .B1(n_354), .B2(n_361), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_389), .B(n_361), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_353), .B1(n_350), .B2(n_379), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_409), .B(n_350), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_350), .B1(n_122), .B2(n_16), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_404), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_388), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g444 ( .A1(n_422), .A2(n_17), .B(n_264), .C(n_161), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_433), .Y(n_446) );
AND3x1_ASAP7_75t_L g447 ( .A(n_413), .B(n_264), .C(n_122), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_427), .B(n_122), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_387), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_390), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_403), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_430), .B(n_249), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_395), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_414), .B(n_249), .Y(n_455) );
OAI22xp33_ASAP7_75t_L g456 ( .A1(n_405), .A2(n_212), .B1(n_230), .B2(n_198), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_415), .B(n_256), .Y(n_457) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_428), .A2(n_18), .B(n_20), .Y(n_458) );
INVxp67_ASAP7_75t_L g459 ( .A(n_386), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_410), .A2(n_256), .B(n_198), .Y(n_460) );
NAND2xp33_ASAP7_75t_SL g461 ( .A(n_393), .B(n_212), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_401), .B(n_24), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_432), .B(n_25), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_388), .B(n_429), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_398), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_420), .B(n_154), .C(n_159), .Y(n_466) );
OA21x2_ASAP7_75t_L g467 ( .A1(n_400), .A2(n_161), .B(n_156), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_397), .B(n_26), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_406), .B(n_28), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_434), .B(n_33), .Y(n_470) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_417), .A2(n_161), .B1(n_156), .B2(n_155), .C(n_159), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_423), .A2(n_156), .B1(n_155), .B2(n_159), .C(n_154), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_436), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_402), .B(n_35), .Y(n_474) );
OAI22xp5_ASAP7_75t_SL g475 ( .A1(n_421), .A2(n_212), .B1(n_198), .B2(n_185), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_400), .Y(n_476) );
OAI21xp5_ASAP7_75t_SL g477 ( .A1(n_421), .A2(n_212), .B(n_44), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_386), .B(n_38), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_399), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_419), .Y(n_480) );
INVxp67_ASAP7_75t_L g481 ( .A(n_399), .Y(n_481) );
AOI21xp33_ASAP7_75t_L g482 ( .A1(n_425), .A2(n_48), .B(n_49), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_402), .B(n_52), .Y(n_483) );
NAND2xp33_ASAP7_75t_SL g484 ( .A(n_443), .B(n_412), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g485 ( .A1(n_473), .A2(n_416), .B1(n_435), .B2(n_419), .C(n_385), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_449), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_453), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_437), .B(n_396), .Y(n_488) );
XNOR2xp5_ASAP7_75t_L g489 ( .A(n_464), .B(n_418), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_481), .A2(n_408), .B1(n_392), .B2(n_431), .C(n_418), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_451), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_454), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_461), .B(n_392), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_465), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_438), .B(n_405), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_442), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_477), .A2(n_405), .B(n_391), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_447), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_448), .Y(n_500) );
OAI221xp5_ASAP7_75t_L g501 ( .A1(n_459), .A2(n_481), .B1(n_444), .B2(n_461), .C(n_466), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_459), .B(n_426), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_476), .B(n_53), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_450), .B(n_55), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_479), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_439), .B(n_230), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_476), .B(n_56), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_446), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_479), .Y(n_509) );
OAI31xp33_ASAP7_75t_L g510 ( .A1(n_441), .A2(n_57), .A3(n_59), .B(n_61), .Y(n_510) );
OAI322xp33_ASAP7_75t_L g511 ( .A1(n_480), .A2(n_159), .A3(n_154), .B1(n_65), .B2(n_67), .C1(n_68), .C2(n_69), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g512 ( .A1(n_469), .A2(n_212), .B(n_64), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_446), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_450), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_455), .B(n_63), .Y(n_515) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_484), .A2(n_469), .B(n_458), .C(n_482), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_491), .A2(n_468), .B1(n_456), .B2(n_462), .Y(n_517) );
OAI21xp5_ASAP7_75t_SL g518 ( .A1(n_512), .A2(n_456), .B(n_478), .Y(n_518) );
AOI311xp33_ASAP7_75t_L g519 ( .A1(n_488), .A2(n_471), .A3(n_460), .B(n_472), .C(n_483), .Y(n_519) );
AOI21xp33_ASAP7_75t_SL g520 ( .A1(n_498), .A2(n_475), .B(n_467), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_484), .A2(n_474), .B(n_440), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_486), .Y(n_522) );
OAI21xp33_ASAP7_75t_L g523 ( .A1(n_488), .A2(n_457), .B(n_452), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_485), .B(n_467), .Y(n_524) );
CKINVDCx16_ASAP7_75t_R g525 ( .A(n_491), .Y(n_525) );
AOI211xp5_ASAP7_75t_L g526 ( .A1(n_499), .A2(n_463), .B(n_470), .C(n_467), .Y(n_526) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_501), .A2(n_70), .B(n_71), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_506), .A2(n_185), .B(n_198), .C(n_77), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_500), .B(n_154), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_490), .A2(n_154), .B1(n_159), .B2(n_502), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_495), .A2(n_154), .B1(n_159), .B2(n_508), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_510), .B(n_493), .C(n_497), .Y(n_532) );
AOI22x1_ASAP7_75t_L g533 ( .A1(n_489), .A2(n_508), .B1(n_504), .B2(n_514), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_505), .Y(n_534) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_520), .A2(n_487), .B1(n_492), .B2(n_494), .C(n_496), .Y(n_535) );
INVxp67_ASAP7_75t_L g536 ( .A(n_532), .Y(n_536) );
OAI21xp33_ASAP7_75t_SL g537 ( .A1(n_521), .A2(n_493), .B(n_504), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_517), .A2(n_505), .B1(n_509), .B2(n_513), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_522), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_517), .A2(n_509), .B1(n_515), .B2(n_503), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_534), .Y(n_541) );
INVx1_ASAP7_75t_SL g542 ( .A(n_525), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g543 ( .A(n_527), .B(n_511), .C(n_507), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_524), .B(n_523), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g545 ( .A1(n_530), .A2(n_516), .B(n_533), .C(n_518), .Y(n_545) );
OAI21x1_ASAP7_75t_SL g546 ( .A1(n_535), .A2(n_526), .B(n_531), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_539), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_542), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_538), .B(n_519), .Y(n_549) );
NOR2xp33_ASAP7_75t_SL g550 ( .A(n_537), .B(n_528), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_536), .B(n_529), .C(n_545), .Y(n_551) );
INVx3_ASAP7_75t_L g552 ( .A(n_548), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_547), .B(n_544), .Y(n_553) );
OR4x2_ASAP7_75t_L g554 ( .A(n_546), .B(n_540), .C(n_543), .D(n_541), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_552), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_552), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_555), .Y(n_557) );
OA22x2_ASAP7_75t_L g558 ( .A1(n_556), .A2(n_552), .B1(n_549), .B2(n_553), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_557), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g560 ( .A1(n_559), .A2(n_552), .B1(n_553), .B2(n_554), .C1(n_558), .C2(n_550), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_560), .A2(n_551), .B1(n_553), .B2(n_554), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_561), .A2(n_551), .B(n_553), .Y(n_562) );
endmodule