module fake_jpeg_6892_n_209 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_8),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_38),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_14),
.B1(n_12),
.B2(n_23),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_25),
.B1(n_24),
.B2(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_25),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_19),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_47),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_32),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_56),
.A2(n_57),
.B1(n_28),
.B2(n_30),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_36),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_32),
.Y(n_59)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_39),
.Y(n_70)
);

XOR2x2_ASAP7_75t_SL g87 ( 
.A(n_70),
.B(n_47),
.Y(n_87)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_28),
.B1(n_30),
.B2(n_55),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_80),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_54),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_73),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_51),
.B1(n_56),
.B2(n_45),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_84),
.B1(n_88),
.B2(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_71),
.B(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI21x1_ASAP7_75t_L g92 ( 
.A1(n_87),
.A2(n_63),
.B(n_54),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_56),
.B1(n_48),
.B2(n_29),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_48),
.B(n_54),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_69),
.B(n_63),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_77),
.A2(n_74),
.B1(n_71),
.B2(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_94),
.B1(n_105),
.B2(n_90),
.Y(n_112)
);

XOR2x1_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_87),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_63),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_101),
.C(n_81),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_103),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_85),
.B(n_67),
.C(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_33),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_110),
.B(n_19),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_88),
.B1(n_77),
.B2(n_84),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_108),
.A2(n_111),
.B1(n_122),
.B2(n_27),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_87),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_105),
.A2(n_88),
.B1(n_80),
.B2(n_81),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_38),
.B1(n_31),
.B2(n_27),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_68),
.B1(n_89),
.B2(n_62),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_119),
.B1(n_61),
.B2(n_72),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_94),
.C(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_101),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_120),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_68),
.B1(n_53),
.B2(n_64),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_86),
.B1(n_68),
.B2(n_78),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_137),
.C(n_138),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_128),
.B1(n_139),
.B2(n_22),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_93),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_127),
.B(n_132),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_103),
.B1(n_99),
.B2(n_104),
.Y(n_128)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_112),
.A2(n_64),
.B1(n_16),
.B2(n_22),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_64),
.B1(n_16),
.B2(n_22),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_72),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_121),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_115),
.Y(n_143)
);

XOR2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_61),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_136),
.B(n_19),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_64),
.C(n_27),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_27),
.C(n_31),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_27),
.C(n_31),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_31),
.C(n_65),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_121),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_117),
.B1(n_115),
.B2(n_122),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_144),
.A2(n_133),
.B(n_130),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_19),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_110),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_147),
.A2(n_151),
.B(n_138),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_140),
.C(n_137),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_132),
.Y(n_159)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_154),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_20),
.B1(n_21),
.B2(n_13),
.Y(n_155)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_155),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_161),
.B(n_162),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_164),
.Y(n_173)
);

NOR2xp67_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_123),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_167),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_145),
.B(n_134),
.Y(n_160)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_148),
.B(n_129),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_146),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_165),
.A2(n_152),
.B1(n_162),
.B2(n_166),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_21),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_176),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_177),
.B(n_174),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_163),
.A2(n_149),
.A3(n_142),
.B1(n_150),
.B2(n_65),
.C1(n_31),
.C2(n_21),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_159),
.B(n_142),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_179),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_181),
.B(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

AOI21x1_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_156),
.B(n_10),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_188),
.B(n_7),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_21),
.B(n_20),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_186),
.A2(n_65),
.B(n_20),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_187),
.Y(n_192)
);

AOI31xp33_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_8),
.A3(n_10),
.B(n_7),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_185),
.B(n_169),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_194),
.B(n_186),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_187),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_172),
.C(n_7),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_0),
.C(n_1),
.Y(n_201)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_196),
.A2(n_199),
.A3(n_200),
.B1(n_1),
.B2(n_4),
.C1(n_5),
.C2(n_40),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_15),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_201),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_192),
.A2(n_52),
.A3(n_15),
.B1(n_40),
.B2(n_3),
.C1(n_0),
.C2(n_5),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_52),
.B(n_40),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_199),
.A2(n_52),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_205),
.A2(n_4),
.B(n_5),
.Y(n_206)
);

OAI211xp5_ASAP7_75t_L g208 ( 
.A1(n_206),
.A2(n_202),
.B(n_4),
.C(n_5),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_207),
.Y(n_209)
);


endmodule