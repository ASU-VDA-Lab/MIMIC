module fake_ariane_3167_n_2055 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2055);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2055;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_363;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_1003;
wire n_701;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_1102;
wire n_719;
wire n_263;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_132),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_177),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_90),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_77),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_105),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_47),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_113),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_166),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_49),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_6),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_51),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_38),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_15),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_8),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_110),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_111),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_46),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_30),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_123),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_101),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_106),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_179),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_40),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_108),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_0),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_33),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_181),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_139),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_71),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_30),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_26),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_12),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_72),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_104),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_130),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_6),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_86),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_73),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_22),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_203),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_63),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_155),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_14),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_89),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_52),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_114),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_138),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_141),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_124),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_45),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_50),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_9),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_125),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_121),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_23),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_5),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_109),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_201),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_41),
.Y(n_277)
);

BUFx2_ASAP7_75t_SL g278 ( 
.A(n_41),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_22),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_87),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_163),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_9),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_100),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_159),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_84),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_39),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_128),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_53),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_147),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_92),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_129),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_98),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_133),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_117),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_78),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_127),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_99),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_185),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_198),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_172),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_17),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_171),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_205),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_26),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_192),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_75),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_103),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_10),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_173),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_93),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_8),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_169),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_19),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_74),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_44),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_42),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_49),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_152),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_33),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_11),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_34),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_20),
.Y(n_323)
);

CKINVDCx14_ASAP7_75t_R g324 ( 
.A(n_44),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_23),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_137),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_119),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_50),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_19),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_66),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_20),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_95),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_183),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_112),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_88),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_91),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_13),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_48),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_68),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_134),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_62),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_15),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_153),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_160),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_13),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_40),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_187),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_188),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_54),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_202),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_118),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_76),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_43),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_148),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_10),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_170),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_161),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_154),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_97),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_69),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_64),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_12),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_189),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_175),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_11),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_83),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_42),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_149),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_200),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_196),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_70),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_27),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_37),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_102),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_167),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_37),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_58),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_136),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_156),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_58),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_151),
.Y(n_381)
);

BUFx5_ASAP7_75t_L g382 ( 
.A(n_145),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_157),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_80),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_48),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_31),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_62),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_57),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_180),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_35),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_60),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_67),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_197),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_120),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_107),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_27),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_56),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_142),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_34),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_2),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_94),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_7),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_126),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_184),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_43),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_122),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_164),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_60),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_17),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_116),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_57),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_55),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_402),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_213),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_324),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_213),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_224),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_267),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_362),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_224),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_400),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_402),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_360),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_217),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_217),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_392),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_226),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_400),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_220),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_407),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_402),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_232),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_226),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_266),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_308),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_405),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_405),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_405),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_405),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_209),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_232),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_261),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_323),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_209),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_355),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_355),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_223),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_247),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_260),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_269),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_270),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_261),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_283),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_274),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_283),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_277),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_287),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_305),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_312),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_258),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_327),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_314),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_221),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_281),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_318),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g469 ( 
.A(n_317),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_325),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_281),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_377),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_329),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_327),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_346),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_373),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_332),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_288),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_221),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_385),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_377),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_386),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_253),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_250),
.Y(n_485)
);

INVxp67_ASAP7_75t_SL g486 ( 
.A(n_253),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_294),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_258),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_332),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_258),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_371),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_371),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_278),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_225),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_378),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_221),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_286),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_225),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_286),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_378),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_286),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_288),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_299),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_297),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_403),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_297),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_339),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_403),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_408),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_299),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_299),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_219),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_408),
.Y(n_514)
);

INVxp33_ASAP7_75t_SL g515 ( 
.A(n_228),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_304),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_304),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_304),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_334),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_339),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_422),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_487),
.B(n_291),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_413),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_433),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_413),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_432),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_432),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_435),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_455),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_455),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_444),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_433),
.B(n_291),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_435),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_424),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_438),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_439),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_440),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_441),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_441),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_486),
.B(n_481),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_464),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_485),
.A2(n_219),
.B1(n_268),
.B2(n_236),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_504),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_476),
.B(n_334),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_507),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_507),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_508),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

BUFx2_ASAP7_75t_L g556 ( 
.A(n_415),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_502),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_502),
.B(n_354),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_520),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_520),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_464),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_210),
.Y(n_562)
);

OAI21x1_ASAP7_75t_L g563 ( 
.A1(n_431),
.A2(n_294),
.B(n_212),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_444),
.B(n_294),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_485),
.A2(n_268),
.B1(n_337),
.B2(n_236),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_443),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_474),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g569 ( 
.A(n_419),
.B(n_256),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_425),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_467),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_490),
.B(n_272),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_447),
.Y(n_573)
);

OA21x2_ASAP7_75t_L g574 ( 
.A1(n_447),
.A2(n_218),
.B(n_211),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_414),
.B(n_334),
.Y(n_575)
);

AND2x6_ASAP7_75t_L g576 ( 
.A(n_467),
.B(n_254),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_497),
.B(n_222),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_448),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_448),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_416),
.B(n_228),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_471),
.B(n_354),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_427),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_449),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_449),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_472),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_417),
.B(n_230),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_472),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_499),
.B(n_271),
.Y(n_588)
);

INVxp33_ASAP7_75t_SL g589 ( 
.A(n_423),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_471),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_478),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_478),
.Y(n_592)
);

AND2x4_ASAP7_75t_L g593 ( 
.A(n_501),
.B(n_381),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_429),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_503),
.B(n_242),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_450),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_512),
.B(n_381),
.Y(n_597)
);

AND2x4_ASAP7_75t_L g598 ( 
.A(n_517),
.B(n_272),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_451),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_452),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_420),
.B(n_364),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_453),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_457),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_421),
.B(n_230),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_428),
.B(n_484),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_459),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_545),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_551),
.B(n_511),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_551),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_535),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_524),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_524),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_545),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_545),
.Y(n_616)
);

NAND3xp33_ASAP7_75t_L g617 ( 
.A(n_603),
.B(n_493),
.C(n_436),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_525),
.B(n_518),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_526),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_546),
.B(n_519),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_527),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_536),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_546),
.B(n_519),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_524),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_536),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_602),
.B(n_463),
.Y(n_627)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_564),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_524),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_564),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_557),
.B(n_437),
.Y(n_632)
);

AND2x6_ASAP7_75t_L g633 ( 
.A(n_575),
.B(n_254),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_537),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_537),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_526),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_539),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_525),
.B(n_423),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_557),
.B(n_511),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_575),
.B(n_516),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_522),
.B(n_516),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_524),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_526),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_539),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_602),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_524),
.Y(n_647)
);

INVx4_ASAP7_75t_L g648 ( 
.A(n_564),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_572),
.A2(n_515),
.B1(n_436),
.B2(n_498),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_522),
.B(n_426),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_541),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_541),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_522),
.B(n_426),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_522),
.B(n_430),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_528),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_528),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_602),
.B(n_430),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_533),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_542),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_530),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_R g662 ( 
.A(n_531),
.B(n_474),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_528),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_538),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_564),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_564),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_538),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_538),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_525),
.B(n_515),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_540),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_602),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_580),
.B(n_466),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_598),
.B(n_506),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_580),
.B(n_479),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_588),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_598),
.B(n_514),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_533),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_540),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_603),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_542),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_540),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_543),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_586),
.B(n_496),
.Y(n_684)
);

BUFx3_ASAP7_75t_L g685 ( 
.A(n_603),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_523),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_523),
.Y(n_687)
);

INVx11_ASAP7_75t_L g688 ( 
.A(n_564),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_554),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_554),
.Y(n_691)
);

INVxp33_ASAP7_75t_L g692 ( 
.A(n_569),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_583),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_586),
.B(n_510),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_590),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_590),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_R g699 ( 
.A(n_589),
.B(n_489),
.Y(n_699)
);

INVxp33_ASAP7_75t_L g700 ( 
.A(n_548),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_576),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_591),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_591),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_533),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_591),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_529),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_554),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_533),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_554),
.Y(n_709)
);

AO21x2_ASAP7_75t_L g710 ( 
.A1(n_563),
.A2(n_255),
.B(n_251),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_549),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_529),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_603),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_605),
.B(n_498),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_529),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_598),
.B(n_494),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_574),
.A2(n_469),
.B1(n_446),
.B2(n_418),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_548),
.A2(n_572),
.B1(n_396),
.B2(n_337),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_605),
.B(n_207),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_583),
.Y(n_720)
);

INVx5_ASAP7_75t_L g721 ( 
.A(n_576),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_547),
.Y(n_722)
);

BUFx10_ASAP7_75t_L g723 ( 
.A(n_598),
.Y(n_723)
);

NAND3xp33_ASAP7_75t_L g724 ( 
.A(n_603),
.B(n_276),
.C(n_263),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_529),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_572),
.B(n_460),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_549),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_561),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_529),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_572),
.B(n_461),
.Y(n_730)
);

OR2x6_ASAP7_75t_L g731 ( 
.A(n_572),
.B(n_462),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_534),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_558),
.B(n_465),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_593),
.B(n_468),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_583),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_534),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_534),
.Y(n_737)
);

BUFx3_ASAP7_75t_L g738 ( 
.A(n_603),
.Y(n_738)
);

INVx3_ASAP7_75t_L g739 ( 
.A(n_534),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_534),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_549),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_558),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_534),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_550),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_544),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_564),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_564),
.Y(n_747)
);

NAND3xp33_ASAP7_75t_L g748 ( 
.A(n_604),
.B(n_301),
.C(n_293),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_544),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_544),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_544),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_558),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_593),
.B(n_470),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_544),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_574),
.A2(n_388),
.B1(n_391),
.B2(n_475),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_558),
.B(n_473),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_621),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_655),
.B(n_692),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_723),
.B(n_556),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_610),
.B(n_593),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_610),
.B(n_593),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_726),
.B(n_597),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_730),
.B(n_597),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_627),
.B(n_597),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_627),
.B(n_597),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_621),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_611),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_628),
.A2(n_574),
.B1(n_396),
.B2(n_594),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_694),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_734),
.B(n_601),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_717),
.B(n_567),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_753),
.B(n_601),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_633),
.B(n_601),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_L g774 ( 
.A(n_744),
.B(n_604),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_633),
.B(n_618),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_633),
.B(n_601),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_622),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_633),
.B(n_562),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_L g779 ( 
.A(n_744),
.B(n_604),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_633),
.B(n_577),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_622),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_633),
.B(n_595),
.Y(n_782)
);

NAND3x1_ASAP7_75t_L g783 ( 
.A(n_718),
.B(n_513),
.C(n_445),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_SL g784 ( 
.A1(n_700),
.A2(n_456),
.B1(n_458),
.B2(n_434),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_623),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_686),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_646),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_653),
.B(n_604),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_687),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_723),
.B(n_604),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_661),
.B(n_489),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_623),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_633),
.B(n_659),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_654),
.B(n_599),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_608),
.A2(n_599),
.B(n_607),
.C(n_560),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_620),
.B(n_624),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_626),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_723),
.B(n_550),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_642),
.B(n_606),
.Y(n_799)
);

AO22x2_ASAP7_75t_L g800 ( 
.A1(n_649),
.A2(n_477),
.B1(n_495),
.B2(n_581),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_608),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_723),
.B(n_550),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_626),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_659),
.B(n_571),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_662),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_619),
.Y(n_806)
);

NAND3x1_ASAP7_75t_L g807 ( 
.A(n_673),
.B(n_492),
.C(n_491),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_678),
.B(n_571),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_731),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_678),
.B(n_571),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_661),
.B(n_491),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_704),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_722),
.B(n_571),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_617),
.B(n_500),
.C(n_492),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_731),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_704),
.B(n_581),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_634),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_676),
.B(n_550),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_676),
.B(n_609),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_619),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_636),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_676),
.B(n_560),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_708),
.B(n_581),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_634),
.Y(n_824)
);

NOR2x1p5_ASAP7_75t_L g825 ( 
.A(n_722),
.B(n_505),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_676),
.B(n_560),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_629),
.B(n_560),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_635),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_635),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_708),
.B(n_581),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_617),
.B(n_606),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_742),
.B(n_592),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_637),
.Y(n_833)
);

AOI22xp5_ASAP7_75t_L g834 ( 
.A1(n_731),
.A2(n_596),
.B1(n_600),
.B2(n_594),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_637),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_SL g836 ( 
.A(n_728),
.B(n_238),
.Y(n_836)
);

AND2x6_ASAP7_75t_L g837 ( 
.A(n_646),
.B(n_552),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_742),
.B(n_592),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_752),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_645),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_629),
.B(n_563),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_629),
.B(n_631),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_645),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_752),
.B(n_638),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_629),
.B(n_207),
.Y(n_845)
);

NOR2x1p5_ASAP7_75t_L g846 ( 
.A(n_728),
.B(n_505),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_658),
.A2(n_606),
.B1(n_509),
.B2(n_553),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_646),
.B(n_552),
.Y(n_848)
);

OR2x6_ASAP7_75t_L g849 ( 
.A(n_672),
.B(n_606),
.Y(n_849)
);

AND2x6_ASAP7_75t_SL g850 ( 
.A(n_716),
.B(n_480),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_694),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_641),
.B(n_553),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_677),
.B(n_509),
.Y(n_853)
);

BUFx4_ASAP7_75t_L g854 ( 
.A(n_699),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_639),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_671),
.B(n_555),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_636),
.Y(n_857)
);

OAI221xp5_ASAP7_75t_L g858 ( 
.A1(n_733),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.C(n_238),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_650),
.B(n_669),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_674),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_SL g861 ( 
.A(n_631),
.B(n_570),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_644),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_631),
.B(n_227),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_644),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_719),
.B(n_555),
.Y(n_865)
);

INVx5_ASAP7_75t_L g866 ( 
.A(n_631),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_671),
.B(n_559),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_651),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_671),
.B(n_566),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_755),
.B(n_566),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_684),
.B(n_584),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_714),
.Y(n_872)
);

NAND3xp33_ASAP7_75t_L g873 ( 
.A(n_696),
.B(n_409),
.C(n_240),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_711),
.A2(n_574),
.B1(n_583),
.B2(n_573),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_648),
.B(n_227),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_756),
.B(n_584),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_651),
.A2(n_240),
.B1(n_411),
.B2(n_412),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_656),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_652),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_652),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_648),
.B(n_231),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_727),
.B(n_585),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_657),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_727),
.B(n_587),
.Y(n_884)
);

AOI22xp5_ASAP7_75t_L g885 ( 
.A1(n_660),
.A2(n_364),
.B1(n_231),
.B2(n_233),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_741),
.B(n_587),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_657),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_694),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_694),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_660),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_741),
.A2(n_583),
.B1(n_573),
.B2(n_579),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_648),
.B(n_233),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_614),
.B(n_583),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_681),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_632),
.B(n_215),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_681),
.B(n_582),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_663),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_683),
.A2(n_579),
.B1(n_578),
.B2(n_573),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_648),
.B(n_234),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_665),
.B(n_234),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_665),
.B(n_235),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_683),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_693),
.A2(n_241),
.B1(n_239),
.B2(n_235),
.Y(n_903)
);

OAI21xp33_ASAP7_75t_L g904 ( 
.A1(n_693),
.A2(n_248),
.B(n_246),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_614),
.B(n_568),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_615),
.A2(n_579),
.B(n_578),
.C(n_568),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_615),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_616),
.B(n_568),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_612),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_616),
.B(n_482),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_663),
.A2(n_483),
.B(n_319),
.C(n_315),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_612),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_664),
.Y(n_913)
);

NOR2xp67_ASAP7_75t_L g914 ( 
.A(n_724),
.B(n_532),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_664),
.Y(n_915)
);

INVx5_ASAP7_75t_L g916 ( 
.A(n_837),
.Y(n_916)
);

INVxp67_ASAP7_75t_SL g917 ( 
.A(n_809),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_757),
.B(n_766),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_777),
.B(n_697),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_758),
.B(n_791),
.Y(n_920)
);

NOR3xp33_ASAP7_75t_L g921 ( 
.A(n_811),
.B(n_273),
.C(n_262),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_819),
.A2(n_859),
.B1(n_855),
.B2(n_796),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_801),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_837),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_781),
.B(n_697),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_785),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_792),
.B(n_797),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_809),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_815),
.B(n_665),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_767),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_803),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_817),
.B(n_824),
.Y(n_932)
);

BUFx3_ASAP7_75t_L g933 ( 
.A(n_896),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_819),
.A2(n_666),
.B1(n_746),
.B2(n_665),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_784),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_828),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_829),
.B(n_698),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_768),
.A2(n_667),
.B1(n_670),
.B2(n_668),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_833),
.B(n_698),
.Y(n_939)
);

BUFx6f_ASAP7_75t_L g940 ( 
.A(n_769),
.Y(n_940)
);

NOR2xp67_ASAP7_75t_L g941 ( 
.A(n_814),
.B(n_724),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_835),
.B(n_702),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_815),
.B(n_666),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_786),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_789),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_840),
.B(n_702),
.Y(n_946)
);

NAND2xp33_ASAP7_75t_SL g947 ( 
.A(n_805),
.B(n_666),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_759),
.B(n_612),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_843),
.B(n_703),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_868),
.B(n_703),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_759),
.B(n_612),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_831),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_879),
.B(n_705),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_853),
.B(n_705),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_880),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_849),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_825),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_762),
.B(n_694),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_837),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_859),
.B(n_613),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_806),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_890),
.B(n_667),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_849),
.B(n_666),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_894),
.B(n_668),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_820),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_854),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_771),
.B(n_670),
.Y(n_967)
);

OAI22xp33_ASAP7_75t_L g968 ( 
.A1(n_763),
.A2(n_282),
.B1(n_289),
.B2(n_279),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_902),
.B(n_679),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_768),
.A2(n_682),
.B1(n_679),
.B2(n_746),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_876),
.B(n_682),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_821),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_796),
.A2(n_747),
.B1(n_746),
.B2(n_685),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_769),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_836),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_910),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_850),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_893),
.A2(n_709),
.B(n_707),
.Y(n_978)
);

NOR3xp33_ASAP7_75t_SL g979 ( 
.A(n_858),
.B(n_309),
.C(n_302),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_837),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_860),
.B(n_613),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_876),
.B(n_707),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_872),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_872),
.B(n_613),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_844),
.B(n_839),
.Y(n_985)
);

NAND2x1p5_ASAP7_75t_L g986 ( 
.A(n_866),
.B(n_746),
.Y(n_986)
);

OR2x2_ASAP7_75t_L g987 ( 
.A(n_849),
.B(n_689),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_907),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_L g989 ( 
.A1(n_770),
.A2(n_709),
.B(n_647),
.C(n_750),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_813),
.B(n_839),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_846),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_847),
.B(n_720),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_882),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_884),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_886),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_800),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_832),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_895),
.B(n_625),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_838),
.Y(n_999)
);

OR2x6_ASAP7_75t_L g1000 ( 
.A(n_800),
.B(n_747),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_804),
.Y(n_1001)
);

AND2x2_ASAP7_75t_SL g1002 ( 
.A(n_861),
.B(n_747),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_831),
.A2(n_695),
.B(n_691),
.C(n_690),
.Y(n_1003)
);

AND3x1_ASAP7_75t_L g1004 ( 
.A(n_852),
.B(n_630),
.C(n_625),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_857),
.Y(n_1005)
);

CKINVDCx20_ASAP7_75t_R g1006 ( 
.A(n_877),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_794),
.B(n_316),
.Y(n_1007)
);

INVx1_ASAP7_75t_SL g1008 ( 
.A(n_783),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_866),
.B(n_720),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_764),
.B(n_625),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_808),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_862),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_810),
.Y(n_1013)
);

NAND2x1_ASAP7_75t_L g1014 ( 
.A(n_787),
.B(n_747),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_794),
.B(n_689),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_765),
.B(n_680),
.Y(n_1016)
);

OR2x2_ASAP7_75t_SL g1017 ( 
.A(n_873),
.B(n_748),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_SL g1018 ( 
.A(n_772),
.B(n_625),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_912),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_848),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_866),
.B(n_720),
.Y(n_1021)
);

AND3x2_ASAP7_75t_SL g1022 ( 
.A(n_807),
.B(n_691),
.C(n_690),
.Y(n_1022)
);

INVx5_ASAP7_75t_L g1023 ( 
.A(n_769),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_788),
.B(n_695),
.Y(n_1024)
);

AND3x1_ASAP7_75t_L g1025 ( 
.A(n_852),
.B(n_643),
.C(n_630),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_866),
.B(n_720),
.Y(n_1026)
);

INVxp67_ASAP7_75t_L g1027 ( 
.A(n_799),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_856),
.Y(n_1028)
);

AND2x6_ASAP7_75t_SL g1029 ( 
.A(n_871),
.B(n_306),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_864),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_867),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_760),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_841),
.A2(n_715),
.B(n_712),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_788),
.B(n_865),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_869),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_905),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_903),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_865),
.B(n_630),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_SL g1039 ( 
.A(n_871),
.B(n_640),
.Y(n_1039)
);

NOR2xp67_ASAP7_75t_L g1040 ( 
.A(n_885),
.B(n_748),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_878),
.B(n_643),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_883),
.B(n_643),
.Y(n_1042)
);

NAND2xp33_ASAP7_75t_SL g1043 ( 
.A(n_761),
.B(n_643),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_908),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_887),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_816),
.Y(n_1046)
);

INVx5_ASAP7_75t_L g1047 ( 
.A(n_769),
.Y(n_1047)
);

INVx4_ASAP7_75t_L g1048 ( 
.A(n_787),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_823),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_834),
.B(n_680),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_773),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_897),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_812),
.A2(n_685),
.B1(n_738),
.B2(n_713),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_830),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_913),
.B(n_647),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_915),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_909),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_851),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_904),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_795),
.Y(n_1060)
);

INVxp67_ASAP7_75t_SL g1061 ( 
.A(n_851),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_870),
.B(n_647),
.Y(n_1062)
);

INVx8_ASAP7_75t_L g1063 ( 
.A(n_851),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_776),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_851),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_827),
.B(n_647),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_889),
.Y(n_1067)
);

BUFx3_ASAP7_75t_L g1068 ( 
.A(n_889),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_906),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_889),
.Y(n_1070)
);

AND3x1_ASAP7_75t_SL g1071 ( 
.A(n_818),
.B(n_321),
.C(n_320),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_775),
.B(n_735),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_798),
.A2(n_680),
.B1(n_685),
.B2(n_713),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_889),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_778),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_780),
.Y(n_1076)
);

INVx2_ASAP7_75t_SL g1077 ( 
.A(n_818),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_798),
.B(n_713),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_SL g1079 ( 
.A(n_822),
.B(n_640),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_906),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_898),
.B(n_675),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_782),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_891),
.A2(n_845),
.B1(n_875),
.B2(n_863),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_793),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_898),
.B(n_675),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_822),
.B(n_706),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_790),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_826),
.B(n_735),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_888),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_790),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_891),
.A2(n_738),
.B1(n_710),
.B2(n_754),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_1063),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_1063),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_933),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_926),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_952),
.A2(n_826),
.B(n_802),
.C(n_901),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_SL g1097 ( 
.A(n_1037),
.B(n_328),
.C(n_322),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_922),
.B(n_802),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_952),
.A2(n_331),
.B1(n_399),
.B2(n_397),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1034),
.A2(n_874),
.B1(n_892),
.B2(n_901),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_923),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1063),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_929),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1034),
.A2(n_874),
.B1(n_881),
.B2(n_900),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1027),
.A2(n_875),
.B(n_863),
.C(n_900),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1007),
.B(n_845),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_971),
.A2(n_841),
.B(n_842),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_920),
.B(n_881),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_968),
.A2(n_911),
.B(n_779),
.C(n_774),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_931),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1027),
.B(n_892),
.Y(n_1111)
);

BUFx2_ASAP7_75t_R g1112 ( 
.A(n_935),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1032),
.B(n_899),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_936),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_971),
.A2(n_842),
.B(n_899),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_955),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1040),
.A2(n_911),
.B(n_738),
.C(n_706),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_993),
.A2(n_688),
.B1(n_706),
.B2(n_732),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_983),
.B(n_338),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_994),
.A2(n_732),
.B1(n_739),
.B2(n_750),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_976),
.B(n_732),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_916),
.B(n_739),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_918),
.A2(n_739),
.B1(n_750),
.B2(n_353),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_930),
.B(n_739),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_998),
.A2(n_989),
.B(n_1010),
.C(n_921),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_1006),
.B(n_1029),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1015),
.A2(n_982),
.B(n_1024),
.Y(n_1127)
);

NAND2x1p5_ASAP7_75t_L g1128 ( 
.A(n_916),
.B(n_640),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_956),
.B(n_341),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_928),
.Y(n_1130)
);

CKINVDCx6p67_ASAP7_75t_R g1131 ( 
.A(n_957),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_916),
.B(n_237),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_995),
.B(n_712),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_997),
.B(n_715),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_SL g1135 ( 
.A(n_959),
.B(n_914),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_916),
.B(n_237),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_960),
.A2(n_754),
.B(n_751),
.C(n_749),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1015),
.A2(n_710),
.B(n_725),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_924),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_940),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_924),
.B(n_239),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_966),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_929),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_928),
.B(n_975),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_917),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_956),
.B(n_342),
.Y(n_1146)
);

A2O1A1Ixp33_ASAP7_75t_SL g1147 ( 
.A1(n_989),
.A2(n_921),
.B(n_1060),
.C(n_951),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_924),
.B(n_241),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1033),
.A2(n_729),
.B(n_725),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_959),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_940),
.Y(n_1151)
);

INVx4_ASAP7_75t_L g1152 ( 
.A(n_924),
.Y(n_1152)
);

BUFx12f_ASAP7_75t_L g1153 ( 
.A(n_957),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_999),
.B(n_729),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_991),
.Y(n_1155)
);

NOR2xp67_ASAP7_75t_L g1156 ( 
.A(n_1023),
.B(n_736),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_954),
.B(n_737),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_944),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_990),
.B(n_737),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_977),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_917),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_1019),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_982),
.A2(n_710),
.B(n_740),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_985),
.B(n_743),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1024),
.A2(n_745),
.B(n_743),
.Y(n_1165)
);

AOI22x1_ASAP7_75t_L g1166 ( 
.A1(n_1048),
.A2(n_751),
.B1(n_749),
.B2(n_745),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_968),
.A2(n_404),
.B(n_395),
.C(n_311),
.Y(n_1167)
);

BUFx4f_ASAP7_75t_L g1168 ( 
.A(n_963),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1038),
.A2(n_978),
.B(n_925),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_967),
.B(n_345),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_945),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_940),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1000),
.B(n_349),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_918),
.A2(n_358),
.B(n_366),
.C(n_326),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_948),
.A2(n_344),
.B(n_369),
.C(n_359),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1000),
.B(n_365),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1038),
.A2(n_229),
.B(n_214),
.Y(n_1177)
);

AO21x1_ASAP7_75t_L g1178 ( 
.A1(n_1018),
.A2(n_343),
.B(n_357),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1000),
.B(n_367),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_978),
.A2(n_361),
.B(n_368),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_943),
.B(n_372),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_943),
.Y(n_1182)
);

BUFx6f_ASAP7_75t_L g1183 ( 
.A(n_974),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_927),
.A2(n_376),
.B1(n_380),
.B2(n_387),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1046),
.B(n_532),
.Y(n_1185)
);

INVx3_ASAP7_75t_SL g1186 ( 
.A(n_1059),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_974),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_988),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_961),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_965),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_963),
.Y(n_1191)
);

OAI21xp33_ASAP7_75t_L g1192 ( 
.A1(n_979),
.A2(n_244),
.B(n_208),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_979),
.A2(n_544),
.B(n_532),
.C(n_521),
.Y(n_1193)
);

AO32x2_ASAP7_75t_L g1194 ( 
.A1(n_1077),
.A2(n_521),
.A3(n_532),
.B1(n_576),
.B2(n_4),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_927),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_972),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_980),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1005),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_932),
.A2(n_532),
.B1(n_245),
.B2(n_330),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1071),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_974),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_932),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_919),
.A2(n_243),
.B(n_406),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1012),
.Y(n_1204)
);

AND2x4_ASAP7_75t_L g1205 ( 
.A(n_980),
.B(n_640),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_984),
.B(n_216),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1030),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_919),
.A2(n_937),
.B(n_925),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1045),
.Y(n_1209)
);

INVx3_ASAP7_75t_SL g1210 ( 
.A(n_1017),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1052),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1056),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1087),
.B(n_249),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1074),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1049),
.A2(n_532),
.B(n_521),
.C(n_336),
.Y(n_1215)
);

INVx5_ASAP7_75t_L g1216 ( 
.A(n_1074),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1020),
.A2(n_5),
.B(n_14),
.C(n_16),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_987),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_937),
.A2(n_335),
.B1(n_257),
.B2(n_259),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1079),
.A2(n_16),
.B(n_18),
.C(n_21),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_939),
.A2(n_252),
.B1(n_264),
.B2(n_275),
.Y(n_1221)
);

O2A1O1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1028),
.A2(n_18),
.B(n_21),
.C(n_24),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1050),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_939),
.A2(n_379),
.B1(n_300),
.B2(n_298),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1057),
.B(n_280),
.Y(n_1225)
);

A2O1A1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1054),
.A2(n_521),
.B(n_284),
.C(n_285),
.Y(n_1226)
);

INVx4_ASAP7_75t_L g1227 ( 
.A(n_1023),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_962),
.Y(n_1228)
);

AO32x2_ASAP7_75t_L g1229 ( 
.A1(n_1022),
.A2(n_521),
.A3(n_576),
.B1(n_28),
.B2(n_29),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_942),
.A2(n_389),
.B1(n_295),
.B2(n_292),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_1002),
.B(n_254),
.Y(n_1231)
);

INVxp67_ASAP7_75t_SL g1232 ( 
.A(n_1061),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1031),
.B(n_24),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1035),
.B(n_25),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_981),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1058),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1074),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1087),
.B(n_290),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1068),
.Y(n_1239)
);

INVx4_ASAP7_75t_L g1240 ( 
.A(n_1023),
.Y(n_1240)
);

OR2x6_ASAP7_75t_L g1241 ( 
.A(n_1050),
.B(n_521),
.Y(n_1241)
);

AO32x2_ASAP7_75t_L g1242 ( 
.A1(n_1100),
.A2(n_1022),
.A3(n_1070),
.B1(n_1051),
.B2(n_1064),
.Y(n_1242)
);

INVx3_ASAP7_75t_SL g1243 ( 
.A(n_1131),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1210),
.B(n_1008),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1195),
.A2(n_1231),
.B1(n_1208),
.B2(n_1106),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1127),
.A2(n_1061),
.B(n_946),
.Y(n_1246)
);

AOI221xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1217),
.A2(n_953),
.B1(n_946),
.B2(n_942),
.C(n_950),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1099),
.A2(n_1098),
.B1(n_1206),
.B2(n_1228),
.Y(n_1248)
);

AOI21xp33_ASAP7_75t_L g1249 ( 
.A1(n_1125),
.A2(n_1167),
.B(n_1174),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1160),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1130),
.B(n_996),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1144),
.B(n_1235),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1095),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1153),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1100),
.A2(n_1003),
.B(n_1081),
.Y(n_1255)
);

AOI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1138),
.A2(n_1072),
.B(n_958),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1149),
.A2(n_1080),
.B(n_1069),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1145),
.B(n_1001),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1169),
.A2(n_1062),
.B(n_1086),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1110),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1163),
.A2(n_1062),
.B(n_1086),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1107),
.A2(n_1088),
.B(n_1025),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1115),
.A2(n_950),
.B(n_949),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1103),
.B(n_1023),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1165),
.A2(n_1004),
.B(n_969),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1104),
.A2(n_949),
.B(n_953),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1104),
.A2(n_1043),
.B(n_962),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1214),
.Y(n_1268)
);

AO22x2_ASAP7_75t_L g1269 ( 
.A1(n_1173),
.A2(n_1011),
.B1(n_1013),
.B2(n_1075),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1166),
.A2(n_969),
.B(n_964),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1092),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1161),
.B(n_1036),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1108),
.B(n_1048),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1092),
.Y(n_1274)
);

BUFx3_ASAP7_75t_L g1275 ( 
.A(n_1162),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1186),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1119),
.B(n_1044),
.Y(n_1277)
);

OA21x2_ASAP7_75t_L g1278 ( 
.A1(n_1117),
.A2(n_1083),
.B(n_1091),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1094),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1175),
.A2(n_941),
.B(n_947),
.C(n_973),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1218),
.B(n_1076),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1223),
.B(n_1082),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1105),
.A2(n_1085),
.A3(n_1090),
.B(n_1089),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1118),
.A2(n_1042),
.B(n_1041),
.Y(n_1284)
);

OAI22x1_ASAP7_75t_L g1285 ( 
.A1(n_1126),
.A2(n_1071),
.B1(n_992),
.B2(n_1078),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1168),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1143),
.B(n_1067),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1092),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1178),
.A2(n_1055),
.A3(n_1041),
.B(n_1066),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1158),
.Y(n_1290)
);

AOI221x1_ASAP7_75t_L g1291 ( 
.A1(n_1193),
.A2(n_1096),
.B1(n_1192),
.B2(n_1123),
.C(n_1111),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1222),
.B(n_1016),
.C(n_1073),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1171),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1114),
.Y(n_1294)
);

NAND3x1_ASAP7_75t_L g1295 ( 
.A(n_1179),
.B(n_1067),
.C(n_1053),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1147),
.A2(n_1021),
.B(n_1009),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1112),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1143),
.B(n_1182),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1236),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1137),
.A2(n_1078),
.B(n_934),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1116),
.Y(n_1301)
);

AOI21xp33_ASAP7_75t_L g1302 ( 
.A1(n_1109),
.A2(n_1123),
.B(n_1202),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1220),
.A2(n_1026),
.B(n_1014),
.C(n_1065),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1170),
.B(n_938),
.Y(n_1304)
);

OAI221xp5_ASAP7_75t_L g1305 ( 
.A1(n_1099),
.A2(n_1097),
.B1(n_1192),
.B2(n_1181),
.C(n_1184),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1189),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1188),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1182),
.B(n_1047),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_SL g1309 ( 
.A1(n_1233),
.A2(n_1047),
.B(n_1070),
.C(n_1016),
.Y(n_1309)
);

AO32x2_ASAP7_75t_L g1310 ( 
.A1(n_1120),
.A2(n_1016),
.A3(n_970),
.B1(n_1047),
.B2(n_1084),
.Y(n_1310)
);

OAI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1234),
.A2(n_1215),
.B(n_1226),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1135),
.A2(n_1039),
.B(n_986),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_SL g1313 ( 
.A1(n_1122),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1191),
.B(n_986),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1133),
.A2(n_382),
.B(n_79),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1113),
.B(n_1129),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1177),
.A2(n_356),
.B(n_296),
.C(n_303),
.Y(n_1317)
);

O2A1O1Ixp33_ASAP7_75t_SL g1318 ( 
.A1(n_1132),
.A2(n_32),
.B(n_35),
.C(n_36),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1232),
.A2(n_254),
.B(n_265),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_SL g1320 ( 
.A1(n_1227),
.A2(n_32),
.B(n_36),
.Y(n_1320)
);

BUFx3_ASAP7_75t_L g1321 ( 
.A(n_1155),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1134),
.A2(n_576),
.B(n_310),
.Y(n_1322)
);

AND2x2_ASAP7_75t_SL g1323 ( 
.A(n_1168),
.B(n_265),
.Y(n_1323)
);

INVx6_ASAP7_75t_SL g1324 ( 
.A(n_1241),
.Y(n_1324)
);

CKINVDCx9p33_ASAP7_75t_R g1325 ( 
.A(n_1159),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1154),
.A2(n_1185),
.B(n_1197),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1150),
.B(n_374),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1200),
.A2(n_38),
.B1(n_39),
.B2(n_45),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1180),
.A2(n_1199),
.A3(n_1101),
.B(n_1196),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1207),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1199),
.A2(n_1141),
.B(n_1148),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1190),
.A2(n_382),
.A3(n_576),
.B(n_640),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1239),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1191),
.B(n_382),
.Y(n_1334)
);

NOR2xp67_ASAP7_75t_L g1335 ( 
.A(n_1214),
.B(n_194),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1128),
.A2(n_382),
.B(n_115),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1164),
.A2(n_370),
.B(n_313),
.Y(n_1337)
);

AOI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1136),
.A2(n_382),
.B(n_307),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1142),
.Y(n_1339)
);

NAND2x1p5_ASAP7_75t_L g1340 ( 
.A(n_1150),
.B(n_721),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1211),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1139),
.A2(n_265),
.B(n_307),
.Y(n_1342)
);

NAND2xp33_ASAP7_75t_L g1343 ( 
.A(n_1093),
.B(n_382),
.Y(n_1343)
);

INVxp67_ASAP7_75t_SL g1344 ( 
.A(n_1157),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1219),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_1345)
);

OAI21xp33_ASAP7_75t_L g1346 ( 
.A1(n_1219),
.A2(n_383),
.B(n_333),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1203),
.A2(n_375),
.B(n_340),
.C(n_347),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1236),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1152),
.A2(n_307),
.B(n_410),
.Y(n_1349)
);

O2A1O1Ixp33_ASAP7_75t_SL g1350 ( 
.A1(n_1213),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_1350)
);

A2O1A1Ixp33_ASAP7_75t_L g1351 ( 
.A1(n_1225),
.A2(n_384),
.B(n_348),
.C(n_350),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1152),
.A2(n_307),
.B(n_410),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1093),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1221),
.A2(n_59),
.B1(n_61),
.B2(n_410),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1221),
.A2(n_394),
.B(n_352),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1198),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_SL g1357 ( 
.A1(n_1238),
.A2(n_410),
.B(n_351),
.C(n_398),
.Y(n_1357)
);

AOI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1156),
.A2(n_410),
.B(n_701),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1224),
.A2(n_59),
.B(n_61),
.C(n_401),
.Y(n_1359)
);

OR2x2_ASAP7_75t_L g1360 ( 
.A(n_1176),
.B(n_393),
.Y(n_1360)
);

NOR2xp67_ASAP7_75t_L g1361 ( 
.A(n_1214),
.B(n_65),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1241),
.A2(n_363),
.B(n_721),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1216),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1241),
.A2(n_721),
.B(n_701),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1204),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1124),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1224),
.A2(n_721),
.B(n_701),
.Y(n_1367)
);

BUFx2_ASAP7_75t_L g1368 ( 
.A(n_1146),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1216),
.B(n_81),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1230),
.A2(n_721),
.B(n_701),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1230),
.A2(n_701),
.B1(n_85),
.B2(n_96),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1093),
.B(n_82),
.Y(n_1372)
);

NOR2xp67_ASAP7_75t_L g1373 ( 
.A(n_1240),
.B(n_140),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1102),
.B(n_143),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1121),
.A2(n_146),
.B(n_150),
.Y(n_1375)
);

AO31x2_ASAP7_75t_L g1376 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1229),
.B(n_1194),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_1102),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1102),
.A2(n_158),
.B1(n_162),
.B2(n_165),
.Y(n_1378)
);

INVx4_ASAP7_75t_L g1379 ( 
.A(n_1227),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1240),
.A2(n_174),
.B1(n_178),
.B2(n_186),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1140),
.A2(n_190),
.B(n_191),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1194),
.A2(n_204),
.B(n_1229),
.Y(n_1382)
);

NAND2x1p5_ASAP7_75t_L g1383 ( 
.A(n_1140),
.B(n_1151),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1140),
.B(n_1151),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1151),
.B(n_1172),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1172),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1172),
.B(n_1183),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1237),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1183),
.B(n_1187),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1183),
.Y(n_1390)
);

BUFx8_ASAP7_75t_L g1391 ( 
.A(n_1229),
.Y(n_1391)
);

AOI221x1_ASAP7_75t_L g1392 ( 
.A1(n_1187),
.A2(n_1201),
.B1(n_1237),
.B2(n_1194),
.C(n_1205),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1187),
.B(n_1201),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1201),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1237),
.A2(n_1195),
.B1(n_922),
.B2(n_1231),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1205),
.A2(n_1149),
.B(n_1033),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1127),
.A2(n_1208),
.B(n_1034),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1195),
.B(n_922),
.Y(n_1398)
);

AO21x2_ASAP7_75t_L g1399 ( 
.A1(n_1138),
.A2(n_1163),
.B(n_1127),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1286),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1339),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1261),
.A2(n_1246),
.B(n_1257),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1286),
.Y(n_1404)
);

OAI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1248),
.A2(n_1302),
.B(n_1266),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1377),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_SL g1407 ( 
.A1(n_1248),
.A2(n_1359),
.B(n_1398),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1252),
.B(n_1279),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1354),
.A2(n_1305),
.B1(n_1328),
.B2(n_1323),
.Y(n_1409)
);

INVxp67_ASAP7_75t_L g1410 ( 
.A(n_1366),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1392),
.A2(n_1291),
.A3(n_1397),
.B(n_1245),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1253),
.Y(n_1412)
);

INVx8_ASAP7_75t_L g1413 ( 
.A(n_1372),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1260),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1251),
.B(n_1368),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1396),
.A2(n_1263),
.B(n_1265),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1294),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1275),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1391),
.A2(n_1328),
.B1(n_1382),
.B2(n_1395),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1267),
.A2(n_1312),
.B(n_1399),
.Y(n_1420)
);

BUFx2_ASAP7_75t_L g1421 ( 
.A(n_1279),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1285),
.A2(n_1296),
.A3(n_1280),
.B(n_1319),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1273),
.B(n_1269),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1301),
.Y(n_1424)
);

OR2x6_ASAP7_75t_L g1425 ( 
.A(n_1295),
.B(n_1269),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1297),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1307),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1277),
.B(n_1316),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1255),
.A2(n_1247),
.B(n_1262),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1354),
.A2(n_1345),
.B1(n_1371),
.B2(n_1249),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_SL g1431 ( 
.A1(n_1345),
.A2(n_1249),
.B(n_1347),
.C(n_1327),
.Y(n_1431)
);

INVx6_ASAP7_75t_L g1432 ( 
.A(n_1377),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1371),
.A2(n_1304),
.B1(n_1302),
.B2(n_1292),
.Y(n_1433)
);

BUFx2_ASAP7_75t_L g1434 ( 
.A(n_1299),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1330),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1270),
.A2(n_1315),
.B(n_1284),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1272),
.B(n_1344),
.Y(n_1437)
);

NOR2xp67_ASAP7_75t_L g1438 ( 
.A(n_1333),
.B(n_1348),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1341),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1244),
.B(n_1360),
.Y(n_1440)
);

AOI21xp33_ASAP7_75t_L g1441 ( 
.A1(n_1247),
.A2(n_1391),
.B(n_1255),
.Y(n_1441)
);

INVx3_ASAP7_75t_SL g1442 ( 
.A(n_1254),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1290),
.Y(n_1443)
);

AOI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1370),
.A2(n_1338),
.B(n_1331),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1358),
.A2(n_1336),
.B(n_1300),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1293),
.Y(n_1446)
);

BUFx16f_ASAP7_75t_R g1447 ( 
.A(n_1372),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1342),
.A2(n_1349),
.B(n_1311),
.Y(n_1448)
);

NOR2xp67_ASAP7_75t_L g1449 ( 
.A(n_1268),
.B(n_1363),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1306),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1356),
.Y(n_1451)
);

INVx8_ASAP7_75t_L g1452 ( 
.A(n_1271),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1292),
.A2(n_1258),
.B1(n_1375),
.B2(n_1380),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1365),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1394),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1346),
.A2(n_1355),
.B(n_1317),
.C(n_1351),
.Y(n_1456)
);

AOI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1337),
.A2(n_1334),
.B(n_1278),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1314),
.A2(n_1357),
.B(n_1367),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1282),
.B(n_1281),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1367),
.A2(n_1381),
.B(n_1322),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1346),
.A2(n_1355),
.B1(n_1337),
.B2(n_1324),
.Y(n_1461)
);

BUFx2_ASAP7_75t_L g1462 ( 
.A(n_1353),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1321),
.B(n_1276),
.Y(n_1463)
);

AND2x4_ASAP7_75t_L g1464 ( 
.A(n_1268),
.B(n_1363),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1287),
.A2(n_1380),
.B(n_1389),
.Y(n_1465)
);

OAI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1298),
.A2(n_1324),
.B1(n_1308),
.B2(n_1378),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1383),
.A2(n_1364),
.B(n_1352),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1243),
.B(n_1288),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1320),
.A2(n_1388),
.B1(n_1386),
.B2(n_1390),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1379),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1325),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1376),
.B(n_1384),
.Y(n_1472)
);

CKINVDCx6p67_ASAP7_75t_R g1473 ( 
.A(n_1271),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1376),
.B(n_1283),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1309),
.A2(n_1303),
.B(n_1343),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1399),
.A2(n_1374),
.B1(n_1274),
.B2(n_1288),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1379),
.A2(n_1393),
.B1(n_1387),
.B2(n_1385),
.Y(n_1477)
);

AO22x2_ASAP7_75t_L g1478 ( 
.A1(n_1242),
.A2(n_1310),
.B1(n_1283),
.B2(n_1289),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1329),
.B(n_1289),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1350),
.B(n_1313),
.C(n_1318),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1274),
.B(n_1335),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1373),
.A2(n_1340),
.B(n_1362),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1340),
.A2(n_1361),
.B(n_1369),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1329),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1329),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1310),
.Y(n_1486)
);

INVx6_ASAP7_75t_L g1487 ( 
.A(n_1310),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1242),
.A2(n_1248),
.B1(n_1231),
.B2(n_1210),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1332),
.B(n_1398),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1332),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1279),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1248),
.B(n_1359),
.C(n_1345),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1297),
.Y(n_1493)
);

NAND3xp33_ASAP7_75t_L g1494 ( 
.A(n_1248),
.B(n_1359),
.C(n_1345),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1253),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1275),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1283),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1253),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1251),
.B(n_1252),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1253),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1391),
.A2(n_1000),
.B1(n_800),
.B2(n_996),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1253),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1253),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1251),
.B(n_1252),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1253),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1253),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1398),
.B(n_1195),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1253),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1328),
.A2(n_1006),
.B1(n_1126),
.B2(n_1200),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1398),
.B(n_1195),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1253),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1252),
.B(n_661),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1397),
.A2(n_1266),
.B(n_1208),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1398),
.B(n_1195),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1248),
.B(n_1273),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1286),
.B(n_1264),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1321),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1397),
.A2(n_1266),
.B(n_1208),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1522)
);

INVx5_ASAP7_75t_L g1523 ( 
.A(n_1286),
.Y(n_1523)
);

AO31x2_ASAP7_75t_L g1524 ( 
.A1(n_1392),
.A2(n_1291),
.A3(n_1266),
.B(n_1397),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1295),
.B(n_1241),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1253),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1321),
.Y(n_1529)
);

AOI21xp33_ASAP7_75t_L g1530 ( 
.A1(n_1248),
.A2(n_1247),
.B(n_1231),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1531)
);

OAI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1248),
.A2(n_1302),
.B(n_1266),
.Y(n_1532)
);

OAI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1328),
.A2(n_628),
.B1(n_1210),
.B2(n_922),
.Y(n_1533)
);

AND2x4_ASAP7_75t_L g1534 ( 
.A(n_1286),
.B(n_1264),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1251),
.B(n_1252),
.Y(n_1535)
);

INVxp67_ASAP7_75t_SL g1536 ( 
.A(n_1261),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1253),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1539)
);

OAI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1248),
.A2(n_1302),
.B(n_1266),
.Y(n_1540)
);

OR2x6_ASAP7_75t_L g1541 ( 
.A(n_1295),
.B(n_1241),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_SL g1542 ( 
.A1(n_1328),
.A2(n_1006),
.B1(n_1126),
.B2(n_1200),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_1250),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1253),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1256),
.A2(n_1326),
.B(n_1259),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1286),
.B(n_1264),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1286),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1253),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1248),
.A2(n_1328),
.B(n_1249),
.C(n_1345),
.Y(n_1549)
);

OA21x2_ASAP7_75t_L g1550 ( 
.A1(n_1420),
.A2(n_1532),
.B(n_1405),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1437),
.B(n_1509),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1518),
.B(n_1466),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1492),
.A2(n_1494),
.B1(n_1549),
.B2(n_1409),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1412),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1492),
.A2(n_1494),
.B1(n_1549),
.B2(n_1409),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1556)
);

CKINVDCx16_ASAP7_75t_R g1557 ( 
.A(n_1543),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1410),
.Y(n_1558)
);

O2A1O1Ixp33_ASAP7_75t_L g1559 ( 
.A1(n_1533),
.A2(n_1456),
.B(n_1407),
.C(n_1430),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1529),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_L g1561 ( 
.A1(n_1405),
.A2(n_1532),
.B(n_1540),
.C(n_1530),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1410),
.B(n_1535),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1509),
.B(n_1512),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1434),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1415),
.B(n_1491),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1425),
.B(n_1421),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1418),
.Y(n_1567)
);

AOI221x1_ASAP7_75t_SL g1568 ( 
.A1(n_1430),
.A2(n_1514),
.B1(n_1530),
.B2(n_1441),
.C(n_1408),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1401),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1419),
.A2(n_1540),
.B1(n_1433),
.B2(n_1453),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1428),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1414),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1511),
.A2(n_1542),
.B1(n_1488),
.B2(n_1419),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1455),
.Y(n_1574)
);

NOR2xp67_ASAP7_75t_L g1575 ( 
.A(n_1423),
.B(n_1520),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1431),
.A2(n_1433),
.B(n_1441),
.C(n_1488),
.Y(n_1576)
);

OAI31xp33_ASAP7_75t_L g1577 ( 
.A1(n_1466),
.A2(n_1501),
.A3(n_1480),
.B(n_1461),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1512),
.B(n_1516),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1417),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1401),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1496),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1459),
.B(n_1423),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1436),
.A2(n_1416),
.B(n_1402),
.Y(n_1583)
);

NOR2xp67_ASAP7_75t_L g1584 ( 
.A(n_1468),
.B(n_1477),
.Y(n_1584)
);

O2A1O1Ixp33_ASAP7_75t_L g1585 ( 
.A1(n_1480),
.A2(n_1516),
.B(n_1455),
.C(n_1477),
.Y(n_1585)
);

O2A1O1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1475),
.A2(n_1400),
.B(n_1404),
.C(n_1547),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1504),
.A2(n_1527),
.B(n_1517),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1440),
.B(n_1424),
.Y(n_1588)
);

NAND2x1p5_ASAP7_75t_L g1589 ( 
.A(n_1523),
.B(n_1465),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1463),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1486),
.A2(n_1471),
.B1(n_1487),
.B2(n_1413),
.Y(n_1591)
);

BUFx3_ASAP7_75t_L g1592 ( 
.A(n_1462),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1506),
.A2(n_1531),
.B(n_1545),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1427),
.B(n_1495),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_L g1595 ( 
.A1(n_1498),
.A2(n_1538),
.B(n_1548),
.C(n_1507),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1472),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1500),
.B(n_1502),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1503),
.B(n_1508),
.Y(n_1598)
);

OAI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1487),
.A2(n_1413),
.B1(n_1429),
.B2(n_1447),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1510),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1536),
.A2(n_1460),
.B(n_1429),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1513),
.B(n_1526),
.Y(n_1602)
);

O2A1O1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1544),
.A2(n_1469),
.B(n_1439),
.C(n_1435),
.Y(n_1603)
);

O2A1O1Ixp5_ASAP7_75t_L g1604 ( 
.A1(n_1489),
.A2(n_1457),
.B(n_1479),
.C(n_1470),
.Y(n_1604)
);

OAI22xp5_ASAP7_75t_L g1605 ( 
.A1(n_1487),
.A2(n_1447),
.B1(n_1523),
.B2(n_1525),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1523),
.A2(n_1541),
.B1(n_1476),
.B2(n_1470),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1523),
.A2(n_1541),
.B1(n_1406),
.B2(n_1432),
.Y(n_1607)
);

O2A1O1Ixp5_ASAP7_75t_L g1608 ( 
.A1(n_1479),
.A2(n_1481),
.B(n_1474),
.C(n_1444),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1519),
.B(n_1534),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1519),
.B(n_1546),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1442),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1449),
.A2(n_1426),
.B(n_1493),
.Y(n_1612)
);

O2A1O1Ixp5_ASAP7_75t_L g1613 ( 
.A1(n_1484),
.A2(n_1490),
.B(n_1485),
.C(n_1497),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1478),
.B(n_1411),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1473),
.B(n_1451),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1443),
.B(n_1446),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1450),
.B(n_1454),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1406),
.A2(n_1432),
.B1(n_1478),
.B2(n_1452),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1406),
.A2(n_1432),
.B1(n_1478),
.B2(n_1452),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1452),
.A2(n_1524),
.B1(n_1411),
.B2(n_1422),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1411),
.B(n_1524),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1448),
.A2(n_1458),
.B1(n_1445),
.B2(n_1482),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1522),
.A2(n_1528),
.B(n_1537),
.C(n_1539),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1403),
.B(n_1483),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1467),
.A2(n_1492),
.B1(n_1494),
.B2(n_1549),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1410),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1409),
.A2(n_1549),
.B(n_1453),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1420),
.A2(n_1392),
.B(n_1405),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1412),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1631)
);

BUFx2_ASAP7_75t_L g1632 ( 
.A(n_1421),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1420),
.A2(n_1392),
.B(n_1405),
.Y(n_1633)
);

OA21x2_ASAP7_75t_L g1634 ( 
.A1(n_1420),
.A2(n_1392),
.B(n_1405),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1491),
.B(n_1438),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1464),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1437),
.B(n_1509),
.Y(n_1637)
);

INVxp67_ASAP7_75t_L g1638 ( 
.A(n_1408),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1409),
.A2(n_1549),
.B(n_1453),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1409),
.A2(n_1549),
.B(n_1453),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1409),
.A2(n_1549),
.B(n_1453),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1412),
.Y(n_1642)
);

O2A1O1Ixp5_ASAP7_75t_L g1643 ( 
.A1(n_1409),
.A2(n_1530),
.B(n_1532),
.C(n_1405),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1492),
.A2(n_1494),
.B1(n_1549),
.B2(n_1409),
.Y(n_1644)
);

O2A1O1Ixp5_ASAP7_75t_L g1645 ( 
.A1(n_1409),
.A2(n_1530),
.B(n_1532),
.C(n_1405),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1412),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1410),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1410),
.Y(n_1648)
);

BUFx12f_ASAP7_75t_L g1649 ( 
.A(n_1426),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1650)
);

AOI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1409),
.A2(n_1328),
.B(n_1549),
.C(n_1533),
.Y(n_1651)
);

O2A1O1Ixp5_ASAP7_75t_L g1652 ( 
.A1(n_1409),
.A2(n_1530),
.B(n_1532),
.C(n_1405),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1549),
.A2(n_1494),
.B(n_1492),
.C(n_1409),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1491),
.B(n_1438),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1409),
.A2(n_1549),
.B(n_1453),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1499),
.B(n_1505),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1409),
.A2(n_1391),
.B1(n_1000),
.B2(n_800),
.Y(n_1657)
);

AOI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1515),
.A2(n_1521),
.B(n_1453),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1515),
.A2(n_1521),
.B(n_1453),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1492),
.A2(n_1494),
.B1(n_1549),
.B2(n_1409),
.Y(n_1660)
);

O2A1O1Ixp33_ASAP7_75t_L g1661 ( 
.A1(n_1533),
.A2(n_1549),
.B(n_1409),
.C(n_1456),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1437),
.B(n_1509),
.Y(n_1662)
);

OA21x2_ASAP7_75t_L g1663 ( 
.A1(n_1420),
.A2(n_1392),
.B(n_1405),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1437),
.B(n_1509),
.Y(n_1664)
);

OA21x2_ASAP7_75t_L g1665 ( 
.A1(n_1420),
.A2(n_1392),
.B(n_1405),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1409),
.A2(n_1549),
.B(n_1453),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1550),
.B(n_1629),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1657),
.A2(n_1570),
.B1(n_1573),
.B2(n_1660),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1554),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1550),
.B(n_1629),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1592),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1614),
.B(n_1621),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1600),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1558),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1572),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1579),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_SL g1677 ( 
.A1(n_1661),
.A2(n_1559),
.B(n_1570),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1633),
.B(n_1634),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1553),
.A2(n_1555),
.B1(n_1644),
.B2(n_1660),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1626),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1551),
.B(n_1637),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1647),
.Y(n_1682)
);

OAI21xp5_ASAP7_75t_L g1683 ( 
.A1(n_1627),
.A2(n_1640),
.B(n_1639),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1552),
.A2(n_1555),
.B1(n_1553),
.B2(n_1644),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1551),
.B(n_1662),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1633),
.B(n_1634),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1630),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1642),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1648),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1574),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1665),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1663),
.B(n_1665),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1563),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1577),
.A2(n_1625),
.B1(n_1651),
.B2(n_1638),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1658),
.B(n_1659),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1614),
.B(n_1565),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1564),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1646),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1595),
.Y(n_1699)
);

BUFx2_ASAP7_75t_L g1700 ( 
.A(n_1589),
.Y(n_1700)
);

AO21x2_ASAP7_75t_L g1701 ( 
.A1(n_1601),
.A2(n_1620),
.B(n_1561),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1613),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1583),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1598),
.B(n_1588),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1587),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1587),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1594),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1624),
.B(n_1636),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1596),
.B(n_1582),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1653),
.A2(n_1576),
.B(n_1585),
.Y(n_1710)
);

INVxp67_ASAP7_75t_R g1711 ( 
.A(n_1599),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1593),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1597),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1593),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1602),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1604),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1563),
.Y(n_1717)
);

AO21x2_ASAP7_75t_L g1718 ( 
.A1(n_1622),
.A2(n_1666),
.B(n_1641),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1608),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1578),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1632),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1581),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1655),
.B(n_1606),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1556),
.B(n_1628),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_R g1725 ( 
.A(n_1557),
.B(n_1649),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1575),
.A2(n_1617),
.B1(n_1566),
.B2(n_1591),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1578),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1643),
.A2(n_1652),
.B(n_1645),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1616),
.Y(n_1729)
);

OA21x2_ASAP7_75t_L g1730 ( 
.A1(n_1618),
.A2(n_1619),
.B(n_1606),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1603),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1618),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1567),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1623),
.Y(n_1734)
);

INVxp67_ASAP7_75t_L g1735 ( 
.A(n_1719),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1704),
.B(n_1631),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1667),
.B(n_1650),
.Y(n_1737)
);

OAI221xp5_ASAP7_75t_SL g1738 ( 
.A1(n_1679),
.A2(n_1668),
.B1(n_1677),
.B2(n_1694),
.C(n_1710),
.Y(n_1738)
);

INVxp67_ASAP7_75t_SL g1739 ( 
.A(n_1667),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1717),
.B(n_1568),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1717),
.B(n_1568),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1704),
.B(n_1656),
.Y(n_1742)
);

OAI21xp33_ASAP7_75t_L g1743 ( 
.A1(n_1679),
.A2(n_1562),
.B(n_1567),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1709),
.B(n_1571),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1669),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1704),
.B(n_1584),
.Y(n_1746)
);

NOR2x1_ASAP7_75t_SL g1747 ( 
.A(n_1723),
.B(n_1607),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1696),
.B(n_1591),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1673),
.Y(n_1749)
);

INVx3_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

NAND2x1_ASAP7_75t_L g1751 ( 
.A(n_1723),
.B(n_1654),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1720),
.B(n_1635),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1673),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1709),
.B(n_1560),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1709),
.B(n_1605),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1669),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1720),
.B(n_1586),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1727),
.B(n_1615),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1675),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1674),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1670),
.B(n_1610),
.Y(n_1761)
);

NAND2x1p5_ASAP7_75t_L g1762 ( 
.A(n_1728),
.B(n_1700),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1676),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1724),
.B(n_1609),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1671),
.B(n_1611),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1727),
.B(n_1590),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1678),
.B(n_1686),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1678),
.B(n_1569),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1678),
.B(n_1580),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1708),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1705),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1708),
.B(n_1612),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1745),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1740),
.A2(n_1683),
.B1(n_1668),
.B2(n_1718),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1745),
.Y(n_1775)
);

BUFx2_ASAP7_75t_L g1776 ( 
.A(n_1768),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1767),
.B(n_1722),
.Y(n_1777)
);

OAI33xp33_ASAP7_75t_L g1778 ( 
.A1(n_1740),
.A2(n_1684),
.A3(n_1685),
.B1(n_1681),
.B2(n_1693),
.B3(n_1715),
.Y(n_1778)
);

AOI221xp5_ASAP7_75t_L g1779 ( 
.A1(n_1741),
.A2(n_1684),
.B1(n_1694),
.B2(n_1699),
.C(n_1731),
.Y(n_1779)
);

OAI21x1_ASAP7_75t_L g1780 ( 
.A1(n_1762),
.A2(n_1712),
.B(n_1703),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1768),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1749),
.B(n_1672),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1749),
.B(n_1674),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1753),
.B(n_1680),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1767),
.B(n_1722),
.Y(n_1785)
);

AO21x2_ASAP7_75t_L g1786 ( 
.A1(n_1735),
.A2(n_1686),
.B(n_1691),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1760),
.Y(n_1787)
);

AO21x1_ASAP7_75t_SL g1788 ( 
.A1(n_1757),
.A2(n_1734),
.B(n_1683),
.Y(n_1788)
);

OAI33xp33_ASAP7_75t_L g1789 ( 
.A1(n_1741),
.A2(n_1685),
.A3(n_1681),
.B1(n_1693),
.B2(n_1715),
.B3(n_1713),
.Y(n_1789)
);

NAND2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1751),
.B(n_1725),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1737),
.B(n_1733),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1766),
.B(n_1733),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1769),
.A2(n_1718),
.B1(n_1723),
.B2(n_1731),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1756),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1738),
.A2(n_1699),
.B1(n_1723),
.B2(n_1726),
.C(n_1728),
.Y(n_1795)
);

NAND2xp33_ASAP7_75t_R g1796 ( 
.A(n_1772),
.B(n_1730),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1760),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1738),
.A2(n_1691),
.B1(n_1686),
.B2(n_1692),
.C(n_1719),
.Y(n_1798)
);

OAI221xp5_ASAP7_75t_L g1799 ( 
.A1(n_1735),
.A2(n_1723),
.B1(n_1728),
.B2(n_1719),
.C(n_1702),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1753),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1744),
.B(n_1680),
.Y(n_1801)
);

NAND2xp33_ASAP7_75t_R g1802 ( 
.A(n_1772),
.B(n_1730),
.Y(n_1802)
);

INVx3_ASAP7_75t_L g1803 ( 
.A(n_1750),
.Y(n_1803)
);

OAI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1755),
.A2(n_1723),
.B1(n_1711),
.B2(n_1728),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1744),
.B(n_1737),
.Y(n_1805)
);

AOI221xp5_ASAP7_75t_L g1806 ( 
.A1(n_1743),
.A2(n_1692),
.B1(n_1691),
.B2(n_1716),
.C(n_1734),
.Y(n_1806)
);

INVx1_ASAP7_75t_SL g1807 ( 
.A(n_1754),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1737),
.B(n_1689),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1743),
.A2(n_1711),
.B1(n_1728),
.B2(n_1695),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1757),
.B(n_1682),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1769),
.A2(n_1718),
.B1(n_1730),
.B2(n_1732),
.Y(n_1811)
);

OAI332xp33_ASAP7_75t_L g1812 ( 
.A1(n_1739),
.A2(n_1702),
.A3(n_1707),
.B1(n_1732),
.B2(n_1713),
.B3(n_1698),
.C1(n_1687),
.C2(n_1688),
.Y(n_1812)
);

AO21x2_ASAP7_75t_L g1813 ( 
.A1(n_1771),
.A2(n_1692),
.B(n_1714),
.Y(n_1813)
);

AOI33xp33_ASAP7_75t_L g1814 ( 
.A1(n_1746),
.A2(n_1698),
.A3(n_1688),
.B1(n_1687),
.B2(n_1707),
.B3(n_1729),
.Y(n_1814)
);

OA211x2_ASAP7_75t_L g1815 ( 
.A1(n_1751),
.A2(n_1765),
.B(n_1766),
.C(n_1758),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1759),
.Y(n_1816)
);

O2A1O1Ixp33_ASAP7_75t_SL g1817 ( 
.A1(n_1754),
.A2(n_1721),
.B(n_1697),
.C(n_1718),
.Y(n_1817)
);

OAI21xp33_ASAP7_75t_L g1818 ( 
.A1(n_1798),
.A2(n_1762),
.B(n_1758),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1773),
.Y(n_1819)
);

OA21x2_ASAP7_75t_L g1820 ( 
.A1(n_1780),
.A2(n_1806),
.B(n_1811),
.Y(n_1820)
);

NAND3xp33_ASAP7_75t_SL g1821 ( 
.A(n_1779),
.B(n_1762),
.C(n_1690),
.Y(n_1821)
);

HB1xp67_ASAP7_75t_L g1822 ( 
.A(n_1787),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1775),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1786),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1813),
.Y(n_1826)
);

AOI21x1_ASAP7_75t_L g1827 ( 
.A1(n_1809),
.A2(n_1706),
.B(n_1714),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1797),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1790),
.B(n_1772),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1814),
.B(n_1763),
.Y(n_1830)
);

BUFx6f_ASAP7_75t_L g1831 ( 
.A(n_1788),
.Y(n_1831)
);

NAND3xp33_ASAP7_75t_SL g1832 ( 
.A(n_1774),
.B(n_1795),
.C(n_1799),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1794),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1786),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1800),
.Y(n_1835)
);

HB1xp67_ASAP7_75t_L g1836 ( 
.A(n_1783),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1813),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1813),
.Y(n_1838)
);

HB1xp67_ASAP7_75t_L g1839 ( 
.A(n_1783),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1784),
.Y(n_1840)
);

NOR2xp33_ASAP7_75t_L g1841 ( 
.A(n_1812),
.B(n_1736),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1791),
.B(n_1770),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1791),
.B(n_1770),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1777),
.B(n_1762),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1784),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1816),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1782),
.Y(n_1847)
);

NOR2x1p5_ASAP7_75t_L g1848 ( 
.A(n_1810),
.B(n_1671),
.Y(n_1848)
);

AO21x2_ASAP7_75t_L g1849 ( 
.A1(n_1817),
.A2(n_1702),
.B(n_1701),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1814),
.B(n_1763),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1782),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1801),
.Y(n_1852)
);

BUFx2_ASAP7_75t_L g1853 ( 
.A(n_1790),
.Y(n_1853)
);

BUFx3_ASAP7_75t_L g1854 ( 
.A(n_1803),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1833),
.Y(n_1855)
);

AO22x1_ASAP7_75t_L g1856 ( 
.A1(n_1831),
.A2(n_1772),
.B1(n_1778),
.B2(n_1817),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1833),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1853),
.B(n_1848),
.Y(n_1858)
);

NAND2xp33_ASAP7_75t_SL g1859 ( 
.A(n_1853),
.B(n_1776),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1830),
.B(n_1736),
.Y(n_1860)
);

INVxp67_ASAP7_75t_SL g1861 ( 
.A(n_1831),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1853),
.B(n_1777),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1848),
.B(n_1747),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1831),
.B(n_1785),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1831),
.B(n_1785),
.Y(n_1865)
);

NOR2xp33_ASAP7_75t_L g1866 ( 
.A(n_1831),
.B(n_1789),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1834),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1830),
.B(n_1801),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1829),
.B(n_1747),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1833),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1831),
.Y(n_1871)
);

HB1xp67_ASAP7_75t_L g1872 ( 
.A(n_1822),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1831),
.B(n_1781),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1831),
.B(n_1844),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1846),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1834),
.Y(n_1876)
);

INVx1_ASAP7_75t_SL g1877 ( 
.A(n_1822),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1846),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1846),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1841),
.B(n_1742),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1829),
.B(n_1803),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1842),
.B(n_1805),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1842),
.B(n_1742),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1850),
.B(n_1808),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1841),
.B(n_1807),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1819),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1819),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1828),
.Y(n_1889)
);

AOI221xp5_ASAP7_75t_L g1890 ( 
.A1(n_1832),
.A2(n_1804),
.B1(n_1793),
.B2(n_1752),
.C(n_1748),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1850),
.B(n_1792),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1832),
.B(n_1764),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1823),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1842),
.B(n_1808),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1843),
.B(n_1761),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1823),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1887),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1880),
.B(n_1836),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1855),
.Y(n_1899)
);

INVx2_ASAP7_75t_L g1900 ( 
.A(n_1882),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1882),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1873),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1867),
.Y(n_1903)
);

OAI211xp5_ASAP7_75t_SL g1904 ( 
.A1(n_1886),
.A2(n_1818),
.B(n_1824),
.C(n_1825),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1887),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1862),
.B(n_1847),
.Y(n_1906)
);

INVx3_ASAP7_75t_SL g1907 ( 
.A(n_1877),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1891),
.B(n_1836),
.Y(n_1908)
);

NAND2x1p5_ASAP7_75t_L g1909 ( 
.A(n_1869),
.B(n_1871),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_SL g1910 ( 
.A1(n_1869),
.A2(n_1821),
.B(n_1834),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1855),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1877),
.B(n_1839),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1862),
.B(n_1847),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1857),
.Y(n_1914)
);

NAND2x1p5_ASAP7_75t_L g1915 ( 
.A(n_1869),
.B(n_1834),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1858),
.B(n_1851),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1892),
.B(n_1866),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1857),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1858),
.B(n_1851),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1884),
.B(n_1839),
.Y(n_1920)
);

NAND3xp33_ASAP7_75t_L g1921 ( 
.A(n_1856),
.B(n_1820),
.C(n_1818),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1872),
.B(n_1840),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1867),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1884),
.B(n_1840),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1860),
.B(n_1852),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.Y(n_1926)
);

NAND4xp25_ASAP7_75t_L g1927 ( 
.A(n_1859),
.B(n_1821),
.C(n_1815),
.D(n_1854),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1888),
.Y(n_1928)
);

INVxp67_ASAP7_75t_L g1929 ( 
.A(n_1889),
.Y(n_1929)
);

AOI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1856),
.A2(n_1802),
.B1(n_1796),
.B2(n_1820),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1888),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1883),
.B(n_1873),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1860),
.B(n_1868),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1871),
.Y(n_1934)
);

INVx1_ASAP7_75t_SL g1935 ( 
.A(n_1874),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_1907),
.B(n_1863),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1912),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1932),
.B(n_1883),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1899),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1932),
.B(n_1874),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1907),
.B(n_1894),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1900),
.Y(n_1942)
);

NOR2xp33_ASAP7_75t_L g1943 ( 
.A(n_1898),
.B(n_1863),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1900),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1899),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1920),
.B(n_1864),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1921),
.A2(n_1820),
.B1(n_1890),
.B2(n_1849),
.Y(n_1947)
);

INVx1_ASAP7_75t_SL g1948 ( 
.A(n_1935),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1902),
.B(n_1869),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1929),
.B(n_1863),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1902),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1911),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1911),
.Y(n_1953)
);

AND2x2_ASAP7_75t_L g1954 ( 
.A(n_1920),
.B(n_1864),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1916),
.B(n_1894),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1901),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1916),
.B(n_1868),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_SL g1958 ( 
.A1(n_1917),
.A2(n_1820),
.B1(n_1849),
.B2(n_1824),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1901),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1924),
.B(n_1865),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1924),
.B(n_1865),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1919),
.B(n_1895),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1922),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1939),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1939),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_SL g1966 ( 
.A1(n_1963),
.A2(n_1908),
.B1(n_1861),
.B2(n_1863),
.Y(n_1966)
);

NOR3xp33_ASAP7_75t_L g1967 ( 
.A(n_1936),
.B(n_1904),
.C(n_1927),
.Y(n_1967)
);

OAI21x1_ASAP7_75t_L g1968 ( 
.A1(n_1941),
.A2(n_1909),
.B(n_1915),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1949),
.Y(n_1969)
);

OAI21xp5_ASAP7_75t_SL g1970 ( 
.A1(n_1947),
.A2(n_1930),
.B(n_1909),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1945),
.Y(n_1971)
);

AOI211xp5_ASAP7_75t_L g1972 ( 
.A1(n_1963),
.A2(n_1910),
.B(n_1937),
.C(n_1942),
.Y(n_1972)
);

OAI221xp5_ASAP7_75t_SL g1973 ( 
.A1(n_1958),
.A2(n_1910),
.B1(n_1933),
.B2(n_1885),
.C(n_1925),
.Y(n_1973)
);

AOI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1943),
.A2(n_1820),
.B1(n_1849),
.B2(n_1919),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1942),
.B(n_1906),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1957),
.A2(n_1820),
.B1(n_1849),
.B2(n_1933),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1945),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_L g1978 ( 
.A(n_1948),
.B(n_1909),
.Y(n_1978)
);

AOI222xp33_ASAP7_75t_L g1979 ( 
.A1(n_1944),
.A2(n_1824),
.B1(n_1825),
.B2(n_1838),
.C1(n_1826),
.C2(n_1837),
.Y(n_1979)
);

NAND2xp33_ASAP7_75t_SL g1980 ( 
.A(n_1940),
.B(n_1906),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1944),
.B(n_1913),
.Y(n_1981)
);

AOI322xp5_ASAP7_75t_L g1982 ( 
.A1(n_1956),
.A2(n_1824),
.A3(n_1825),
.B1(n_1913),
.B2(n_1876),
.C1(n_1838),
.C2(n_1837),
.Y(n_1982)
);

OAI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1951),
.A2(n_1827),
.B(n_1915),
.Y(n_1983)
);

AOI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1950),
.A2(n_1849),
.B1(n_1824),
.B2(n_1825),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1938),
.B(n_1895),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1938),
.B(n_1956),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1985),
.B(n_1946),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1975),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1969),
.B(n_1959),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_SL g1990 ( 
.A(n_1972),
.B(n_1959),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1986),
.B(n_1946),
.Y(n_1991)
);

NOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1975),
.B(n_1952),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1981),
.B(n_1954),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1981),
.Y(n_1994)
);

AND2x2_ASAP7_75t_SL g1995 ( 
.A(n_1967),
.B(n_1949),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1978),
.B(n_1954),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1964),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1973),
.B(n_1980),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1966),
.B(n_1960),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1965),
.Y(n_2000)
);

AOI21xp5_ASAP7_75t_L g2001 ( 
.A1(n_1990),
.A2(n_1970),
.B(n_1983),
.Y(n_2001)
);

AND3x1_ASAP7_75t_L g2002 ( 
.A(n_1998),
.B(n_1940),
.C(n_1971),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_1990),
.A2(n_1968),
.B(n_1974),
.C(n_1977),
.Y(n_2003)
);

NOR4xp25_ASAP7_75t_L g2004 ( 
.A(n_1989),
.B(n_1976),
.C(n_1952),
.D(n_1953),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1987),
.B(n_1955),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1995),
.A2(n_1984),
.B1(n_1949),
.B2(n_1960),
.Y(n_2006)
);

OAI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1998),
.A2(n_1982),
.B(n_1949),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1992),
.A2(n_1934),
.B(n_1953),
.Y(n_2008)
);

NAND3xp33_ASAP7_75t_SL g2009 ( 
.A(n_1999),
.B(n_1915),
.C(n_1961),
.Y(n_2009)
);

OR2x2_ASAP7_75t_L g2010 ( 
.A(n_1993),
.B(n_1962),
.Y(n_2010)
);

AOI21xp5_ASAP7_75t_L g2011 ( 
.A1(n_1995),
.A2(n_1934),
.B(n_1961),
.Y(n_2011)
);

AOI221xp5_ASAP7_75t_L g2012 ( 
.A1(n_1988),
.A2(n_1825),
.B1(n_1876),
.B2(n_1923),
.C(n_1926),
.Y(n_2012)
);

INVxp67_ASAP7_75t_L g2013 ( 
.A(n_2002),
.Y(n_2013)
);

AOI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_2004),
.A2(n_1991),
.B1(n_1994),
.B2(n_1996),
.Y(n_2014)
);

INVxp67_ASAP7_75t_L g2015 ( 
.A(n_2005),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_2010),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_L g2017 ( 
.A(n_2009),
.B(n_1987),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2011),
.B(n_1997),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_2008),
.B(n_2000),
.Y(n_2019)
);

NOR2x1_ASAP7_75t_L g2020 ( 
.A(n_2007),
.B(n_1903),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2006),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_2016),
.B(n_2001),
.Y(n_2022)
);

INVxp67_ASAP7_75t_L g2023 ( 
.A(n_2017),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_2015),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2018),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_2020),
.B(n_2003),
.Y(n_2026)
);

AOI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_2019),
.A2(n_2012),
.B(n_1923),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_2013),
.B(n_1897),
.Y(n_2028)
);

INVxp67_ASAP7_75t_SL g2029 ( 
.A(n_2014),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2025),
.B(n_2021),
.Y(n_2030)
);

HB1xp67_ASAP7_75t_L g2031 ( 
.A(n_2026),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2022),
.Y(n_2032)
);

INVx2_ASAP7_75t_SL g2033 ( 
.A(n_2024),
.Y(n_2033)
);

NOR2x1_ASAP7_75t_L g2034 ( 
.A(n_2028),
.B(n_1903),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_2023),
.B(n_1926),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2030),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2032),
.B(n_2029),
.Y(n_2037)
);

A2O1A1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_2031),
.A2(n_2027),
.B(n_1876),
.C(n_1931),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2035),
.A2(n_1918),
.B(n_1914),
.C(n_1928),
.Y(n_2039)
);

NOR2xp67_ASAP7_75t_L g2040 ( 
.A(n_2036),
.B(n_2033),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_2037),
.B(n_2034),
.Y(n_2041)
);

NOR3xp33_ASAP7_75t_L g2042 ( 
.A(n_2041),
.B(n_2031),
.C(n_2038),
.Y(n_2042)
);

AOI221xp5_ASAP7_75t_L g2043 ( 
.A1(n_2040),
.A2(n_2039),
.B1(n_1914),
.B2(n_1918),
.C(n_1905),
.Y(n_2043)
);

AOI21xp5_ASAP7_75t_L g2044 ( 
.A1(n_2042),
.A2(n_1925),
.B(n_1979),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_2043),
.B(n_1870),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2045),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2044),
.B(n_1885),
.Y(n_2047)
);

OAI22xp5_ASAP7_75t_SL g2048 ( 
.A1(n_2046),
.A2(n_1881),
.B1(n_1870),
.B2(n_1875),
.Y(n_2048)
);

CKINVDCx20_ASAP7_75t_R g2049 ( 
.A(n_2047),
.Y(n_2049)
);

O2A1O1Ixp33_ASAP7_75t_L g2050 ( 
.A1(n_2049),
.A2(n_1879),
.B(n_1878),
.C(n_1875),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_R g2051 ( 
.A(n_2050),
.B(n_2048),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2051),
.B(n_1878),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2052),
.A2(n_1879),
.B1(n_1896),
.B2(n_1893),
.Y(n_2053)
);

AOI22xp5_ASAP7_75t_L g2054 ( 
.A1(n_2053),
.A2(n_1896),
.B1(n_1893),
.B2(n_1845),
.Y(n_2054)
);

AOI211xp5_ASAP7_75t_L g2055 ( 
.A1(n_2054),
.A2(n_1828),
.B(n_1835),
.C(n_1881),
.Y(n_2055)
);


endmodule