module fake_jpeg_28248_n_162 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx6f_ASAP7_75t_SL g52 ( 
.A(n_24),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_12),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_0),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_58),
.B1(n_52),
.B2(n_62),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_71),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_75),
.B(n_55),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_59),
.B1(n_62),
.B2(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_77),
.Y(n_98)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_81),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx6f_ASAP7_75t_SL g86 ( 
.A(n_83),
.Y(n_86)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_76),
.B(n_53),
.Y(n_89)
);

NOR2x1_ASAP7_75t_R g113 ( 
.A(n_89),
.B(n_64),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_73),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_92),
.A2(n_59),
.B1(n_85),
.B2(n_79),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_95),
.Y(n_104)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_82),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_100),
.B(n_56),
.Y(n_105)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_105),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_64),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_43),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_60),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_111),
.B(n_45),
.Y(n_124)
);

NOR3xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_96),
.C(n_94),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_116),
.B(n_118),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_113),
.B(n_96),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_104),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_56),
.B(n_51),
.C(n_87),
.D(n_63),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_42),
.C(n_57),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_54),
.C(n_49),
.Y(n_127)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_121),
.Y(n_132)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_101),
.B1(n_99),
.B2(n_98),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_106),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_123),
.A2(n_112),
.B1(n_86),
.B2(n_55),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_114),
.A2(n_112),
.B1(n_99),
.B2(n_98),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_133),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_127),
.C(n_128),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_63),
.C(n_108),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_129),
.A2(n_130),
.B1(n_136),
.B2(n_11),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_47),
.B1(n_44),
.B2(n_54),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_115),
.A2(n_44),
.B1(n_47),
.B2(n_4),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_131),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_1),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_139),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_10),
.Y(n_138)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_10),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_11),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.C(n_142),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_28),
.B1(n_39),
.B2(n_13),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_129),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_130),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_149),
.A2(n_144),
.B1(n_139),
.B2(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_146),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_145),
.B(n_148),
.C(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_149),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_31),
.B(n_14),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_156),
.Y(n_157)
);

OAI21x1_ASAP7_75t_SL g158 ( 
.A1(n_157),
.A2(n_33),
.B(n_15),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_34),
.C(n_16),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_36),
.C(n_18),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_37),
.B(n_20),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_21),
.Y(n_162)
);


endmodule