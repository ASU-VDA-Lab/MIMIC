module fake_jpeg_5809_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_17),
.Y(n_69)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_17),
.Y(n_49)
);

AO22x1_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_17),
.B1(n_33),
.B2(n_19),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_29),
.B1(n_18),
.B2(n_21),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_56),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_18),
.B1(n_30),
.B2(n_21),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_66),
.B1(n_67),
.B2(n_33),
.Y(n_89)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_36),
.B(n_32),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_69),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_0),
.Y(n_90)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_41),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_32),
.B1(n_19),
.B2(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_25),
.B1(n_17),
.B2(n_22),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_22),
.B(n_19),
.C(n_33),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_65),
.B(n_60),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_52),
.B(n_57),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_73),
.B(n_47),
.C(n_7),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_34),
.B(n_25),
.C(n_10),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_67),
.B(n_49),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_76),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_79),
.Y(n_102)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_80),
.Y(n_113)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_34),
.C(n_25),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_51),
.C(n_62),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_25),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_77),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_55),
.B1(n_66),
.B2(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_48),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_105),
.B(n_111),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_94),
.A2(n_112),
.B1(n_74),
.B2(n_75),
.Y(n_126)
);

OAI22x1_ASAP7_75t_L g134 ( 
.A1(n_95),
.A2(n_92),
.B1(n_94),
.B2(n_103),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_101),
.B(n_107),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_69),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_103),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_56),
.B(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_45),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_130),
.B1(n_93),
.B2(n_113),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_80),
.B(n_88),
.C(n_74),
.D(n_75),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_121),
.B(n_109),
.Y(n_154)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_123),
.Y(n_160)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_124),
.B(n_127),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_102),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_45),
.B1(n_53),
.B2(n_85),
.Y(n_161)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_91),
.B1(n_60),
.B2(n_68),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_76),
.B(n_78),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_98),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_136),
.B(n_108),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_98),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_113),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_141),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_145),
.B(n_118),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_115),
.C(n_116),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_146),
.B(n_58),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_95),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_154),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_150),
.B(n_158),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_107),
.B1(n_93),
.B2(n_112),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_151),
.A2(n_121),
.B1(n_63),
.B2(n_58),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_164),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_60),
.B1(n_106),
.B2(n_79),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_156),
.A2(n_140),
.B1(n_86),
.B2(n_122),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_128),
.A2(n_134),
.B(n_119),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_157),
.A2(n_168),
.B(n_166),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_99),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_163),
.B1(n_118),
.B2(n_53),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_126),
.A2(n_84),
.B1(n_86),
.B2(n_85),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_84),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_76),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_131),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_142),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_176),
.B(n_144),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_188),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_133),
.B1(n_136),
.B2(n_120),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_175),
.A2(n_190),
.B1(n_159),
.B2(n_1),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_168),
.A2(n_160),
.B(n_128),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_177),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_117),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_180),
.B(n_186),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_161),
.B1(n_167),
.B2(n_146),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_58),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_189),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_141),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_1),
.C(n_2),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_158),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_53),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_76),
.B1(n_78),
.B2(n_63),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_148),
.B(n_8),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_8),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_176),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_172),
.B(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_190),
.B1(n_150),
.B2(n_151),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_213),
.B1(n_194),
.B2(n_2),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_208),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_211),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_173),
.A2(n_153),
.B1(n_148),
.B2(n_143),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_206),
.A2(n_207),
.B1(n_214),
.B2(n_174),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_153),
.B1(n_169),
.B2(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_165),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_149),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_210),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_149),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_184),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_187),
.C(n_175),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_180),
.Y(n_219)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_210),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_182),
.C(n_170),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_223),
.C(n_224),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_192),
.Y(n_224)
);

XOR2x1_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_192),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_205),
.B1(n_207),
.B2(n_196),
.Y(n_235)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_193),
.B(n_179),
.C(n_171),
.D(n_189),
.Y(n_227)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_208),
.C(n_198),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_229),
.B(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_233),
.B1(n_216),
.B2(n_214),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_9),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_231),
.B(n_215),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_3),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_234),
.B(n_199),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_244),
.C(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_243),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_227),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_198),
.B(n_203),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_248),
.B(n_228),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_225),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_222),
.B(n_216),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_250),
.C(n_256),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_218),
.C(n_232),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_239),
.A2(n_200),
.B1(n_211),
.B2(n_223),
.Y(n_251)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_221),
.C(n_231),
.Y(n_256)
);

NOR4xp25_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_200),
.C(n_224),
.D(n_211),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_260),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_242),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_247),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_259),
.A2(n_245),
.B(n_6),
.Y(n_268)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_241),
.B(n_204),
.CI(n_209),
.CON(n_260),
.SN(n_260)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_262),
.B(n_268),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_242),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_263),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_5),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_269),
.A2(n_254),
.B(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_266),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_7),
.B(n_9),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_272),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_256),
.C(n_260),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.C(n_6),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_5),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_279),
.A2(n_280),
.B(n_281),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_10),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_277),
.A2(n_273),
.B(n_276),
.Y(n_282)
);

AOI321xp33_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_274),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C(n_16),
.Y(n_286)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_284),
.B(n_12),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_11),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_290)
);


endmodule