module fake_jpeg_15011_n_26 (n_3, n_2, n_1, n_0, n_4, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx11_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

INVx8_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx13_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_11),
.Y(n_14)
);

CKINVDCx9p33_ASAP7_75t_R g11 ( 
.A(n_5),
.Y(n_11)
);

AOI22xp33_ASAP7_75t_SL g12 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g15 ( 
.A(n_12),
.B(n_0),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_8),
.B1(n_5),
.B2(n_6),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_13),
.B(n_9),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_18),
.Y(n_20)
);

FAx1_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_14),
.CI(n_6),
.CON(n_21),
.SN(n_21)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_7),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_6),
.Y(n_19)
);

MAJx2_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_10),
.C(n_6),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_10),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_7),
.B(n_2),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_1),
.B1(n_4),
.B2(n_12),
.Y(n_26)
);


endmodule