module fake_netlist_1_2250_n_29 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
BUFx6f_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
AND2x6_ASAP7_75t_L g13 ( .A(n_3), .B(n_9), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_3), .B(n_0), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_6), .Y(n_15) );
BUFx6f_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_12), .B(n_15), .Y(n_18) );
AO21x2_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_14), .B(n_13), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_19), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
AOI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_20), .B1(n_19), .B2(n_16), .C(n_12), .Y(n_23) );
NOR2x1_ASAP7_75t_L g24 ( .A(n_23), .B(n_16), .Y(n_24) );
NAND4xp75_ASAP7_75t_L g25 ( .A(n_24), .B(n_13), .C(n_2), .D(n_1), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_1), .Y(n_26) );
OAI22xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_12), .B1(n_13), .B2(n_2), .Y(n_27) );
O2A1O1Ixp33_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_25), .B(n_5), .C(n_7), .Y(n_28) );
OAI21xp33_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_4), .B(n_8), .Y(n_29) );
endmodule