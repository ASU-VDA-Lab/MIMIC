module fake_jpeg_19393_n_176 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_176);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_42),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_12),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_17),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_27),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_68),
.Y(n_84)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_68),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_93),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_66),
.B(n_77),
.C(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_99),
.Y(n_103)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_56),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_95),
.A2(n_97),
.B1(n_58),
.B2(n_62),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_100),
.Y(n_122)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_101),
.A2(n_109),
.B1(n_111),
.B2(n_98),
.Y(n_114)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_63),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_88),
.A2(n_53),
.B1(n_79),
.B2(n_60),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_65),
.B1(n_59),
.B2(n_69),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g112 ( 
.A(n_92),
.B(n_51),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_97),
.C(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_55),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_61),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_128),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_123),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_78),
.B1(n_76),
.B2(n_75),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_72),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_57),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_64),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_100),
.C(n_71),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_45),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_126),
.A2(n_114),
.B1(n_121),
.B2(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_140),
.B1(n_142),
.B2(n_4),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_121),
.A2(n_127),
.B1(n_122),
.B2(n_119),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_69),
.B1(n_2),
.B2(n_3),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_141),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_120),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_136),
.A2(n_26),
.B1(n_44),
.B2(n_43),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_144),
.A2(n_152),
.B1(n_7),
.B2(n_8),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_146),
.B(n_149),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_139),
.A2(n_21),
.B(n_39),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_1),
.Y(n_149)
);

FAx1_ASAP7_75t_SL g150 ( 
.A(n_137),
.B(n_19),
.CI(n_36),
.CON(n_150),
.SN(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_136),
.B(n_31),
.C(n_22),
.D(n_41),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_151),
.A2(n_153),
.B1(n_129),
.B2(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_147),
.B1(n_143),
.B2(n_10),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_161),
.C(n_146),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_158),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_163),
.B(n_164),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_154),
.C(n_159),
.Y(n_164)
);

AOI21x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_145),
.B(n_155),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_150),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_144),
.B1(n_160),
.B2(n_32),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_30),
.C(n_34),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_13),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_33),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_35),
.B(n_9),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_11),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_8),
.Y(n_176)
);


endmodule