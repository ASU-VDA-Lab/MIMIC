module fake_jpeg_21795_n_258 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_258);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_258;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_3),
.B(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_34),
.A2(n_35),
.B(n_26),
.C(n_23),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_31),
.B1(n_25),
.B2(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_42),
.B(n_30),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_35),
.C(n_29),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_46),
.A2(n_51),
.B1(n_40),
.B2(n_20),
.Y(n_64)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NAND2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_49),
.A2(n_42),
.B(n_27),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_25),
.B1(n_31),
.B2(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_40),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_29),
.B1(n_27),
.B2(n_17),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_36),
.B1(n_17),
.B2(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_59),
.B(n_79),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_23),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_69),
.B(n_71),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_64),
.A2(n_66),
.B1(n_68),
.B2(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_42),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_18),
.B1(n_28),
.B2(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_40),
.B1(n_38),
.B2(n_37),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_50),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_74),
.B(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_55),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_52),
.B(n_1),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_15),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_81),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_23),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_40),
.B1(n_32),
.B2(n_22),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_54),
.B1(n_50),
.B2(n_37),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_1),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_50),
.Y(n_104)
);

XOR2x2_ASAP7_75t_L g86 ( 
.A(n_60),
.B(n_71),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_56),
.B(n_58),
.C(n_67),
.D(n_75),
.Y(n_114)
);

BUFx2_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_89),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_90),
.A2(n_84),
.B1(n_62),
.B2(n_83),
.Y(n_126)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_105),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_108),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_93),
.B(n_76),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_63),
.B(n_62),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_59),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_54),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_71),
.B(n_37),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_61),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_37),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_111),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_114),
.A2(n_115),
.B(n_122),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_123),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_57),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_92),
.Y(n_145)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_127),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_79),
.B1(n_83),
.B2(n_87),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_128),
.B(n_134),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_72),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

OR2x4_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_61),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_131),
.B(n_93),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_64),
.B(n_74),
.C(n_68),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_132),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_85),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_135),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_61),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_33),
.B(n_73),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_100),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_106),
.Y(n_141)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

AO22x1_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_108),
.B1(n_100),
.B2(n_109),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_142),
.A2(n_150),
.B1(n_151),
.B2(n_131),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_123),
.A2(n_87),
.B1(n_102),
.B2(n_101),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_143),
.A2(n_147),
.B(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_149),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_111),
.A2(n_87),
.B1(n_102),
.B2(n_101),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_112),
.B1(n_106),
.B2(n_108),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_108),
.B1(n_95),
.B2(n_110),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_154),
.A2(n_161),
.B(n_163),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_122),
.A2(n_83),
.B1(n_94),
.B2(n_109),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_125),
.B1(n_127),
.B2(n_136),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_109),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_114),
.C(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_166),
.C(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_165),
.A2(n_167),
.B1(n_146),
.B2(n_162),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_136),
.C(n_115),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_115),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_153),
.B(n_117),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_175),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_176),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_19),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_116),
.C(n_118),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_128),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_118),
.C(n_73),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_180),
.Y(n_190)
);

INVxp33_ASAP7_75t_SL g179 ( 
.A(n_138),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g203 ( 
.A(n_179),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_33),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_148),
.C(n_150),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_186),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_32),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_152),
.Y(n_185)
);

NOR3xp33_ASAP7_75t_SL g187 ( 
.A(n_185),
.B(n_158),
.C(n_149),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_148),
.B(n_33),
.C(n_32),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_189),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_184),
.A2(n_154),
.B1(n_161),
.B2(n_139),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_200),
.B1(n_169),
.B2(n_172),
.Y(n_210)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_151),
.A3(n_163),
.B1(n_141),
.B2(n_159),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_196),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_2),
.B(n_7),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_22),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_22),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_171),
.B(n_186),
.Y(n_205)
);

AO22x2_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_19),
.B1(n_4),
.B2(n_5),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_206),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_197),
.A2(n_170),
.B1(n_181),
.B2(n_166),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_216),
.B1(n_200),
.B2(n_188),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_215),
.Y(n_227)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_211),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

NOR3xp33_ASAP7_75t_SL g213 ( 
.A(n_187),
.B(n_164),
.C(n_173),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_177),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g221 ( 
.A(n_214),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_201),
.C(n_200),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_222),
.B(n_205),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_190),
.C(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_191),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_216),
.A2(n_218),
.B1(n_207),
.B2(n_217),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_217),
.B1(n_208),
.B2(n_192),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_212),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_232),
.A2(n_234),
.B(n_223),
.Y(n_239)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_235),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_225),
.A2(n_215),
.B(n_213),
.Y(n_234)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_2),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_237),
.B(n_7),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_7),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_227),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_239),
.A2(n_230),
.B(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_9),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_248),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_249),
.B(n_250),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_235),
.Y(n_250)
);

AOI322xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_245),
.A3(n_243),
.B1(n_226),
.B2(n_227),
.C1(n_13),
.C2(n_9),
.Y(n_252)
);

AOI322xp5_ASAP7_75t_L g255 ( 
.A1(n_252),
.A2(n_243),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_14),
.C2(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_251),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_254),
.A2(n_255),
.B(n_10),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_10),
.B(n_11),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_12),
.Y(n_258)
);


endmodule