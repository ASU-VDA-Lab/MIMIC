module real_aes_15573_n_4 (n_0, n_3, n_2, n_1, n_4);
input n_0;
input n_3;
input n_2;
input n_1;
output n_4;
wire n_5;
wire n_7;
wire n_8;
wire n_6;
wire n_9;
wire n_10;
CKINVDCx5p33_ASAP7_75t_R g7 ( .A(n_0), .Y(n_7) );
NOR2xp33_ASAP7_75t_R g9 ( .A(n_0), .B(n_10), .Y(n_9) );
OAI22xp33_ASAP7_75t_SL g4 ( .A1(n_1), .A2(n_2), .B1(n_5), .B2(n_8), .Y(n_4) );
NOR2xp33_ASAP7_75t_R g6 ( .A(n_3), .B(n_7), .Y(n_6) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_3), .Y(n_10) );
INVxp33_ASAP7_75t_SL g5 ( .A(n_6), .Y(n_5) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_9), .Y(n_8) );
endmodule