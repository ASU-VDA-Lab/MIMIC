module real_aes_7028_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_504;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_527;
wire n_505;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_0), .B(n_89), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g461 ( .A(n_0), .Y(n_461) );
INVx1_ASAP7_75t_L g496 ( .A(n_1), .Y(n_496) );
INVx1_ASAP7_75t_L g202 ( .A(n_2), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_3), .A2(n_38), .B1(n_163), .B2(n_526), .Y(n_541) );
AOI21xp33_ASAP7_75t_L g170 ( .A1(n_4), .A2(n_144), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_5), .B(n_137), .Y(n_509) );
AND2x6_ASAP7_75t_L g149 ( .A(n_6), .B(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_7), .A2(n_252), .B(n_253), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g106 ( .A(n_8), .B(n_39), .Y(n_106) );
INVx1_ASAP7_75t_L g177 ( .A(n_9), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_10), .B(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g142 ( .A(n_11), .Y(n_142) );
INVx1_ASAP7_75t_L g490 ( .A(n_12), .Y(n_490) );
INVx1_ASAP7_75t_L g258 ( .A(n_13), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_14), .B(n_185), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_15), .B(n_138), .Y(n_567) );
AO32x2_ASAP7_75t_L g539 ( .A1(n_16), .A2(n_137), .A3(n_182), .B1(n_518), .B2(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g104 ( .A1(n_17), .A2(n_105), .B1(n_112), .B2(n_775), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_18), .A2(n_63), .B1(n_126), .B2(n_127), .Y(n_125) );
INVx1_ASAP7_75t_L g127 ( .A(n_18), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_19), .B(n_163), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_20), .B(n_158), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_21), .B(n_138), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_22), .A2(n_51), .B1(n_163), .B2(n_526), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_23), .B(n_144), .Y(n_214) );
AOI22xp33_ASAP7_75t_SL g527 ( .A1(n_24), .A2(n_80), .B1(n_163), .B2(n_185), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_25), .B(n_163), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_26), .B(n_166), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_27), .A2(n_256), .B(n_257), .C(n_259), .Y(n_255) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_28), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_29), .B(n_179), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_30), .B(n_175), .Y(n_204) );
INVx1_ASAP7_75t_L g191 ( .A(n_31), .Y(n_191) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_32), .A2(n_33), .B1(n_120), .B2(n_121), .Y(n_119) );
INVx1_ASAP7_75t_L g121 ( .A(n_32), .Y(n_121) );
INVxp67_ASAP7_75t_L g120 ( .A(n_33), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_33), .B(n_179), .Y(n_556) );
INVx2_ASAP7_75t_L g147 ( .A(n_34), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g513 ( .A(n_35), .B(n_163), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_36), .B(n_179), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_37), .A2(n_149), .B(n_153), .C(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g189 ( .A(n_40), .Y(n_189) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_41), .A2(n_469), .B1(n_472), .B2(n_473), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_41), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_42), .B(n_175), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_43), .B(n_163), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_44), .A2(n_90), .B1(n_221), .B2(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_45), .B(n_163), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_46), .B(n_163), .Y(n_491) );
CKINVDCx16_ASAP7_75t_R g192 ( .A(n_47), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_48), .A2(n_70), .B1(n_470), .B2(n_471), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_48), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_49), .B(n_495), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_50), .B(n_144), .Y(n_246) );
AOI22xp33_ASAP7_75t_SL g565 ( .A1(n_52), .A2(n_61), .B1(n_163), .B2(n_185), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_53), .A2(n_153), .B1(n_185), .B2(n_187), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_54), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_55), .B(n_163), .Y(n_517) );
CKINVDCx16_ASAP7_75t_R g199 ( .A(n_56), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_57), .B(n_163), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g173 ( .A1(n_58), .A2(n_162), .B(n_174), .C(n_176), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_59), .Y(n_234) );
INVx1_ASAP7_75t_L g172 ( .A(n_60), .Y(n_172) );
INVx1_ASAP7_75t_L g150 ( .A(n_62), .Y(n_150) );
INVx1_ASAP7_75t_L g126 ( .A(n_63), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_64), .B(n_163), .Y(n_497) );
INVx1_ASAP7_75t_L g141 ( .A(n_65), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_66), .Y(n_116) );
AO32x2_ASAP7_75t_L g523 ( .A1(n_67), .A2(n_137), .A3(n_238), .B1(n_518), .B2(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g516 ( .A(n_68), .Y(n_516) );
INVx1_ASAP7_75t_L g551 ( .A(n_69), .Y(n_551) );
INVx1_ASAP7_75t_L g470 ( .A(n_70), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_SL g157 ( .A1(n_71), .A2(n_158), .B(n_159), .C(n_162), .Y(n_157) );
INVxp67_ASAP7_75t_L g160 ( .A(n_72), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_73), .B(n_185), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_74), .A2(n_467), .B1(n_468), .B2(n_474), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_74), .Y(n_467) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g462 ( .A(n_76), .B(n_457), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_77), .A2(n_459), .B1(n_465), .B2(n_770), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_78), .Y(n_195) );
INVx1_ASAP7_75t_L g227 ( .A(n_79), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_81), .A2(n_149), .B(n_153), .C(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_82), .B(n_526), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_83), .B(n_185), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_84), .B(n_203), .Y(n_217) );
INVx2_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_86), .B(n_158), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_87), .B(n_185), .Y(n_505) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_88), .A2(n_149), .B(n_153), .C(n_201), .Y(n_200) );
OR2x2_ASAP7_75t_L g458 ( .A(n_89), .B(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g476 ( .A(n_89), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_91), .A2(n_103), .B1(n_185), .B2(n_186), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_92), .B(n_179), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_93), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_94), .A2(n_149), .B(n_153), .C(n_241), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g248 ( .A(n_95), .Y(n_248) );
INVx1_ASAP7_75t_L g156 ( .A(n_96), .Y(n_156) );
CKINVDCx16_ASAP7_75t_R g254 ( .A(n_97), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_98), .B(n_203), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_99), .B(n_185), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_100), .B(n_137), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_101), .B(n_111), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_102), .A2(n_144), .B(n_151), .Y(n_143) );
INVx1_ASAP7_75t_L g775 ( .A(n_105), .Y(n_775) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
AND2x2_ASAP7_75t_L g460 ( .A(n_106), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_463), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g774 ( .A(n_116), .Y(n_774) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_455), .B(n_462), .Y(n_117) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_122), .B1(n_123), .B2(n_454), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_119), .Y(n_454) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_128), .B2(n_453), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g453 ( .A(n_128), .Y(n_453) );
AOI22xp5_ASAP7_75t_SL g475 ( .A1(n_128), .A2(n_476), .B1(n_477), .B2(n_769), .Y(n_475) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND4x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_371), .C(n_418), .D(n_438), .Y(n_129) );
NOR3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_301), .C(n_326), .Y(n_130) );
OAI211xp5_ASAP7_75t_SL g131 ( .A1(n_132), .A2(n_209), .B(n_261), .C(n_291), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_180), .Y(n_133) );
INVx3_ASAP7_75t_SL g343 ( .A(n_134), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_134), .B(n_274), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_134), .B(n_196), .Y(n_424) );
AND2x2_ASAP7_75t_L g447 ( .A(n_134), .B(n_313), .Y(n_447) );
AND2x4_ASAP7_75t_L g134 ( .A(n_135), .B(n_168), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g265 ( .A(n_136), .B(n_169), .Y(n_265) );
INVx3_ASAP7_75t_L g278 ( .A(n_136), .Y(n_278) );
AND2x2_ASAP7_75t_L g283 ( .A(n_136), .B(n_168), .Y(n_283) );
OR2x2_ASAP7_75t_L g334 ( .A(n_136), .B(n_275), .Y(n_334) );
BUFx2_ASAP7_75t_L g354 ( .A(n_136), .Y(n_354) );
AND2x2_ASAP7_75t_L g364 ( .A(n_136), .B(n_275), .Y(n_364) );
AND2x2_ASAP7_75t_L g370 ( .A(n_136), .B(n_181), .Y(n_370) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_143), .B(n_165), .Y(n_136) );
INVx4_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
OA21x2_ASAP7_75t_L g501 ( .A1(n_137), .A2(n_502), .B(n_509), .Y(n_501) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g182 ( .A(n_138), .Y(n_182) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_139), .B(n_140), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx2_ASAP7_75t_L g252 ( .A(n_144), .Y(n_252) );
AND2x4_ASAP7_75t_L g144 ( .A(n_145), .B(n_149), .Y(n_144) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_145), .B(n_149), .Y(n_193) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
INVx1_ASAP7_75t_L g495 ( .A(n_146), .Y(n_495) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx2_ASAP7_75t_L g154 ( .A(n_147), .Y(n_154) );
INVx1_ASAP7_75t_L g186 ( .A(n_147), .Y(n_186) );
INVx1_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
INVx1_ASAP7_75t_L g158 ( .A(n_148), .Y(n_158) );
INVx3_ASAP7_75t_L g161 ( .A(n_148), .Y(n_161) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_148), .Y(n_175) );
BUFx6f_ASAP7_75t_L g188 ( .A(n_148), .Y(n_188) );
INVx4_ASAP7_75t_SL g164 ( .A(n_149), .Y(n_164) );
OAI21xp5_ASAP7_75t_L g488 ( .A1(n_149), .A2(n_489), .B(n_493), .Y(n_488) );
OAI21xp5_ASAP7_75t_L g502 ( .A1(n_149), .A2(n_503), .B(n_506), .Y(n_502) );
BUFx3_ASAP7_75t_L g518 ( .A(n_149), .Y(n_518) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_149), .A2(n_531), .B(n_535), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_149), .A2(n_550), .B(n_553), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_156), .B(n_157), .C(n_164), .Y(n_151) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_152), .A2(n_164), .B(n_172), .C(n_173), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g253 ( .A1(n_152), .A2(n_164), .B(n_254), .C(n_255), .Y(n_253) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_154), .Y(n_163) );
BUFx3_ASAP7_75t_L g221 ( .A(n_154), .Y(n_221) );
INVx1_ASAP7_75t_L g526 ( .A(n_154), .Y(n_526) );
INVx1_ASAP7_75t_L g534 ( .A(n_158), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_161), .B(n_177), .Y(n_176) );
INVx5_ASAP7_75t_L g203 ( .A(n_161), .Y(n_203) );
OAI22xp5_ASAP7_75t_SL g524 ( .A1(n_161), .A2(n_175), .B1(n_525), .B2(n_527), .Y(n_524) );
O2A1O1Ixp5_ASAP7_75t_SL g550 ( .A1(n_162), .A2(n_203), .B(n_551), .C(n_552), .Y(n_550) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_163), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_164), .A2(n_184), .B1(n_192), .B2(n_193), .Y(n_183) );
OA21x2_ASAP7_75t_L g169 ( .A1(n_166), .A2(n_170), .B(n_178), .Y(n_169) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_SL g223 ( .A(n_167), .B(n_224), .Y(n_223) );
AO21x1_ASAP7_75t_L g562 ( .A1(n_167), .A2(n_563), .B(n_566), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_167), .B(n_518), .C(n_563), .Y(n_581) );
INVx1_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_169), .B(n_275), .Y(n_289) );
INVx2_ASAP7_75t_L g299 ( .A(n_169), .Y(n_299) );
AND2x2_ASAP7_75t_L g312 ( .A(n_169), .B(n_278), .Y(n_312) );
OR2x2_ASAP7_75t_L g323 ( .A(n_169), .B(n_275), .Y(n_323) );
AND2x2_ASAP7_75t_SL g369 ( .A(n_169), .B(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g381 ( .A(n_169), .Y(n_381) );
AND2x2_ASAP7_75t_L g427 ( .A(n_169), .B(n_181), .Y(n_427) );
O2A1O1Ixp5_ASAP7_75t_L g515 ( .A1(n_174), .A2(n_494), .B(n_516), .C(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_174), .A2(n_536), .B(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g244 ( .A(n_175), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_175), .A2(n_498), .B1(n_541), .B2(n_542), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_175), .A2(n_498), .B1(n_564), .B2(n_565), .Y(n_563) );
INVx1_ASAP7_75t_L g208 ( .A(n_179), .Y(n_208) );
INVx2_ASAP7_75t_L g238 ( .A(n_179), .Y(n_238) );
OA21x2_ASAP7_75t_L g250 ( .A1(n_179), .A2(n_251), .B(n_260), .Y(n_250) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_179), .A2(n_530), .B(n_538), .Y(n_529) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_179), .A2(n_549), .B(n_556), .Y(n_548) );
INVx3_ASAP7_75t_SL g300 ( .A(n_180), .Y(n_300) );
OR2x2_ASAP7_75t_L g353 ( .A(n_180), .B(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_196), .Y(n_180) );
INVx3_ASAP7_75t_L g275 ( .A(n_181), .Y(n_275) );
AND2x2_ASAP7_75t_L g342 ( .A(n_181), .B(n_197), .Y(n_342) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_181), .Y(n_410) );
AOI33xp33_ASAP7_75t_L g414 ( .A1(n_181), .A2(n_343), .A3(n_350), .B1(n_359), .B2(n_415), .B3(n_416), .Y(n_414) );
AO21x2_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_194), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_182), .B(n_195), .Y(n_194) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_182), .A2(n_198), .B(n_206), .Y(n_197) );
INVx2_ASAP7_75t_L g222 ( .A(n_182), .Y(n_222) );
INVx2_ASAP7_75t_L g205 ( .A(n_185), .Y(n_205) );
INVx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OAI22xp5_ASAP7_75t_SL g187 ( .A1(n_188), .A2(n_189), .B1(n_190), .B2(n_191), .Y(n_187) );
INVx2_ASAP7_75t_L g190 ( .A(n_188), .Y(n_190) );
INVx4_ASAP7_75t_L g256 ( .A(n_188), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g198 ( .A1(n_193), .A2(n_199), .B(n_200), .Y(n_198) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_193), .A2(n_227), .B(n_228), .Y(n_226) );
INVx1_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_196), .B(n_278), .Y(n_277) );
NOR3xp33_ASAP7_75t_L g337 ( .A(n_196), .B(n_338), .C(n_340), .Y(n_337) );
AND2x2_ASAP7_75t_L g363 ( .A(n_196), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_196), .B(n_370), .Y(n_373) );
AND2x2_ASAP7_75t_L g426 ( .A(n_196), .B(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g282 ( .A(n_197), .Y(n_282) );
OR2x2_ASAP7_75t_L g376 ( .A(n_197), .B(n_275), .Y(n_376) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_203), .B(n_204), .C(n_205), .Y(n_201) );
INVx2_ASAP7_75t_L g498 ( .A(n_203), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_203), .A2(n_504), .B(n_505), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_203), .A2(n_513), .B(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_205), .A2(n_490), .B(n_491), .C(n_492), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_208), .B(n_234), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_208), .B(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_235), .Y(n_209) );
AOI32xp33_ASAP7_75t_L g327 ( .A1(n_210), .A2(n_328), .A3(n_330), .B1(n_332), .B2(n_335), .Y(n_327) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_210), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g430 ( .A(n_210), .Y(n_430) );
INVx4_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g362 ( .A(n_211), .B(n_346), .Y(n_362) );
AND2x2_ASAP7_75t_L g382 ( .A(n_211), .B(n_308), .Y(n_382) );
AND2x2_ASAP7_75t_L g450 ( .A(n_211), .B(n_368), .Y(n_450) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_225), .Y(n_211) );
INVx3_ASAP7_75t_L g271 ( .A(n_212), .Y(n_271) );
AND2x2_ASAP7_75t_L g285 ( .A(n_212), .B(n_269), .Y(n_285) );
OR2x2_ASAP7_75t_L g290 ( .A(n_212), .B(n_268), .Y(n_290) );
INVx1_ASAP7_75t_L g297 ( .A(n_212), .Y(n_297) );
AND2x2_ASAP7_75t_L g305 ( .A(n_212), .B(n_279), .Y(n_305) );
AND2x2_ASAP7_75t_L g307 ( .A(n_212), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_212), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g360 ( .A(n_212), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_212), .B(n_445), .Y(n_444) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_223), .Y(n_212) );
AOI21xp5_ASAP7_75t_SL g213 ( .A1(n_214), .A2(n_215), .B(n_222), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_219), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_219), .A2(n_230), .B(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g259 ( .A(n_221), .Y(n_259) );
INVx1_ASAP7_75t_L g232 ( .A(n_222), .Y(n_232) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_222), .A2(n_488), .B(n_499), .Y(n_487) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_222), .A2(n_511), .B(n_519), .Y(n_510) );
INVx2_ASAP7_75t_L g269 ( .A(n_225), .Y(n_269) );
AND2x2_ASAP7_75t_L g315 ( .A(n_225), .B(n_236), .Y(n_315) );
AND2x2_ASAP7_75t_L g325 ( .A(n_225), .B(n_250), .Y(n_325) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_232), .B(n_233), .Y(n_225) );
INVx2_ASAP7_75t_L g445 ( .A(n_235), .Y(n_445) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_249), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_236), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g286 ( .A(n_236), .Y(n_286) );
AND2x2_ASAP7_75t_L g330 ( .A(n_236), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g346 ( .A(n_236), .B(n_309), .Y(n_346) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g294 ( .A(n_237), .Y(n_294) );
AND2x2_ASAP7_75t_L g308 ( .A(n_237), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g359 ( .A(n_237), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_237), .B(n_269), .Y(n_391) );
AO21x2_ASAP7_75t_L g237 ( .A1(n_238), .A2(n_239), .B(n_247), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_240), .B(n_246), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_245), .Y(n_241) );
AND2x2_ASAP7_75t_L g270 ( .A(n_249), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g331 ( .A(n_249), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_249), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g368 ( .A(n_249), .Y(n_368) );
INVx1_ASAP7_75t_L g401 ( .A(n_249), .Y(n_401) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g279 ( .A(n_250), .B(n_269), .Y(n_279) );
INVx1_ASAP7_75t_L g309 ( .A(n_250), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_256), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g492 ( .A(n_256), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_256), .A2(n_554), .B(n_555), .Y(n_553) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_266), .B1(n_272), .B2(n_279), .C(n_280), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_263), .B(n_283), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_263), .B(n_346), .Y(n_423) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_265), .B(n_313), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_265), .B(n_274), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_265), .B(n_288), .Y(n_417) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g339 ( .A(n_269), .Y(n_339) );
AND2x2_ASAP7_75t_L g314 ( .A(n_270), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g392 ( .A(n_270), .Y(n_392) );
AND2x2_ASAP7_75t_L g324 ( .A(n_271), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_271), .B(n_294), .Y(n_340) );
AND2x2_ASAP7_75t_L g404 ( .A(n_271), .B(n_330), .Y(n_404) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g313 ( .A(n_275), .B(n_282), .Y(n_313) );
AND2x2_ASAP7_75t_L g409 ( .A(n_276), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_278), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_279), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_279), .B(n_286), .Y(n_374) );
AND2x2_ASAP7_75t_L g394 ( .A(n_279), .B(n_294), .Y(n_394) );
AND2x2_ASAP7_75t_L g415 ( .A(n_279), .B(n_359), .Y(n_415) );
OAI32xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_284), .A3(n_286), .B1(n_287), .B2(n_290), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_SL g288 ( .A(n_282), .Y(n_288) );
NAND2x1_ASAP7_75t_L g329 ( .A(n_282), .B(n_312), .Y(n_329) );
OR2x2_ASAP7_75t_L g333 ( .A(n_282), .B(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_282), .B(n_381), .Y(n_434) );
INVx1_ASAP7_75t_L g302 ( .A(n_283), .Y(n_302) );
OAI221xp5_ASAP7_75t_SL g420 ( .A1(n_284), .A2(n_375), .B1(n_421), .B2(n_424), .C(n_425), .Y(n_420) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g292 ( .A(n_285), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g335 ( .A(n_285), .B(n_308), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_285), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g413 ( .A(n_285), .B(n_346), .Y(n_413) );
INVxp67_ASAP7_75t_L g349 ( .A(n_286), .Y(n_349) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
AND2x2_ASAP7_75t_L g419 ( .A(n_288), .B(n_406), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_288), .B(n_369), .Y(n_442) );
INVx1_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_290), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g435 ( .A(n_290), .B(n_436), .Y(n_435) );
OAI21xp5_ASAP7_75t_SL g291 ( .A1(n_292), .A2(n_295), .B(n_298), .Y(n_291) );
AND2x2_ASAP7_75t_L g304 ( .A(n_293), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g388 ( .A(n_297), .B(n_308), .Y(n_388) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x2_ASAP7_75t_L g406 ( .A(n_299), .B(n_364), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_299), .B(n_363), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_300), .B(n_312), .Y(n_386) );
OAI211xp5_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_303), .B(n_306), .C(n_316), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_302), .A2(n_337), .B1(n_341), .B2(n_344), .C(n_347), .Y(n_336) );
AOI31xp33_ASAP7_75t_L g431 ( .A1(n_302), .A2(n_432), .A3(n_433), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_310), .B1(n_312), .B2(n_314), .Y(n_306) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g432 ( .A(n_312), .Y(n_432) );
INVx1_ASAP7_75t_L g395 ( .A(n_313), .Y(n_395) );
O2A1O1Ixp33_ASAP7_75t_L g438 ( .A1(n_315), .A2(n_439), .B(n_441), .C(n_443), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_320), .B2(n_324), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_321), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI221xp5_ASAP7_75t_SL g411 ( .A1(n_323), .A2(n_357), .B1(n_376), .B2(n_412), .C(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g407 ( .A(n_324), .Y(n_407) );
INVx1_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
NAND3xp33_ASAP7_75t_SL g326 ( .A(n_327), .B(n_336), .C(n_351), .Y(n_326) );
OAI21xp33_ASAP7_75t_L g377 ( .A1(n_328), .A2(n_378), .B(n_382), .Y(n_377) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_330), .B(n_430), .Y(n_429) );
INVxp67_ASAP7_75t_L g437 ( .A(n_331), .Y(n_437) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g375 ( .A(n_338), .B(n_358), .Y(n_375) );
INVx1_ASAP7_75t_L g350 ( .A(n_339), .Y(n_350) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVx1_ASAP7_75t_L g348 ( .A(n_342), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_342), .B(n_380), .Y(n_379) );
NOR4xp25_ASAP7_75t_L g347 ( .A(n_343), .B(n_348), .C(n_349), .D(n_350), .Y(n_347) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AOI222xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_356), .B1(n_362), .B2(n_363), .C1(n_365), .C2(n_369), .Y(n_351) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g449 ( .A(n_353), .Y(n_449) );
INVx1_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_365), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_370), .A2(n_426), .B(n_428), .Y(n_425) );
NOR4xp25_ASAP7_75t_L g371 ( .A(n_372), .B(n_383), .C(n_396), .D(n_411), .Y(n_371) );
OAI221xp5_ASAP7_75t_SL g372 ( .A1(n_373), .A2(n_374), .B1(n_375), .B2(n_376), .C(n_377), .Y(n_372) );
INVx1_ASAP7_75t_L g452 ( .A(n_373), .Y(n_452) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_380), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_SL g380 ( .A(n_381), .Y(n_380) );
OAI222xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B1(n_389), .B2(n_390), .C1(n_393), .C2(n_395), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI211xp5_ASAP7_75t_L g418 ( .A1(n_388), .A2(n_419), .B(n_420), .C(n_431), .Y(n_418) );
OR2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_402), .B1(n_403), .B2(n_405), .C1(n_407), .C2(n_408), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_413), .A2(n_416), .B1(n_449), .B2(n_450), .Y(n_448) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g443 ( .A1(n_444), .A2(n_446), .B(n_448), .C(n_451), .Y(n_443) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2x2_ASAP7_75t_L g772 ( .A(n_459), .B(n_476), .Y(n_772) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_462), .A2(n_464), .B(n_773), .Y(n_463) );
XNOR2xp5_ASAP7_75t_L g465 ( .A(n_466), .B(n_475), .Y(n_465) );
INVx1_ASAP7_75t_L g474 ( .A(n_468), .Y(n_474) );
INVx1_ASAP7_75t_L g472 ( .A(n_469), .Y(n_472) );
INVx2_ASAP7_75t_L g769 ( .A(n_476), .Y(n_769) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_SL g478 ( .A(n_479), .B(n_735), .Y(n_478) );
NOR3xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_639), .C(n_723), .Y(n_479) );
NAND4xp25_ASAP7_75t_L g480 ( .A(n_481), .B(n_582), .C(n_604), .D(n_620), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_520), .B1(n_543), .B2(n_561), .C(n_568), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_500), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_484), .B(n_561), .Y(n_594) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_484), .B(n_622), .C(n_635), .D(n_637), .Y(n_634) );
INVxp67_ASAP7_75t_L g751 ( .A(n_484), .Y(n_751) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OR2x2_ASAP7_75t_L g633 ( .A(n_485), .B(n_571), .Y(n_633) );
AND2x2_ASAP7_75t_L g657 ( .A(n_485), .B(n_500), .Y(n_657) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g624 ( .A(n_486), .B(n_560), .Y(n_624) );
AND2x2_ASAP7_75t_L g664 ( .A(n_486), .B(n_645), .Y(n_664) );
AND2x2_ASAP7_75t_L g681 ( .A(n_486), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_486), .B(n_501), .Y(n_705) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g559 ( .A(n_487), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g576 ( .A(n_487), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g588 ( .A(n_487), .B(n_501), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_487), .B(n_510), .Y(n_610) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_496), .B(n_497), .C(n_498), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_498), .A2(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g591 ( .A(n_500), .B(n_592), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_500), .A2(n_641), .B1(n_644), .B2(n_646), .C(n_650), .Y(n_640) );
AND2x2_ASAP7_75t_L g699 ( .A(n_500), .B(n_664), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_500), .B(n_681), .Y(n_733) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
INVx3_ASAP7_75t_L g560 ( .A(n_501), .Y(n_560) );
AND2x2_ASAP7_75t_L g608 ( .A(n_501), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g662 ( .A(n_501), .B(n_577), .Y(n_662) );
AND2x2_ASAP7_75t_L g720 ( .A(n_501), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g561 ( .A(n_510), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g577 ( .A(n_510), .Y(n_577) );
INVx1_ASAP7_75t_L g632 ( .A(n_510), .Y(n_632) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_510), .Y(n_638) );
AND2x2_ASAP7_75t_L g683 ( .A(n_510), .B(n_560), .Y(n_683) );
OR2x2_ASAP7_75t_L g722 ( .A(n_510), .B(n_562), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_515), .B(n_518), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_520), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_528), .Y(n_520) );
AND2x2_ASAP7_75t_L g718 ( .A(n_521), .B(n_715), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_521), .B(n_700), .Y(n_750) );
BUFx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g649 ( .A(n_522), .B(n_573), .Y(n_649) );
AND2x2_ASAP7_75t_L g698 ( .A(n_522), .B(n_546), .Y(n_698) );
INVx1_ASAP7_75t_L g744 ( .A(n_522), .Y(n_744) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_523), .Y(n_558) );
AND2x2_ASAP7_75t_L g599 ( .A(n_523), .B(n_573), .Y(n_599) );
INVx1_ASAP7_75t_L g616 ( .A(n_523), .Y(n_616) );
AND2x2_ASAP7_75t_L g622 ( .A(n_523), .B(n_539), .Y(n_622) );
AND2x2_ASAP7_75t_L g690 ( .A(n_528), .B(n_598), .Y(n_690) );
INVx2_ASAP7_75t_L g755 ( .A(n_528), .Y(n_755) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_539), .Y(n_528) );
AND2x2_ASAP7_75t_L g572 ( .A(n_529), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g585 ( .A(n_529), .B(n_547), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_529), .B(n_546), .Y(n_613) );
INVx1_ASAP7_75t_L g619 ( .A(n_529), .Y(n_619) );
INVx1_ASAP7_75t_L g636 ( .A(n_529), .Y(n_636) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_529), .Y(n_648) );
INVx2_ASAP7_75t_L g716 ( .A(n_529), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_534), .Y(n_531) );
INVx2_ASAP7_75t_L g573 ( .A(n_539), .Y(n_573) );
BUFx2_ASAP7_75t_L g670 ( .A(n_539), .Y(n_670) );
AND2x2_ASAP7_75t_L g715 ( .A(n_539), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_557), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_545), .B(n_652), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_545), .A2(n_714), .B(n_728), .Y(n_738) );
AND2x2_ASAP7_75t_L g763 ( .A(n_545), .B(n_649), .Y(n_763) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g685 ( .A(n_547), .Y(n_685) );
AND2x2_ASAP7_75t_L g714 ( .A(n_547), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_548), .Y(n_598) );
INVx2_ASAP7_75t_L g617 ( .A(n_548), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_548), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx2_ASAP7_75t_L g571 ( .A(n_558), .Y(n_571) );
OR2x2_ASAP7_75t_L g584 ( .A(n_558), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g652 ( .A(n_558), .B(n_648), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_558), .B(n_748), .Y(n_747) );
OR2x2_ASAP7_75t_L g753 ( .A(n_558), .B(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_558), .B(n_690), .Y(n_765) );
AND2x2_ASAP7_75t_L g644 ( .A(n_559), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g667 ( .A(n_559), .B(n_561), .Y(n_667) );
INVx2_ASAP7_75t_L g579 ( .A(n_560), .Y(n_579) );
AND2x2_ASAP7_75t_L g607 ( .A(n_560), .B(n_580), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_560), .B(n_632), .Y(n_688) );
AND2x2_ASAP7_75t_L g602 ( .A(n_561), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g749 ( .A(n_561), .Y(n_749) );
AND2x2_ASAP7_75t_L g761 ( .A(n_561), .B(n_624), .Y(n_761) );
AND2x2_ASAP7_75t_L g587 ( .A(n_562), .B(n_577), .Y(n_587) );
INVx1_ASAP7_75t_L g682 ( .A(n_562), .Y(n_682) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x4_ASAP7_75t_L g580 ( .A(n_567), .B(n_581), .Y(n_580) );
INVxp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_574), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_571), .B(n_618), .Y(n_627) );
OR2x2_ASAP7_75t_L g759 ( .A(n_571), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g676 ( .A(n_572), .B(n_617), .Y(n_676) );
AND2x2_ASAP7_75t_L g684 ( .A(n_572), .B(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g743 ( .A(n_572), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g767 ( .A(n_572), .B(n_614), .Y(n_767) );
NOR2xp67_ASAP7_75t_L g725 ( .A(n_573), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g754 ( .A(n_573), .B(n_617), .Y(n_754) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
AND2x2_ASAP7_75t_L g606 ( .A(n_576), .B(n_607), .Y(n_606) );
INVxp67_ASAP7_75t_L g768 ( .A(n_576), .Y(n_768) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx1_ASAP7_75t_L g603 ( .A(n_579), .Y(n_603) );
AND2x2_ASAP7_75t_L g654 ( .A(n_579), .B(n_587), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_579), .B(n_722), .Y(n_748) );
INVx2_ASAP7_75t_L g593 ( .A(n_580), .Y(n_593) );
INVx3_ASAP7_75t_L g645 ( .A(n_580), .Y(n_645) );
OR2x2_ASAP7_75t_L g673 ( .A(n_580), .B(n_674), .Y(n_673) );
AOI311xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_586), .A3(n_588), .B(n_589), .C(n_600), .Y(n_582) );
O2A1O1Ixp33_ASAP7_75t_L g620 ( .A1(n_583), .A2(n_621), .B(n_623), .C(n_625), .Y(n_620) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_SL g605 ( .A(n_585), .Y(n_605) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g623 ( .A(n_587), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_587), .B(n_603), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_587), .B(n_588), .Y(n_756) );
AND2x2_ASAP7_75t_L g678 ( .A(n_588), .B(n_592), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_594), .B(n_595), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g736 ( .A(n_592), .B(n_624), .Y(n_736) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_593), .B(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g630 ( .A(n_593), .Y(n_630) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
AND2x2_ASAP7_75t_L g621 ( .A(n_597), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g666 ( .A(n_599), .Y(n_666) );
AND2x4_ASAP7_75t_L g728 ( .A(n_599), .B(n_697), .Y(n_728) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_602), .A2(n_668), .B1(n_680), .B2(n_684), .C1(n_686), .C2(n_690), .Y(n_679) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B(n_608), .C(n_611), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_605), .B(n_649), .Y(n_672) );
INVx1_ASAP7_75t_L g694 ( .A(n_607), .Y(n_694) );
INVx1_ASAP7_75t_L g628 ( .A(n_609), .Y(n_628) );
OR2x2_ASAP7_75t_L g693 ( .A(n_610), .B(n_694), .Y(n_693) );
OAI21xp33_ASAP7_75t_SL g611 ( .A1(n_612), .A2(n_614), .B(n_618), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_612), .B(n_630), .C(n_631), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_612), .A2(n_649), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_616), .Y(n_669) );
AND2x2_ASAP7_75t_SL g635 ( .A(n_617), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g726 ( .A(n_617), .Y(n_726) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_617), .Y(n_742) );
INVx2_ASAP7_75t_L g700 ( .A(n_618), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_622), .B(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g674 ( .A(n_624), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B1(n_629), .B2(n_633), .C(n_634), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_628), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_SL g762 ( .A(n_628), .Y(n_762) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g643 ( .A(n_635), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_635), .B(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g701 ( .A(n_635), .B(n_649), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_635), .B(n_711), .Y(n_710) );
AND2x2_ASAP7_75t_L g734 ( .A(n_635), .B(n_669), .Y(n_734) );
BUFx3_ASAP7_75t_L g697 ( .A(n_636), .Y(n_697) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND5xp2_ASAP7_75t_L g639 ( .A(n_640), .B(n_658), .C(n_679), .D(n_691), .E(n_706), .Y(n_639) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AOI32xp33_ASAP7_75t_L g731 ( .A1(n_643), .A2(n_670), .A3(n_686), .B1(n_732), .B2(n_734), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_645), .B(n_704), .Y(n_703) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g655 ( .A(n_649), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_665), .B1(n_667), .B2(n_668), .C(n_671), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g660 ( .A(n_661), .B(n_663), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g730 ( .A(n_662), .B(n_681), .Y(n_730) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g745 ( .A1(n_667), .A2(n_728), .B1(n_746), .B2(n_751), .C(n_752), .Y(n_745) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g711 ( .A(n_670), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_673), .B1(n_675), .B2(n_677), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
INVx1_ASAP7_75t_L g689 ( .A(n_681), .Y(n_689) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OR2x2_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
AOI222xp33_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_695), .B1(n_699), .B2(n_700), .C1(n_701), .C2(n_702), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g746 ( .A1(n_700), .A2(n_747), .B1(n_749), .B2(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_SL g704 ( .A(n_705), .Y(n_704) );
AOI21xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_713), .A2(n_717), .B(n_719), .Y(n_712) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g760 ( .A(n_715), .Y(n_760) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_724), .A2(n_727), .B(n_729), .C(n_731), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI211xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_737), .B(n_739), .C(n_764), .Y(n_735) );
CKINVDCx16_ASAP7_75t_R g740 ( .A(n_736), .Y(n_740) );
INVxp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI211xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_745), .C(n_757), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
AOI21xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_755), .B(n_756), .Y(n_752) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_761), .B1(n_762), .B2(n_763), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
AOI21xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B(n_768), .Y(n_764) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
endmodule