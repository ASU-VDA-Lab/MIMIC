module real_jpeg_4475_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_1),
.A2(n_22),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_1),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_1),
.A2(n_36),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_1),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_151),
.B1(n_214),
.B2(n_217),
.Y(n_213)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_1),
.A2(n_253),
.B(n_256),
.C(n_259),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_1),
.B(n_267),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_1),
.B(n_55),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_1),
.B(n_75),
.C(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_1),
.B(n_112),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_1),
.B(n_108),
.C(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_1),
.B(n_29),
.Y(n_327)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_2),
.A2(n_78),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_2),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_2),
.A2(n_83),
.B1(n_114),
.B2(n_118),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_2),
.A2(n_26),
.B1(n_83),
.B2(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_2),
.A2(n_83),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_3),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_3),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_3),
.A2(n_89),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_3),
.A2(n_89),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_3),
.A2(n_89),
.B1(n_194),
.B2(n_198),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_4),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_5),
.Y(n_405)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_6),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_7),
.Y(n_267)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_8),
.Y(n_255)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_10),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_10),
.A2(n_24),
.B1(n_143),
.B2(n_146),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_10),
.A2(n_24),
.B1(n_183),
.B2(n_187),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_10),
.A2(n_24),
.B1(n_164),
.B2(n_265),
.Y(n_264)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_11),
.Y(n_261)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_12),
.Y(n_403)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_13),
.Y(n_75)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_402),
.B(n_404),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_131),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_129),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_18),
.B(n_126),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.C(n_124),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_19),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.C(n_84),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_20),
.A2(n_177),
.B1(n_178),
.B2(n_189),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_20),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_20),
.B(n_138),
.C(n_178),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_20),
.B(n_234),
.C(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_20),
.A2(n_189),
.B1(n_234),
.B2(n_328),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_20),
.A2(n_189),
.B1(n_374),
.B2(n_375),
.Y(n_373)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g222 ( 
.A1(n_21),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_222)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_28),
.A2(n_48),
.B1(n_51),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_28),
.A2(n_51),
.B1(n_121),
.B2(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_28),
.A2(n_48),
.B(n_51),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_30),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_31),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_31),
.Y(n_181)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_36),
.Y(n_258)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_44),
.B2(n_46),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_45),
.Y(n_122)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_52),
.A2(n_84),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_52),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_52),
.B(n_222),
.C(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_52),
.A2(n_377),
.B1(n_379),
.B2(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_80),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_53),
.B(n_148),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_68),
.Y(n_53)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_54),
.A2(n_68),
.B1(n_141),
.B2(n_147),
.Y(n_140)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_55),
.A2(n_193),
.B(n_199),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_55),
.B(n_142),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_55),
.A2(n_69),
.B1(n_80),
.B2(n_193),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_59),
.B1(n_62),
.B2(n_66),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g160 ( 
.A(n_61),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_61),
.Y(n_216)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_65),
.Y(n_172)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_69),
.B(n_148),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_72),
.Y(n_145)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_72),
.Y(n_291)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_82),
.Y(n_198)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_84),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_91),
.B1(n_112),
.B2(n_113),
.Y(n_84)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_85),
.Y(n_380)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_88),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_91),
.B(n_221),
.Y(n_381)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_103),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_92),
.A2(n_103),
.B1(n_179),
.B2(n_182),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g234 ( 
.A1(n_92),
.A2(n_103),
.B1(n_179),
.B2(n_182),
.Y(n_234)
);

NAND2x1_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_98),
.B1(n_100),
.B2(n_102),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_99),
.Y(n_310)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_103),
.A2(n_380),
.B(n_381),
.Y(n_379)
);

AOI22x1_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_106),
.Y(n_312)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_120),
.B(n_124),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_125),
.B(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_397),
.B(n_401),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_368),
.B(n_394),
.Y(n_132)
);

OAI211xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_268),
.B(n_362),
.C(n_367),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_239),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g362 ( 
.A1(n_135),
.A2(n_239),
.B(n_363),
.C(n_366),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_223),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_136),
.B(n_223),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_190),
.C(n_206),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_137),
.B(n_190),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_176),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_156),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_139),
.A2(n_140),
.B1(n_156),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_139),
.A2(n_140),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_139),
.A2(n_140),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_140),
.B(n_263),
.C(n_300),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_140),
.B(n_320),
.C(n_322),
.Y(n_333)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_162),
.B1(n_167),
.B2(n_173),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_163),
.A2(n_213),
.B1(n_264),
.B2(n_267),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_163),
.A2(n_213),
.B1(n_264),
.B2(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_164),
.Y(n_279)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_168),
.B(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_170),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_170),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_177),
.A2(n_178),
.B1(n_218),
.B2(n_289),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_177),
.B(n_289),
.C(n_307),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_177),
.A2(n_178),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_178),
.B(n_222),
.C(n_338),
.Y(n_355)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_180),
.A2(n_254),
.B(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_201),
.B2(n_205),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_201),
.Y(n_230)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_201),
.A2(n_205),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_201),
.A2(n_229),
.B(n_230),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_202),
.B(n_213),
.Y(n_313)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_203),
.Y(n_282)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_220),
.C(n_222),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_218),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_209),
.A2(n_218),
.B1(n_289),
.B2(n_354),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_216),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_218),
.A2(n_289),
.B1(n_290),
.B2(n_294),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_222),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_222),
.A2(n_246),
.B1(n_336),
.B2(n_337),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_222),
.A2(n_246),
.B1(n_372),
.B2(n_373),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_222),
.A2(n_246),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_222),
.B(n_373),
.C(n_378),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_237),
.B2(n_238),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_231),
.B1(n_232),
.B2(n_236),
.Y(n_225)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_231),
.B(n_236),
.C(n_238),
.Y(n_393)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_234),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_234),
.A2(n_324),
.B1(n_325),
.B2(n_328),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_234),
.Y(n_328)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_235),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_235),
.A2(n_383),
.B1(n_387),
.B2(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_240),
.B(n_242),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_248),
.C(n_250),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_244),
.B(n_248),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_250),
.B(n_361),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_251),
.B(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_262),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_252),
.A2(n_262),
.B1(n_263),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_252),
.Y(n_345)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_262),
.A2(n_263),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_263),
.B(n_284),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_284),
.Y(n_285)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_347),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_332),
.B(n_346),
.Y(n_269)
);

AOI21x1_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_317),
.B(n_331),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_272),
.A2(n_304),
.B(n_316),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_296),
.B(n_303),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_286),
.B(n_295),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_283),
.B(n_285),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_281),
.A2(n_287),
.B1(n_326),
.B2(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_288),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_326),
.C(n_328),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_294),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_290),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_305),
.B(n_306),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_315),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_313),
.B2(n_314),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_314),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_330),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_318),
.B(n_330),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_322),
.B1(n_323),
.B2(n_329),
.Y(n_318)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_333),
.B(n_334),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_340),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_342),
.C(n_343),
.Y(n_356)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_357),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_349),
.B(n_356),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_356),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_350),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_355),
.C(n_359),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_357),
.A2(n_364),
.B(n_365),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_360),
.Y(n_357)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_358),
.B(n_360),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_389),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_369),
.A2(n_395),
.B(n_396),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_382),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_382),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_378),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_387),
.C(n_388),
.Y(n_382)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_393),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_393),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_398),
.B(n_400),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_402),
.B(n_405),
.Y(n_404)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);


endmodule