module fake_jpeg_31044_n_180 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_180);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_6),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_40),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_1),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_81),
.Y(n_94)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_58),
.C(n_53),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_96),
.Y(n_102)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_44),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_88),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_95),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_63),
.B(n_69),
.C(n_62),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_96),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_67),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_44),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_64),
.B1(n_54),
.B2(n_52),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_108),
.B1(n_113),
.B2(n_45),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_5),
.Y(n_133)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_110),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_64),
.B1(n_52),
.B2(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_71),
.Y(n_110)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_111),
.A2(n_8),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_83),
.B(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_114),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_70),
.B1(n_68),
.B2(n_46),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_4),
.Y(n_132)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_61),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_2),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_59),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_1),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_122),
.B1(n_20),
.B2(n_21),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_111),
.A2(n_57),
.B1(n_56),
.B2(n_55),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_101),
.A2(n_55),
.B1(n_2),
.B2(n_4),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_114),
.A2(n_98),
.B1(n_101),
.B2(n_99),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_30),
.B(n_33),
.C(n_34),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_55),
.B1(n_5),
.B2(n_7),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

FAx1_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_141),
.CI(n_29),
.CON(n_158),
.SN(n_158)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_110),
.B(n_10),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_140),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_11),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_110),
.B(n_14),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_16),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_19),
.Y(n_142)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_146),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_137),
.Y(n_146)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_24),
.B(n_28),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_151),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_158),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_159),
.A2(n_123),
.B1(n_125),
.B2(n_128),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_121),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_148),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_167),
.B(n_154),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_152),
.A2(n_142),
.A3(n_127),
.B1(n_132),
.B2(n_135),
.C1(n_41),
.C2(n_42),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_171),
.B1(n_162),
.B2(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

AOI222xp33_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_159),
.B1(n_161),
.B2(n_149),
.C1(n_160),
.C2(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_159),
.C(n_173),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_150),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_144),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_144),
.B(n_164),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_168),
.Y(n_180)
);


endmodule