module real_aes_676_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_635;
wire n_792;
wire n_287;
wire n_386;
wire n_673;
wire n_518;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_656;
wire n_532;
wire n_316;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_782;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_799;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_475;
wire n_554;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_0), .A2(n_145), .B1(n_477), .B2(n_478), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g515 ( .A1(n_1), .A2(n_3), .B1(n_328), .B2(n_398), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_2), .A2(n_767), .B1(n_768), .B2(n_785), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_2), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_4), .A2(n_268), .B1(n_408), .B2(n_633), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_5), .A2(n_80), .B1(n_394), .B2(n_395), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_6), .A2(n_87), .B1(n_415), .B2(n_503), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_7), .A2(n_60), .B1(n_321), .B2(n_394), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_8), .A2(n_97), .B1(n_413), .B2(n_506), .Y(n_505) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_9), .A2(n_197), .B1(n_299), .B2(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g761 ( .A(n_9), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_10), .A2(n_167), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_11), .A2(n_240), .B1(n_394), .B2(n_395), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_12), .A2(n_19), .B1(n_405), .B2(n_406), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_13), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_14), .A2(n_180), .B1(n_406), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_15), .A2(n_35), .B1(n_416), .B2(n_496), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_16), .A2(n_139), .B1(n_481), .B2(n_488), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g743 ( .A1(n_17), .A2(n_245), .B1(n_467), .B2(n_472), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g366 ( .A(n_18), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_20), .B(n_293), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_21), .A2(n_234), .B1(n_477), .B2(n_478), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g495 ( .A1(n_22), .A2(n_148), .B1(n_410), .B2(n_496), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_23), .A2(n_129), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22x1_ASAP7_75t_L g728 ( .A1(n_24), .A2(n_131), .B1(n_368), .B2(n_481), .Y(n_728) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_25), .A2(n_69), .B1(n_299), .B2(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_25), .B(n_760), .Y(n_759) );
AO222x2_ASAP7_75t_L g466 ( .A1(n_26), .A2(n_68), .B1(n_216), .B2(n_427), .C1(n_467), .C2(n_468), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_27), .A2(n_199), .B1(n_371), .B2(n_415), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_28), .A2(n_33), .B1(n_560), .B2(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_SL g476 ( .A1(n_29), .A2(n_217), .B1(n_477), .B2(n_478), .Y(n_476) );
AOI22xp33_ASAP7_75t_SL g497 ( .A1(n_30), .A2(n_101), .B1(n_498), .B2(n_500), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_31), .A2(n_202), .B1(n_394), .B2(n_545), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_32), .A2(n_146), .B1(n_468), .B2(n_560), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_34), .A2(n_249), .B1(n_480), .B2(n_484), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_36), .A2(n_220), .B1(n_529), .B2(n_530), .Y(n_652) );
INVx1_ASAP7_75t_L g311 ( .A(n_37), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_38), .A2(n_223), .B1(n_542), .B2(n_543), .Y(n_541) );
XNOR2xp5_ASAP7_75t_L g712 ( .A(n_39), .B(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_40), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_41), .A2(n_45), .B1(n_481), .B2(n_488), .Y(n_751) );
AOI222xp33_ASAP7_75t_L g783 ( .A1(n_42), .A2(n_61), .B1(n_159), .B2(n_427), .C1(n_696), .C2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g473 ( .A1(n_43), .A2(n_226), .B1(n_432), .B2(n_433), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_44), .A2(n_170), .B1(n_678), .B2(n_679), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_46), .A2(n_128), .B1(n_481), .B2(n_488), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_47), .A2(n_238), .B1(n_372), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_48), .A2(n_118), .B1(n_485), .B2(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_49), .B(n_547), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_50), .A2(n_250), .B1(n_467), .B2(n_585), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_51), .A2(n_186), .B1(n_467), .B2(n_472), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_52), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_53), .A2(n_259), .B1(n_342), .B2(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g509 ( .A(n_54), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_55), .A2(n_267), .B1(n_444), .B2(n_445), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_56), .A2(n_166), .B1(n_532), .B2(n_681), .Y(n_680) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_57), .A2(n_114), .B1(n_471), .B2(n_472), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_58), .A2(n_136), .B1(n_444), .B2(n_681), .Y(n_775) );
CKINVDCx20_ASAP7_75t_R g718 ( .A(n_59), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_62), .A2(n_230), .B1(n_328), .B2(n_332), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_63), .A2(n_212), .B1(n_430), .B2(n_433), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_64), .A2(n_151), .B1(n_450), .B2(n_451), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_65), .A2(n_78), .B1(n_401), .B2(n_517), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_66), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_67), .A2(n_179), .B1(n_527), .B2(n_782), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_70), .A2(n_109), .B1(n_468), .B2(n_471), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g392 ( .A(n_71), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g531 ( .A1(n_72), .A2(n_126), .B1(n_445), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_73), .A2(n_244), .B1(n_415), .B2(n_633), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_74), .A2(n_174), .B1(n_480), .B2(n_481), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_75), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_76), .A2(n_237), .B1(n_484), .B2(n_485), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_77), .A2(n_193), .B1(n_534), .B2(n_535), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g747 ( .A1(n_79), .A2(n_233), .B1(n_477), .B2(n_478), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_81), .A2(n_130), .B1(n_471), .B2(n_699), .Y(n_698) );
OAI22x1_ASAP7_75t_L g791 ( .A1(n_82), .A2(n_769), .B1(n_792), .B2(n_793), .Y(n_791) );
CKINVDCx16_ASAP7_75t_R g793 ( .A(n_82), .Y(n_793) );
INVx3_ASAP7_75t_L g299 ( .A(n_83), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_84), .A2(n_156), .B1(n_487), .B2(n_488), .Y(n_486) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_85), .A2(n_164), .B1(n_400), .B2(n_401), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_86), .A2(n_198), .B1(n_415), .B2(n_416), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_88), .A2(n_177), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_89), .A2(n_133), .B1(n_485), .B2(n_487), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_90), .A2(n_135), .B1(n_400), .B2(n_543), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_91), .A2(n_253), .B1(n_413), .B2(n_506), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_92), .A2(n_147), .B1(n_410), .B2(n_496), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_93), .A2(n_190), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_94), .A2(n_191), .B1(n_437), .B2(n_539), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_95), .A2(n_181), .B1(n_328), .B2(n_332), .Y(n_771) );
OA22x2_ASAP7_75t_L g521 ( .A1(n_96), .A2(n_522), .B1(n_523), .B2(n_548), .Y(n_521) );
INVxp67_ASAP7_75t_L g548 ( .A(n_96), .Y(n_548) );
OA22x2_ASAP7_75t_L g597 ( .A1(n_96), .A2(n_522), .B1(n_523), .B2(n_548), .Y(n_597) );
XNOR2x1_ASAP7_75t_L g551 ( .A(n_98), .B(n_552), .Y(n_551) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_99), .A2(n_203), .B1(n_228), .B2(n_313), .C1(n_547), .C2(n_687), .Y(n_686) );
AO222x2_ASAP7_75t_L g741 ( .A1(n_100), .A2(n_150), .B1(n_173), .B2(n_427), .C1(n_432), .C2(n_696), .Y(n_741) );
OAI22x1_ASAP7_75t_L g621 ( .A1(n_102), .A2(n_622), .B1(n_634), .B2(n_635), .Y(n_621) );
INVx1_ASAP7_75t_L g635 ( .A(n_102), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_103), .A2(n_183), .B1(n_478), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_104), .A2(n_153), .B1(n_471), .B2(n_699), .Y(n_744) );
INVx1_ASAP7_75t_SL g300 ( .A(n_105), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_105), .B(n_140), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_106), .A2(n_169), .B1(n_357), .B2(n_444), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_107), .Y(n_717) );
INVx2_ASAP7_75t_L g279 ( .A(n_108), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_110), .A2(n_185), .B1(n_451), .B2(n_777), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_111), .A2(n_227), .B1(n_408), .B2(n_410), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_112), .A2(n_260), .B1(n_413), .B2(n_573), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_113), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g435 ( .A1(n_115), .A2(n_123), .B1(n_436), .B2(n_437), .Y(n_435) );
OA22x2_ASAP7_75t_L g637 ( .A1(n_116), .A2(n_638), .B1(n_660), .B2(n_661), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_116), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_117), .A2(n_261), .B1(n_371), .B2(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_119), .A2(n_246), .B1(n_485), .B2(n_487), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_120), .A2(n_195), .B1(n_444), .B2(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_121), .B(n_547), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_122), .A2(n_142), .B1(n_413), .B2(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_124), .B(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_125), .A2(n_218), .B1(n_368), .B2(n_447), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_127), .A2(n_272), .B(n_280), .C(n_765), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g593 ( .A(n_132), .Y(n_593) );
OA22x2_ASAP7_75t_L g287 ( .A1(n_134), .A2(n_288), .B1(n_289), .B2(n_384), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_134), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_137), .A2(n_270), .B1(n_585), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_138), .A2(n_144), .B1(n_529), .B2(n_530), .Y(n_528) );
AO22x2_ASAP7_75t_L g302 ( .A1(n_140), .A2(n_207), .B1(n_299), .B2(n_303), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g452 ( .A1(n_141), .A2(n_222), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_143), .A2(n_158), .B1(n_328), .B2(n_398), .Y(n_397) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_149), .A2(n_163), .B1(n_437), .B2(n_539), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_152), .A2(n_236), .B1(n_416), .B2(n_529), .Y(n_606) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_154), .A2(n_215), .B1(n_400), .B2(n_518), .Y(n_647) );
INVx1_ASAP7_75t_L g301 ( .A(n_155), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_157), .A2(n_224), .B1(n_432), .B2(n_696), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_160), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_161), .A2(n_211), .B1(n_408), .B2(n_608), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g748 ( .A1(n_162), .A2(n_178), .B1(n_480), .B2(n_484), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_165), .A2(n_208), .B1(n_439), .B2(n_440), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_168), .A2(n_192), .B1(n_357), .B2(n_444), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g355 ( .A(n_171), .Y(n_355) );
INVx1_ASAP7_75t_L g422 ( .A(n_172), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_175), .A2(n_188), .B1(n_394), .B2(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_176), .B(n_321), .Y(n_320) );
CKINVDCx20_ASAP7_75t_R g380 ( .A(n_182), .Y(n_380) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_184), .A2(n_225), .B1(n_368), .B2(n_453), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_187), .A2(n_205), .B1(n_394), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_189), .A2(n_213), .B1(n_467), .B2(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_194), .B(n_511), .Y(n_624) );
CKINVDCx16_ASAP7_75t_R g710 ( .A(n_196), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_200), .A2(n_262), .B1(n_371), .B2(n_685), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_201), .A2(n_491), .B1(n_492), .B2(n_519), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_201), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_204), .A2(n_219), .B1(n_480), .B2(n_488), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_206), .A2(n_463), .B1(n_464), .B2(n_489), .Y(n_462) );
INVx1_ASAP7_75t_L g489 ( .A(n_206), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_209), .A2(n_266), .B1(n_371), .B2(n_373), .C(n_376), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_210), .A2(n_257), .B1(n_432), .B2(n_433), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_214), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g757 ( .A(n_214), .Y(n_757) );
INVx1_ASAP7_75t_L g276 ( .A(n_221), .Y(n_276) );
AND2x2_ASAP7_75t_R g787 ( .A(n_221), .B(n_757), .Y(n_787) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_229), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_231), .A2(n_254), .B1(n_338), .B2(n_342), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_232), .A2(n_265), .B1(n_328), .B2(n_398), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_235), .A2(n_255), .B1(n_394), .B2(n_395), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_239), .B(n_278), .Y(n_277) );
AO22x2_ASAP7_75t_L g603 ( .A1(n_241), .A2(n_604), .B1(n_617), .B2(n_618), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_241), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_242), .B(n_391), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_243), .A2(n_264), .B1(n_328), .B2(n_398), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_247), .B(n_427), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_248), .A2(n_269), .B1(n_485), .B2(n_708), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_251), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_252), .Y(n_561) );
XNOR2x1_ASAP7_75t_L g386 ( .A(n_256), .B(n_387), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_258), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_263), .Y(n_558) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_274), .B(n_277), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g799 ( .A(n_275), .B(n_277), .Y(n_799) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_276), .B(n_757), .Y(n_756) );
OAI32xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_600), .A3(n_754), .B1(n_763), .B2(n_764), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_520), .B2(n_599), .Y(n_281) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_282), .A2(n_283), .B1(n_520), .B2(n_599), .C(n_755), .Y(n_764) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_457), .B2(n_458), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_419), .B1(n_455), .B2(n_456), .Y(n_285) );
INVx1_ASAP7_75t_L g456 ( .A(n_286), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_385), .B1(n_417), .B2(n_418), .Y(n_286) );
INVx2_ASAP7_75t_L g417 ( .A(n_287), .Y(n_417) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND3x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_346), .C(n_370), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_291), .B(n_326), .Y(n_290) );
OAI221xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_311), .B1(n_312), .B2(n_319), .C(n_320), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx4_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx4_ASAP7_75t_SL g391 ( .A(n_294), .Y(n_391) );
INVx3_ASAP7_75t_SL g512 ( .A(n_294), .Y(n_512) );
INVx3_ASAP7_75t_L g547 ( .A(n_294), .Y(n_547) );
INVx6_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_304), .Y(n_295) );
AND2x4_ASAP7_75t_L g334 ( .A(n_296), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g344 ( .A(n_296), .B(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g427 ( .A(n_296), .B(n_304), .Y(n_427) );
AND2x2_ASAP7_75t_L g467 ( .A(n_296), .B(n_345), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_296), .B(n_335), .Y(n_468) );
AND2x2_ASAP7_75t_L g699 ( .A(n_296), .B(n_335), .Y(n_699) );
AND2x2_ASAP7_75t_L g773 ( .A(n_296), .B(n_345), .Y(n_773) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_302), .Y(n_296) );
AND2x2_ASAP7_75t_L g317 ( .A(n_297), .B(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_297), .Y(n_325) );
INVx2_ASAP7_75t_L g341 ( .A(n_297), .Y(n_341) );
OAI22x1_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_300), .B2(n_301), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g303 ( .A(n_299), .Y(n_303) );
INVx2_ASAP7_75t_L g307 ( .A(n_299), .Y(n_307) );
INVx1_ASAP7_75t_L g310 ( .A(n_299), .Y(n_310) );
INVx2_ASAP7_75t_L g318 ( .A(n_302), .Y(n_318) );
AND2x2_ASAP7_75t_L g340 ( .A(n_302), .B(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g358 ( .A(n_302), .Y(n_358) );
AND2x4_ASAP7_75t_L g364 ( .A(n_304), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g375 ( .A(n_304), .B(n_340), .Y(n_375) );
AND2x4_ASAP7_75t_L g379 ( .A(n_304), .B(n_317), .Y(n_379) );
AND2x2_ASAP7_75t_L g480 ( .A(n_304), .B(n_365), .Y(n_480) );
AND2x6_ASAP7_75t_L g481 ( .A(n_304), .B(n_340), .Y(n_481) );
AND2x2_ASAP7_75t_L g487 ( .A(n_304), .B(n_317), .Y(n_487) );
AND2x2_ASAP7_75t_L g708 ( .A(n_304), .B(n_317), .Y(n_708) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_308), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g316 ( .A(n_306), .B(n_308), .Y(n_316) );
AND2x2_ASAP7_75t_L g324 ( .A(n_306), .B(n_309), .Y(n_324) );
INVx1_ASAP7_75t_L g331 ( .A(n_306), .Y(n_331) );
INVxp67_ASAP7_75t_L g345 ( .A(n_308), .Y(n_345) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g330 ( .A(n_309), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx6f_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx5_ASAP7_75t_L g394 ( .A(n_315), .Y(n_394) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x4_ASAP7_75t_L g339 ( .A(n_316), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g369 ( .A(n_316), .B(n_365), .Y(n_369) );
AND2x4_ASAP7_75t_L g432 ( .A(n_316), .B(n_317), .Y(n_432) );
AND2x2_ASAP7_75t_L g472 ( .A(n_316), .B(n_340), .Y(n_472) );
AND2x2_ASAP7_75t_L g484 ( .A(n_316), .B(n_365), .Y(n_484) );
AND2x2_ASAP7_75t_L g585 ( .A(n_316), .B(n_340), .Y(n_585) );
AND2x2_ASAP7_75t_L g329 ( .A(n_317), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g471 ( .A(n_317), .B(n_330), .Y(n_471) );
AND2x4_ASAP7_75t_L g365 ( .A(n_318), .B(n_341), .Y(n_365) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_321), .Y(n_687) );
INVx3_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g545 ( .A(n_322), .Y(n_545) );
INVx2_ASAP7_75t_L g642 ( .A(n_322), .Y(n_642) );
INVx3_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx12f_ASAP7_75t_L g395 ( .A(n_323), .Y(n_395) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x4_ASAP7_75t_L g357 ( .A(n_324), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g372 ( .A(n_324), .B(n_365), .Y(n_372) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_324), .B(n_325), .Y(n_433) );
AND2x4_ASAP7_75t_L g478 ( .A(n_324), .B(n_358), .Y(n_478) );
AND2x4_ASAP7_75t_L g485 ( .A(n_324), .B(n_365), .Y(n_485) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_324), .B(n_325), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_337), .Y(n_326) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_329), .Y(n_436) );
INVx3_ASAP7_75t_L g540 ( .A(n_329), .Y(n_540) );
AND2x2_ASAP7_75t_L g354 ( .A(n_330), .B(n_340), .Y(n_354) );
AND2x4_ASAP7_75t_L g383 ( .A(n_330), .B(n_365), .Y(n_383) );
AND2x2_ASAP7_75t_SL g477 ( .A(n_330), .B(n_340), .Y(n_477) );
AND2x6_ASAP7_75t_L g488 ( .A(n_330), .B(n_365), .Y(n_488) );
AND2x2_ASAP7_75t_L g704 ( .A(n_330), .B(n_340), .Y(n_704) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_331), .Y(n_336) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx4f_ASAP7_75t_L g398 ( .A(n_334), .Y(n_398) );
BUFx6f_ASAP7_75t_SL g437 ( .A(n_334), .Y(n_437) );
BUFx3_ASAP7_75t_L g673 ( .A(n_334), .Y(n_673) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx4f_ASAP7_75t_SL g517 ( .A(n_338), .Y(n_517) );
INVx1_ASAP7_75t_L g565 ( .A(n_338), .Y(n_565) );
BUFx2_ASAP7_75t_L g675 ( .A(n_338), .Y(n_675) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx3_ASAP7_75t_L g400 ( .A(n_339), .Y(n_400) );
BUFx2_ASAP7_75t_L g439 ( .A(n_339), .Y(n_439) );
BUFx2_ASAP7_75t_L g542 ( .A(n_339), .Y(n_542) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_SL g401 ( .A(n_343), .Y(n_401) );
INVx2_ASAP7_75t_L g440 ( .A(n_343), .Y(n_440) );
INVx2_ASAP7_75t_SL g518 ( .A(n_343), .Y(n_518) );
INVx1_ASAP7_75t_L g543 ( .A(n_343), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_343), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_563) );
INVx6_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_359), .Y(n_346) );
OAI22xp33_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_355), .B2(n_356), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g405 ( .A(n_351), .Y(n_405) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g499 ( .A(n_352), .Y(n_499) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_352), .Y(n_532) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_354), .Y(n_444) );
BUFx3_ASAP7_75t_L g651 ( .A(n_354), .Y(n_651) );
INVx3_ASAP7_75t_L g406 ( .A(n_356), .Y(n_406) );
INVx2_ASAP7_75t_L g500 ( .A(n_356), .Y(n_500) );
INVx5_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
BUFx2_ASAP7_75t_L g445 ( .A(n_357), .Y(n_445) );
BUFx2_ASAP7_75t_L g681 ( .A(n_357), .Y(n_681) );
OAI22xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_361), .B1(n_366), .B2(n_367), .Y(n_359) );
INVx1_ASAP7_75t_L g678 ( .A(n_361), .Y(n_678) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_362), .Y(n_415) );
INVx4_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_SL g453 ( .A(n_363), .Y(n_453) );
INVx2_ASAP7_75t_SL g529 ( .A(n_363), .Y(n_529) );
INVx2_ASAP7_75t_L g782 ( .A(n_363), .Y(n_782) );
INVx8_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g679 ( .A(n_368), .Y(n_679) );
BUFx6f_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx3_ASAP7_75t_L g416 ( .A(n_369), .Y(n_416) );
INVx2_ASAP7_75t_L g504 ( .A(n_369), .Y(n_504) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_369), .Y(n_527) );
BUFx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g454 ( .A(n_372), .Y(n_454) );
BUFx2_ASAP7_75t_SL g506 ( .A(n_372), .Y(n_506) );
INVx2_ASAP7_75t_L g536 ( .A(n_372), .Y(n_536) );
BUFx3_ASAP7_75t_L g656 ( .A(n_372), .Y(n_656) );
BUFx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx3_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
BUFx2_ASAP7_75t_L g777 ( .A(n_375), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B1(n_380), .B2(n_381), .Y(n_376) );
INVx2_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
INVx3_ASAP7_75t_L g534 ( .A(n_378), .Y(n_534) );
INVx2_ASAP7_75t_L g655 ( .A(n_378), .Y(n_655) );
INVx2_ASAP7_75t_L g685 ( .A(n_378), .Y(n_685) );
INVx6_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx3_ASAP7_75t_L g447 ( .A(n_379), .Y(n_447) );
BUFx3_ASAP7_75t_L g780 ( .A(n_379), .Y(n_780) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_SL g410 ( .A(n_382), .Y(n_410) );
INVx2_ASAP7_75t_L g451 ( .A(n_382), .Y(n_451) );
INVx2_ASAP7_75t_L g530 ( .A(n_382), .Y(n_530) );
INVx1_ASAP7_75t_SL g608 ( .A(n_382), .Y(n_608) );
INVx2_ASAP7_75t_L g633 ( .A(n_382), .Y(n_633) );
INVx8_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g418 ( .A(n_385), .Y(n_418) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g387 ( .A(n_388), .B(n_402), .Y(n_387) );
NOR2xp67_ASAP7_75t_L g388 ( .A(n_389), .B(n_396), .Y(n_388) );
OAI21xp5_ASAP7_75t_SL g389 ( .A1(n_390), .A2(n_392), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVxp67_ASAP7_75t_L g562 ( .A(n_398), .Y(n_562) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_403), .B(n_411), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_407), .Y(n_403) );
INVx2_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx3_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
INVx2_ASAP7_75t_SL g496 ( .A(n_409), .Y(n_496) );
INVx2_ASAP7_75t_L g526 ( .A(n_409), .Y(n_526) );
INVx2_ASAP7_75t_L g658 ( .A(n_409), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g455 ( .A(n_419), .Y(n_455) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
XNOR2x1_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
NAND2x1_ASAP7_75t_L g423 ( .A(n_424), .B(n_441), .Y(n_423) );
NOR2xp67_ASAP7_75t_L g424 ( .A(n_425), .B(n_434), .Y(n_424) );
OAI21xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_428), .B(n_429), .Y(n_425) );
OAI222xp33_ASAP7_75t_L g715 ( .A1(n_426), .A2(n_431), .B1(n_716), .B2(n_717), .C1(n_718), .C2(n_719), .Y(n_715) );
INVx2_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_432), .Y(n_784) );
INVxp67_ASAP7_75t_L g719 ( .A(n_433), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_435), .B(n_438), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_448), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_452), .Y(n_448) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
XNOR2x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_490), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_465), .B(n_474), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_469), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_482), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_479), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_SL g519 ( .A(n_492), .Y(n_519) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_507), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_501), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g659 ( .A(n_504), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_514), .Y(n_507) );
OAI21xp33_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_513), .Y(n_508) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx6f_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_549), .B1(n_594), .B2(n_598), .Y(n_520) );
INVx2_ASAP7_75t_SL g522 ( .A(n_523), .Y(n_522) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_537), .Y(n_523) );
NAND4xp25_ASAP7_75t_SL g524 ( .A(n_525), .B(n_528), .C(n_531), .D(n_533), .Y(n_524) );
INVx1_ASAP7_75t_L g574 ( .A(n_527), .Y(n_574) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_SL g610 ( .A(n_536), .Y(n_610) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .C(n_544), .D(n_546), .Y(n_537) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g560 ( .A(n_540), .Y(n_560) );
INVx1_ASAP7_75t_L g598 ( .A(n_549), .Y(n_598) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
XOR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_576), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_567), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_557), .C(n_563), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_555), .B(n_556), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B1(n_561), .B2(n_562), .Y(n_557) );
INVx2_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_568), .B(n_571), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .Y(n_571) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
XOR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_593), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_578), .B(n_586), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_590), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g763 ( .A(n_600), .Y(n_763) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_663), .B1(n_752), .B2(n_753), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_602), .Y(n_752) );
XNOR2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_619), .Y(n_602) );
INVx1_ASAP7_75t_SL g618 ( .A(n_604), .Y(n_618) );
NOR2x1_ASAP7_75t_L g604 ( .A(n_605), .B(n_612), .Y(n_604) );
NAND4xp25_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .C(n_609), .D(n_611), .Y(n_605) );
NAND4xp25_ASAP7_75t_SL g612 ( .A(n_613), .B(n_614), .C(n_615), .D(n_616), .Y(n_612) );
AO22x2_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_636), .B2(n_637), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g634 ( .A(n_622), .Y(n_634) );
OR2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_628), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .C(n_626), .D(n_627), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_630), .C(n_631), .D(n_632), .Y(n_628) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_648), .Y(n_638) );
NOR3xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_644), .C(n_646), .Y(n_639) );
NOR4xp25_ASAP7_75t_L g661 ( .A(n_640), .B(n_649), .C(n_653), .D(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_645), .B(n_647), .Y(n_662) );
INVxp67_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_653), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g753 ( .A(n_663), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_665), .B1(n_734), .B2(n_735), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
AO22x2_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_711), .B1(n_730), .B2(n_731), .Y(n_665) );
INVx2_ASAP7_75t_SL g730 ( .A(n_666), .Y(n_730) );
OA22x2_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_689), .B2(n_690), .Y(n_666) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
XNOR2x1_ASAP7_75t_L g668 ( .A(n_669), .B(n_688), .Y(n_668) );
NAND4xp75_ASAP7_75t_L g669 ( .A(n_670), .B(n_676), .C(n_682), .D(n_686), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_674), .Y(n_670) );
BUFx6f_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_680), .Y(n_676) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
XOR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_710), .Y(n_690) );
NAND2x1p5_ASAP7_75t_L g691 ( .A(n_692), .B(n_701), .Y(n_691) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_697), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
NOR2x1_ASAP7_75t_L g701 ( .A(n_702), .B(n_706), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_705), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
INVx2_ASAP7_75t_L g733 ( .A(n_711), .Y(n_733) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g713 ( .A(n_714), .B(n_723), .Y(n_713) );
NOR2x1_ASAP7_75t_L g714 ( .A(n_715), .B(n_720), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NOR2x1_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
XNOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_745), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_749), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
INVx2_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_758), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_756), .B(n_759), .Y(n_796) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
OAI222xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_786), .B1(n_788), .B2(n_793), .C1(n_794), .C2(n_797), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NAND4xp25_ASAP7_75t_SL g769 ( .A(n_770), .B(n_774), .C(n_778), .D(n_783), .Y(n_769) );
AND4x1_ASAP7_75t_L g792 ( .A(n_770), .B(n_774), .C(n_778), .D(n_783), .Y(n_792) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_772), .Y(n_770) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_SL g794 ( .A(n_795), .Y(n_794) );
CKINVDCx6p67_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
endmodule