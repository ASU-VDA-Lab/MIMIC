module fake_jpeg_18673_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_20),
.Y(n_60)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_44),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx12f_ASAP7_75t_SL g45 ( 
.A(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_50),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_31),
.B1(n_24),
.B2(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_57),
.A2(n_61),
.B1(n_70),
.B2(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_62),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_31),
.B1(n_24),
.B2(n_23),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_20),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_31),
.B1(n_17),
.B2(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_19),
.B1(n_29),
.B2(n_18),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_23),
.B1(n_17),
.B2(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_74),
.Y(n_98)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_37),
.B(n_30),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_17),
.B1(n_48),
.B2(n_40),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_89),
.B(n_100),
.Y(n_129)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_85),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_51),
.C(n_20),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_56),
.C(n_55),
.Y(n_121)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_32),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_SL g135 ( 
.A1(n_80),
.A2(n_81),
.B(n_75),
.Y(n_135)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_62),
.B(n_20),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_103),
.Y(n_113)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_36),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_36),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_91),
.B1(n_95),
.B2(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_66),
.A2(n_32),
.B1(n_19),
.B2(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_88),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_21),
.B(n_25),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_90),
.B(n_97),
.Y(n_125)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_93),
.Y(n_133)
);

BUFx2_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_64),
.A2(n_29),
.B1(n_27),
.B2(n_35),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_20),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_105),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_28),
.B(n_25),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_29),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_27),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_18),
.B1(n_21),
.B2(n_33),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_68),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_33),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_109),
.B1(n_13),
.B2(n_4),
.Y(n_130)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_55),
.A2(n_33),
.B1(n_1),
.B2(n_2),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_111),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_0),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_135),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_122),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_58),
.C(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_124),
.B1(n_130),
.B2(n_102),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_134),
.A2(n_102),
.B1(n_81),
.B2(n_78),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_126),
.B(n_106),
.Y(n_167)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_87),
.B1(n_75),
.B2(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_117),
.B1(n_113),
.B2(n_126),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_98),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_145),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_77),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_146),
.Y(n_161)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_79),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_117),
.B(n_120),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_150),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_77),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_153),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_119),
.A2(n_83),
.B1(n_99),
.B2(n_75),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_152),
.A2(n_129),
.B1(n_122),
.B2(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_83),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_157),
.A2(n_140),
.B1(n_147),
.B2(n_148),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_136),
.B(n_121),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_159),
.B(n_174),
.Y(n_184)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_138),
.Y(n_187)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_143),
.A2(n_129),
.B(n_126),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_173),
.B(n_143),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_172),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_88),
.B(n_123),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_93),
.Y(n_174)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_175),
.Y(n_192)
);

OA21x2_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_179),
.B(n_183),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_177),
.B(n_186),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_182),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_153),
.C(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_139),
.A3(n_141),
.B1(n_152),
.B2(n_154),
.C1(n_148),
.C2(n_144),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_185),
.A2(n_189),
.B1(n_165),
.B2(n_164),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_160),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_169),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_133),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_159),
.B(n_105),
.C(n_132),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_190),
.B(n_174),
.C(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_131),
.Y(n_191)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_205),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_199),
.C(n_204),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_166),
.B(n_172),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_196),
.A2(n_176),
.B(n_187),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_197),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_167),
.C(n_169),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_184),
.B(n_171),
.C(n_158),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_171),
.C(n_166),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_173),
.C(n_92),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_213),
.B(n_214),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_188),
.B1(n_186),
.B2(n_180),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_196),
.B1(n_197),
.B2(n_203),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_182),
.B(n_161),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_193),
.A2(n_189),
.B1(n_170),
.B2(n_181),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_217),
.B1(n_101),
.B2(n_7),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_204),
.B(n_162),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_215),
.B(n_198),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_195),
.C(n_199),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_194),
.A2(n_107),
.B1(n_82),
.B2(n_76),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_224),
.C(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_221),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_198),
.C(n_132),
.Y(n_224)
);

OAI31xp33_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_133),
.A3(n_131),
.B(n_92),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_227),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_226),
.B(n_209),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_232),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_222),
.A2(n_211),
.B(n_208),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_231),
.A2(n_223),
.B(n_220),
.Y(n_234)
);

AOI31xp33_ASAP7_75t_L g233 ( 
.A1(n_225),
.A2(n_217),
.A3(n_216),
.B(n_218),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_233),
.A2(n_212),
.B(n_7),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_236),
.B(n_237),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_230),
.A2(n_227),
.B1(n_224),
.B2(n_219),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_229),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_108),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_238),
.A2(n_3),
.B1(n_9),
.B2(n_11),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_239),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_11),
.B(n_12),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_11),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_244),
.A2(n_245),
.B(n_13),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_13),
.Y(n_247)
);


endmodule