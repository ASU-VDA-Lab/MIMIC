module fake_netlist_6_4826_n_2871 (n_52, n_591, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_590, n_625, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_607, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_595, n_627, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_628, n_557, n_349, n_643, n_233, n_617, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_615, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_639, n_327, n_369, n_597, n_280, n_287, n_353, n_610, n_555, n_389, n_415, n_65, n_230, n_605, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_644, n_621, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_601, n_338, n_522, n_466, n_506, n_56, n_360, n_603, n_119, n_235, n_536, n_622, n_147, n_191, n_340, n_387, n_452, n_616, n_39, n_344, n_73, n_581, n_428, n_609, n_432, n_641, n_101, n_167, n_631, n_174, n_127, n_516, n_153, n_525, n_611, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_647, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_614, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_638, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_648, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_626, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_624, n_279, n_252, n_228, n_565, n_594, n_356, n_577, n_166, n_184, n_552, n_619, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_592, n_323, n_606, n_393, n_411, n_503, n_152, n_623, n_92, n_599, n_513, n_321, n_645, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_608, n_620, n_420, n_630, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_589, n_481, n_325, n_329, n_464, n_600, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_635, n_95, n_311, n_10, n_403, n_253, n_634, n_583, n_596, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_642, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_618, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_612, n_633, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_632, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_604, n_120, n_251, n_301, n_274, n_636, n_110, n_151, n_412, n_640, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_598, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_593, n_514, n_646, n_528, n_391, n_457, n_364, n_637, n_295, n_385, n_629, n_388, n_190, n_262, n_484, n_613, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_602, n_194, n_171, n_192, n_57, n_169, n_51, n_649, n_283, n_2871);

input n_52;
input n_591;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_590;
input n_625;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_607;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_595;
input n_627;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_628;
input n_557;
input n_349;
input n_643;
input n_233;
input n_617;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_615;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_639;
input n_327;
input n_369;
input n_597;
input n_280;
input n_287;
input n_353;
input n_610;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_605;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_644;
input n_621;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_601;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_603;
input n_119;
input n_235;
input n_536;
input n_622;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_616;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_609;
input n_432;
input n_641;
input n_101;
input n_167;
input n_631;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_611;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_647;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_614;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_638;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_648;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_626;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_624;
input n_279;
input n_252;
input n_228;
input n_565;
input n_594;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_619;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_592;
input n_323;
input n_606;
input n_393;
input n_411;
input n_503;
input n_152;
input n_623;
input n_92;
input n_599;
input n_513;
input n_321;
input n_645;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_608;
input n_620;
input n_420;
input n_630;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_589;
input n_481;
input n_325;
input n_329;
input n_464;
input n_600;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_635;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_634;
input n_583;
input n_596;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_642;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_618;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_612;
input n_633;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_632;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_604;
input n_120;
input n_251;
input n_301;
input n_274;
input n_636;
input n_110;
input n_151;
input n_412;
input n_640;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_598;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_593;
input n_514;
input n_646;
input n_528;
input n_391;
input n_457;
input n_364;
input n_637;
input n_295;
input n_385;
input n_629;
input n_388;
input n_190;
input n_262;
input n_484;
input n_613;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_602;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_649;
input n_283;

output n_2871;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_2405;
wire n_1743;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_2838;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2510;
wire n_1954;
wire n_1735;
wire n_2044;
wire n_1541;
wire n_1300;
wire n_2480;
wire n_2739;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_2786;
wire n_1591;
wire n_772;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_1094;
wire n_953;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2735;
wire n_1843;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_2778;
wire n_2850;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_2101;
wire n_2696;
wire n_2059;
wire n_2198;
wire n_2669;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_2692;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2654;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_2355;
wire n_966;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1950;
wire n_1726;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_2641;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2345;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_2347;
wire n_850;
wire n_690;
wire n_1886;
wire n_1801;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_2810;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_696;
wire n_1515;
wire n_961;
wire n_1317;
wire n_1082;
wire n_2733;
wire n_2824;
wire n_687;
wire n_697;
wire n_890;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_2644;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2728;
wire n_2349;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_2691;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_2436;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_1293;
wire n_2693;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_682;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_2590;
wire n_2643;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2650;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2718;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_683;
wire n_1207;
wire n_811;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_1250;
wire n_958;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2552;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_2724;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2502;
wire n_2131;
wire n_2226;
wire n_2801;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_2732;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2720;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_2289;
wire n_1419;
wire n_2863;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_2627;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_2756;
wire n_1871;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_2755;
wire n_923;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2819;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2401;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2716;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_2789;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_776;
wire n_1823;
wire n_2479;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1962;
wire n_1236;
wire n_1794;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_2671;
wire n_2761;
wire n_2793;
wire n_2715;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1929;
wire n_1807;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_823;
wire n_1132;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_2746;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_2736;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_1561;
wire n_2741;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_2743;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2466;
wire n_2111;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_2662;
wire n_753;
wire n_1753;
wire n_2795;
wire n_2471;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_2774;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2632;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_2659;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g650 ( 
.A(n_534),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_526),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_506),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_493),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

BUFx8_ASAP7_75t_SL g655 ( 
.A(n_161),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_377),
.Y(n_656)
);

CKINVDCx20_ASAP7_75t_R g657 ( 
.A(n_401),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_517),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_267),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_437),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_539),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_571),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_256),
.Y(n_663)
);

CKINVDCx14_ASAP7_75t_R g664 ( 
.A(n_147),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_585),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_360),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_80),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_448),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_220),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_633),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_292),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_95),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_524),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_7),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_186),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_456),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_611),
.Y(n_677)
);

BUFx10_ASAP7_75t_L g678 ( 
.A(n_601),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_504),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_565),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_193),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_302),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_605),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_135),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_167),
.Y(n_685)
);

CKINVDCx16_ASAP7_75t_R g686 ( 
.A(n_229),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_556),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_192),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_576),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_594),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_63),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_88),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_480),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_37),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_17),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_471),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_47),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_543),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_595),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_549),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_308),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_342),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_527),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_142),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_172),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_152),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_76),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_472),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_51),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_617),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_318),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_65),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_366),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_315),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_124),
.Y(n_716)
);

BUFx10_ASAP7_75t_L g717 ( 
.A(n_484),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_296),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_346),
.Y(n_719)
);

CKINVDCx20_ASAP7_75t_R g720 ( 
.A(n_148),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_68),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_612),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_528),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_511),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_496),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_649),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_542),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_466),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_155),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_316),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_162),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_154),
.Y(n_732)
);

BUFx10_ASAP7_75t_L g733 ( 
.A(n_513),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_505),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_403),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_215),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_638),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_613),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_364),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_259),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_130),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_553),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_14),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_431),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_149),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_327),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_623),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_320),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_271),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_530),
.Y(n_750)
);

CKINVDCx16_ASAP7_75t_R g751 ( 
.A(n_648),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_202),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_615),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_255),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_488),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_442),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_303),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_141),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_482),
.Y(n_759)
);

CKINVDCx14_ASAP7_75t_R g760 ( 
.A(n_592),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_7),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_521),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_296),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_516),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_218),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_246),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_199),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_415),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_259),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_522),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_1),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_107),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_430),
.Y(n_773)
);

CKINVDCx14_ASAP7_75t_R g774 ( 
.A(n_641),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_341),
.Y(n_775)
);

BUFx8_ASAP7_75t_SL g776 ( 
.A(n_290),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_2),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_264),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_137),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_523),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_369),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_108),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_610),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_111),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_349),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_145),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_344),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_278),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_277),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_310),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_432),
.Y(n_791)
);

BUFx10_ASAP7_75t_L g792 ( 
.A(n_642),
.Y(n_792)
);

BUFx10_ASAP7_75t_L g793 ( 
.A(n_236),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_101),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_163),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_128),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_478),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_559),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_647),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_105),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_152),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_269),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_591),
.Y(n_803)
);

INVx4_ASAP7_75t_R g804 ( 
.A(n_614),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_624),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_551),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_386),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_62),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_277),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_406),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_367),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_48),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_378),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_627),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_96),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_418),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_85),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_168),
.Y(n_818)
);

BUFx10_ASAP7_75t_L g819 ( 
.A(n_78),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_257),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_236),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_620),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_204),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_532),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_515),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_567),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_519),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_454),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_209),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_588),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_548),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_560),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_345),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_397),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_326),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_554),
.Y(n_836)
);

CKINVDCx20_ASAP7_75t_R g837 ( 
.A(n_604),
.Y(n_837)
);

BUFx10_ASAP7_75t_L g838 ( 
.A(n_596),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_439),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_70),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_597),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_577),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_644),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_90),
.Y(n_844)
);

BUFx10_ASAP7_75t_L g845 ( 
.A(n_570),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_60),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_335),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_271),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_68),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_356),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_168),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_166),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_139),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_322),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_192),
.Y(n_855)
);

CKINVDCx20_ASAP7_75t_R g856 ( 
.A(n_49),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_148),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_108),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_310),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_586),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_110),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_128),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_116),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_569),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_238),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_301),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_129),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_440),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_172),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_354),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_132),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_629),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_563),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_228),
.Y(n_874)
);

CKINVDCx20_ASAP7_75t_R g875 ( 
.A(n_35),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_154),
.Y(n_876)
);

CKINVDCx20_ASAP7_75t_R g877 ( 
.A(n_467),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_41),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_602),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_574),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_579),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_269),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_180),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_75),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_123),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_609),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_205),
.Y(n_887)
);

BUFx5_ASAP7_75t_L g888 ( 
.A(n_540),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_196),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_78),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_166),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_179),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_6),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_545),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_158),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_398),
.Y(n_896)
);

BUFx10_ASAP7_75t_L g897 ( 
.A(n_279),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_24),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_474),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_376),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_115),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_459),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_146),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_582),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_27),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_334),
.Y(n_906)
);

CKINVDCx14_ASAP7_75t_R g907 ( 
.A(n_636),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_414),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_443),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_94),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_309),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_137),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_392),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_120),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_51),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_48),
.Y(n_916)
);

CKINVDCx16_ASAP7_75t_R g917 ( 
.A(n_191),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_580),
.Y(n_918)
);

BUFx5_ASAP7_75t_L g919 ( 
.A(n_550),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_312),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_324),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_508),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_1),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_619),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_637),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_47),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_562),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_370),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_357),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_462),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_589),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_220),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_66),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_358),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_173),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_197),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_111),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_274),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_200),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_234),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_42),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_275),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_622),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_546),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_572),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_410),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_643),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_169),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_412),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_388),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_634),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_272),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_57),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_251),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_420),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_514),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_350),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_300),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_213),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_635),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_171),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_127),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_14),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_169),
.Y(n_964)
);

BUFx3_ASAP7_75t_L g965 ( 
.A(n_291),
.Y(n_965)
);

CKINVDCx20_ASAP7_75t_R g966 ( 
.A(n_461),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_290),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_6),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_92),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_9),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_458),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_162),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_628),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_184),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_244),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_409),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_411),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_257),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_198),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_541),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_221),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_72),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_600),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_237),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_330),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_566),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_329),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_37),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_339),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_351),
.Y(n_990)
);

CKINVDCx5p33_ASAP7_75t_R g991 ( 
.A(n_552),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_12),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_533),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_279),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_171),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_138),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_196),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_337),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_616),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_195),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_385),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_191),
.Y(n_1002)
);

CKINVDCx16_ASAP7_75t_R g1003 ( 
.A(n_507),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_238),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_391),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_413),
.Y(n_1006)
);

CKINVDCx14_ASAP7_75t_R g1007 ( 
.A(n_227),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_547),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_525),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_240),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_630),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_446),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_453),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_557),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_593),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_0),
.Y(n_1016)
);

BUFx5_ASAP7_75t_L g1017 ( 
.A(n_336),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_608),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_303),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_5),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_536),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_228),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_30),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_544),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_26),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_626),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_645),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_537),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_487),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_177),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_149),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_272),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_561),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_187),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_230),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_363),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_21),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_22),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_32),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_104),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_311),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_188),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_200),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_435),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_555),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_297),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_234),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_197),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_233),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_502),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_632),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_606),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_113),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_584),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_444),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_132),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_625),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_646),
.Y(n_1058)
);

INVx1_ASAP7_75t_SL g1059 ( 
.A(n_299),
.Y(n_1059)
);

BUFx10_ASAP7_75t_L g1060 ( 
.A(n_538),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_639),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_473),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_323),
.Y(n_1063)
);

CKINVDCx16_ASAP7_75t_R g1064 ( 
.A(n_394),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_590),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_255),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_45),
.Y(n_1067)
);

CKINVDCx20_ASAP7_75t_R g1068 ( 
.A(n_578),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_65),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_190),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_390),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_205),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_361),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_246),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_321),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_535),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_512),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_529),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_603),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_77),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_289),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_343),
.Y(n_1082)
);

CKINVDCx16_ASAP7_75t_R g1083 ( 
.A(n_423),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_18),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_309),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_518),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_501),
.Y(n_1087)
);

BUFx5_ASAP7_75t_L g1088 ( 
.A(n_92),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_510),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_227),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_500),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_621),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_449),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_164),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_598),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_73),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_25),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_304),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_581),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_232),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_464),
.Y(n_1101)
);

CKINVDCx20_ASAP7_75t_R g1102 ( 
.A(n_607),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_84),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_583),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_56),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_69),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_520),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_393),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_489),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_32),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_206),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_306),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_575),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_558),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_150),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_429),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_313),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_287),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_297),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_256),
.Y(n_1120)
);

CKINVDCx14_ASAP7_75t_R g1121 ( 
.A(n_587),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_338),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_631),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_531),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_298),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_305),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_86),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_568),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_331),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_174),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_509),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_207),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_265),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_229),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_564),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_16),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_13),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_193),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_136),
.Y(n_1139)
);

INVx1_ASAP7_75t_SL g1140 ( 
.A(n_248),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_307),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_188),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_179),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_599),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_640),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_295),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_573),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_42),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_198),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_490),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_100),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_239),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_L g1153 ( 
.A(n_752),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_681),
.Y(n_1154)
);

AND2x6_ASAP7_75t_L g1155 ( 
.A(n_670),
.B(n_314),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_928),
.B(n_0),
.Y(n_1156)
);

AND2x6_ASAP7_75t_L g1157 ( 
.A(n_670),
.B(n_317),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_693),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_670),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1088),
.Y(n_1160)
);

INVx4_ASAP7_75t_L g1161 ( 
.A(n_670),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_700),
.Y(n_1162)
);

CKINVDCx11_ASAP7_75t_R g1163 ( 
.A(n_793),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_664),
.B(n_2),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_681),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_664),
.B(n_3),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1007),
.B(n_3),
.Y(n_1167)
);

INVx5_ASAP7_75t_L g1168 ( 
.A(n_700),
.Y(n_1168)
);

INVx5_ASAP7_75t_L g1169 ( 
.A(n_700),
.Y(n_1169)
);

AND2x6_ASAP7_75t_L g1170 ( 
.A(n_700),
.B(n_319),
.Y(n_1170)
);

BUFx12f_ASAP7_75t_L g1171 ( 
.A(n_786),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_752),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_911),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1007),
.B(n_4),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1094),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_703),
.B(n_4),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_752),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1088),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_752),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_678),
.Y(n_1180)
);

BUFx12f_ASAP7_75t_L g1181 ( 
.A(n_786),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1088),
.B(n_5),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_879),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1088),
.Y(n_1184)
);

BUFx8_ASAP7_75t_SL g1185 ( 
.A(n_655),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1088),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_699),
.B(n_8),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1088),
.B(n_8),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1088),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_879),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_879),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_903),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_696),
.B(n_9),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_903),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_903),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_703),
.B(n_735),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_903),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_879),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_963),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_963),
.Y(n_1200)
);

BUFx8_ASAP7_75t_SL g1201 ( 
.A(n_776),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_735),
.B(n_10),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_902),
.Y(n_1203)
);

AND2x4_ASAP7_75t_L g1204 ( 
.A(n_834),
.B(n_10),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_805),
.B(n_11),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_696),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_843),
.B(n_11),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_850),
.B(n_12),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_963),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_891),
.B(n_13),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_834),
.B(n_945),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_902),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_899),
.B(n_15),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_686),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_718),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_891),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_SL g1217 ( 
.A(n_751),
.B(n_15),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_963),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_971),
.B(n_16),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1078),
.B(n_17),
.Y(n_1220)
);

INVx5_ASAP7_75t_L g1221 ( 
.A(n_902),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_651),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_652),
.B(n_18),
.Y(n_1223)
);

BUFx6f_ASAP7_75t_L g1224 ( 
.A(n_1046),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_652),
.B(n_19),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_902),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_654),
.B(n_19),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1046),
.Y(n_1228)
);

INVx5_ASAP7_75t_L g1229 ( 
.A(n_1107),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_945),
.B(n_20),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_654),
.B(n_20),
.Y(n_1231)
);

BUFx6f_ASAP7_75t_L g1232 ( 
.A(n_1046),
.Y(n_1232)
);

INVx5_ASAP7_75t_L g1233 ( 
.A(n_1107),
.Y(n_1233)
);

INVxp67_ASAP7_75t_L g1234 ( 
.A(n_802),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1046),
.Y(n_1235)
);

BUFx12f_ASAP7_75t_L g1236 ( 
.A(n_786),
.Y(n_1236)
);

NOR2x1_ASAP7_75t_L g1237 ( 
.A(n_980),
.B(n_325),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_781),
.B(n_21),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_867),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1003),
.B(n_1064),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_980),
.B(n_22),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1100),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1100),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_965),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1107),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1100),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1107),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_989),
.B(n_23),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_917),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_989),
.B(n_23),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_867),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_867),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1100),
.Y(n_1253)
);

NOR2x1_ASAP7_75t_L g1254 ( 
.A(n_1001),
.B(n_328),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1137),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1001),
.Y(n_1256)
);

AND2x6_ASAP7_75t_L g1257 ( 
.A(n_1018),
.B(n_332),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_SL g1258 ( 
.A(n_1083),
.B(n_24),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1137),
.Y(n_1259)
);

CKINVDCx11_ASAP7_75t_R g1260 ( 
.A(n_793),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_653),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_678),
.Y(n_1262)
);

INVx2_ASAP7_75t_L g1263 ( 
.A(n_1137),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1137),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_660),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_965),
.Y(n_1266)
);

AND2x6_ASAP7_75t_L g1267 ( 
.A(n_1018),
.B(n_333),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_733),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_781),
.B(n_25),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1111),
.B(n_26),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_717),
.Y(n_1271)
);

BUFx6f_ASAP7_75t_L g1272 ( 
.A(n_1111),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_650),
.B(n_27),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1132),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_810),
.B(n_28),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_810),
.B(n_28),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1132),
.Y(n_1277)
);

INVx5_ASAP7_75t_L g1278 ( 
.A(n_717),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_881),
.B(n_29),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_888),
.Y(n_1280)
);

BUFx8_ASAP7_75t_SL g1281 ( 
.A(n_713),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_881),
.B(n_29),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_944),
.B(n_30),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_944),
.B(n_31),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_946),
.B(n_31),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_865),
.Y(n_1286)
);

INVx5_ASAP7_75t_L g1287 ( 
.A(n_717),
.Y(n_1287)
);

INVx5_ASAP7_75t_L g1288 ( 
.A(n_792),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_733),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_946),
.B(n_33),
.Y(n_1290)
);

AND2x4_ASAP7_75t_L g1291 ( 
.A(n_656),
.B(n_33),
.Y(n_1291)
);

INVx5_ASAP7_75t_L g1292 ( 
.A(n_792),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_662),
.Y(n_1293)
);

BUFx6f_ASAP7_75t_L g1294 ( 
.A(n_1139),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1139),
.Y(n_1295)
);

AND2x4_ASAP7_75t_L g1296 ( 
.A(n_658),
.B(n_661),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_947),
.B(n_34),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_669),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1146),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_947),
.B(n_34),
.Y(n_1301)
);

INVxp33_ASAP7_75t_SL g1302 ( 
.A(n_948),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_845),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_976),
.B(n_35),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_669),
.Y(n_1305)
);

INVx4_ASAP7_75t_L g1306 ( 
.A(n_666),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_976),
.B(n_36),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_986),
.B(n_36),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_888),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_986),
.B(n_38),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1004),
.Y(n_1311)
);

INVx5_ASAP7_75t_L g1312 ( 
.A(n_792),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_672),
.B(n_38),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_672),
.B(n_39),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_663),
.Y(n_1315)
);

INVx3_ASAP7_75t_L g1316 ( 
.A(n_819),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_675),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_888),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_695),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1089),
.B(n_39),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_819),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1089),
.B(n_40),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_888),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_665),
.B(n_40),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_838),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1271),
.B(n_760),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1240),
.A2(n_774),
.B1(n_907),
.B2(n_760),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1271),
.B(n_1278),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1217),
.A2(n_853),
.B1(n_887),
.B2(n_745),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1153),
.Y(n_1330)
);

INVx2_ASAP7_75t_SL g1331 ( 
.A(n_1180),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1153),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1302),
.A2(n_907),
.B1(n_1121),
.B2(n_774),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1278),
.B(n_1121),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1281),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1167),
.A2(n_677),
.B1(n_690),
.B2(n_657),
.Y(n_1336)
);

INVxp33_ASAP7_75t_L g1337 ( 
.A(n_1214),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1287),
.B(n_845),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1258),
.A2(n_1059),
.B1(n_1140),
.B2(n_1042),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1192),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1166),
.A2(n_727),
.B1(n_799),
.B2(n_709),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1287),
.B(n_838),
.Y(n_1342)
);

AO22x2_ASAP7_75t_L g1343 ( 
.A1(n_1156),
.A2(n_702),
.B1(n_893),
.B2(n_674),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1288),
.B(n_838),
.Y(n_1344)
);

OAI22xp33_ASAP7_75t_SL g1345 ( 
.A1(n_1164),
.A2(n_667),
.B1(n_671),
.B2(n_659),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1215),
.B(n_1141),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1262),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1166),
.A2(n_837),
.B1(n_847),
.B2(n_803),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1306),
.B(n_704),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1174),
.A2(n_886),
.B1(n_950),
.B2(n_877),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1172),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1195),
.Y(n_1352)
);

AO22x2_ASAP7_75t_L g1353 ( 
.A1(n_1174),
.A2(n_767),
.B1(n_769),
.B2(n_695),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1249),
.A2(n_688),
.B1(n_692),
.B2(n_685),
.Y(n_1354)
);

AO22x2_ASAP7_75t_L g1355 ( 
.A1(n_1176),
.A2(n_769),
.B1(n_784),
.B2(n_767),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1234),
.A2(n_1068),
.B1(n_1101),
.B2(n_966),
.Y(n_1356)
);

OA22x2_ASAP7_75t_L g1357 ( 
.A1(n_1286),
.A2(n_684),
.B1(n_698),
.B2(n_682),
.Y(n_1357)
);

OA22x2_ASAP7_75t_L g1358 ( 
.A1(n_1311),
.A2(n_1158),
.B1(n_1175),
.B2(n_1173),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1158),
.A2(n_794),
.B1(n_808),
.B2(n_720),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1172),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1197),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1173),
.A2(n_1117),
.B1(n_1102),
.B2(n_706),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1175),
.A2(n_710),
.B1(n_716),
.B2(n_705),
.Y(n_1363)
);

AOI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1187),
.A2(n_1205),
.B1(n_1171),
.B2(n_1181),
.Y(n_1364)
);

BUFx16f_ASAP7_75t_R g1365 ( 
.A(n_1202),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1177),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1272),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1199),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1200),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1236),
.A2(n_1239),
.B1(n_1252),
.B2(n_1251),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1222),
.B(n_1093),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1207),
.A2(n_731),
.B1(n_732),
.B2(n_729),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1208),
.A2(n_743),
.B1(n_749),
.B2(n_740),
.Y(n_1373)
);

AO22x2_ASAP7_75t_L g1374 ( 
.A1(n_1204),
.A2(n_789),
.B1(n_920),
.B2(n_784),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_SL g1375 ( 
.A1(n_1268),
.A2(n_875),
.B1(n_912),
.B2(n_856),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1242),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1261),
.B(n_1093),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1177),
.Y(n_1378)
);

AOI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1321),
.A2(n_757),
.B1(n_758),
.B2(n_754),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1288),
.B(n_1060),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1289),
.B(n_841),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1316),
.A2(n_765),
.B1(n_766),
.B2(n_761),
.Y(n_1382)
);

OA22x2_ASAP7_75t_L g1383 ( 
.A1(n_1244),
.A2(n_708),
.B1(n_721),
.B2(n_707),
.Y(n_1383)
);

OAI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1213),
.A2(n_1220),
.B1(n_1219),
.B2(n_1188),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1292),
.B(n_1060),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1303),
.B(n_789),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1182),
.A2(n_778),
.B1(n_779),
.B2(n_771),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1292),
.B(n_1060),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1265),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1312),
.B(n_897),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1312),
.B(n_897),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_SL g1392 ( 
.A(n_1325),
.B(n_782),
.Y(n_1392)
);

AO22x2_ASAP7_75t_L g1393 ( 
.A1(n_1230),
.A2(n_942),
.B1(n_1090),
.B2(n_920),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1325),
.A2(n_1225),
.B1(n_1231),
.B2(n_1223),
.Y(n_1394)
);

OAI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1269),
.A2(n_796),
.B1(n_800),
.B2(n_788),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1293),
.A2(n_809),
.B1(n_812),
.B2(n_801),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1185),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1244),
.B(n_676),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1241),
.A2(n_817),
.B1(n_821),
.B2(n_815),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1274),
.B(n_683),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1274),
.B(n_687),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1196),
.B(n_691),
.Y(n_1402)
);

AOI22x1_ASAP7_75t_L g1403 ( 
.A1(n_1193),
.A2(n_1210),
.B1(n_1270),
.B2(n_1313),
.Y(n_1403)
);

OAI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1276),
.A2(n_829),
.B1(n_846),
.B2(n_823),
.Y(n_1404)
);

OAI22xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1284),
.A2(n_1308),
.B1(n_1320),
.B2(n_1285),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1248),
.A2(n_849),
.B1(n_851),
.B2(n_848),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1250),
.A2(n_1227),
.B1(n_1275),
.B2(n_1238),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1279),
.A2(n_855),
.B1(n_857),
.B2(n_852),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1211),
.B(n_694),
.Y(n_1409)
);

AO22x2_ASAP7_75t_L g1410 ( 
.A1(n_1193),
.A2(n_1270),
.B1(n_1210),
.B2(n_1090),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1256),
.B(n_668),
.Y(n_1411)
);

OR2x2_ASAP7_75t_L g1412 ( 
.A(n_1154),
.B(n_858),
.Y(n_1412)
);

OAI22xp33_ASAP7_75t_R g1413 ( 
.A1(n_1315),
.A2(n_741),
.B1(n_763),
.B2(n_736),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1322),
.A2(n_862),
.B1(n_866),
.B2(n_861),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1282),
.A2(n_874),
.B1(n_878),
.B2(n_871),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1255),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1283),
.A2(n_884),
.B1(n_885),
.B2(n_883),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1165),
.B(n_697),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1179),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1272),
.B(n_1277),
.Y(n_1420)
);

AND2x2_ASAP7_75t_SL g1421 ( 
.A(n_1313),
.B(n_942),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1259),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1290),
.A2(n_892),
.B1(n_895),
.B2(n_890),
.Y(n_1423)
);

AND2x4_ASAP7_75t_SL g1424 ( 
.A(n_1296),
.B(n_940),
.Y(n_1424)
);

OAI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1206),
.A2(n_901),
.B1(n_905),
.B2(n_898),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1297),
.A2(n_914),
.B1(n_915),
.B2(n_910),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1216),
.B(n_711),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1301),
.A2(n_926),
.B1(n_935),
.B2(n_916),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1304),
.A2(n_936),
.B1(n_961),
.B2(n_938),
.Y(n_1429)
);

AO22x2_ASAP7_75t_L g1430 ( 
.A1(n_1314),
.A2(n_777),
.B1(n_790),
.B2(n_772),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1277),
.B(n_795),
.Y(n_1431)
);

AOI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1307),
.A2(n_967),
.B1(n_968),
.B2(n_962),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_974),
.B2(n_970),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1273),
.A2(n_978),
.B1(n_979),
.B2(n_975),
.Y(n_1434)
);

OAI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1294),
.A2(n_992),
.B1(n_994),
.B2(n_984),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1201),
.Y(n_1436)
);

NAND2xp33_ASAP7_75t_SL g1437 ( 
.A(n_1314),
.B(n_953),
.Y(n_1437)
);

AO22x2_ASAP7_75t_L g1438 ( 
.A1(n_1291),
.A2(n_820),
.B1(n_840),
.B2(n_818),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1263),
.Y(n_1439)
);

AOI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1257),
.A2(n_996),
.B1(n_997),
.B2(n_995),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1179),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1257),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1257),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1294),
.Y(n_1444)
);

AO22x2_ASAP7_75t_L g1445 ( 
.A1(n_1324),
.A2(n_859),
.B1(n_863),
.B2(n_844),
.Y(n_1445)
);

OA22x2_ASAP7_75t_L g1446 ( 
.A1(n_1266),
.A2(n_876),
.B1(n_882),
.B2(n_869),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1295),
.Y(n_1447)
);

AO22x2_ASAP7_75t_L g1448 ( 
.A1(n_1300),
.A2(n_923),
.B1(n_932),
.B2(n_889),
.Y(n_1448)
);

OAI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1295),
.A2(n_1010),
.B1(n_1016),
.B2(n_1000),
.Y(n_1449)
);

OR2x2_ASAP7_75t_L g1450 ( 
.A(n_1298),
.B(n_1019),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1159),
.B(n_714),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1218),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1218),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1267),
.A2(n_1163),
.B1(n_1260),
.B2(n_1022),
.Y(n_1454)
);

AO22x2_ASAP7_75t_L g1455 ( 
.A1(n_1317),
.A2(n_937),
.B1(n_939),
.B2(n_933),
.Y(n_1455)
);

INVx3_ASAP7_75t_L g1456 ( 
.A(n_1224),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1224),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1228),
.Y(n_1458)
);

INVx1_ASAP7_75t_SL g1459 ( 
.A(n_1305),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1228),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1305),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1232),
.Y(n_1462)
);

AOI22x1_ASAP7_75t_L g1463 ( 
.A1(n_1299),
.A2(n_952),
.B1(n_954),
.B2(n_941),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1232),
.Y(n_1464)
);

AO22x2_ASAP7_75t_L g1465 ( 
.A1(n_1299),
.A2(n_964),
.B1(n_981),
.B2(n_958),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1243),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1267),
.A2(n_1023),
.B1(n_1030),
.B2(n_1020),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1243),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1246),
.Y(n_1469)
);

AOI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1267),
.A2(n_1035),
.B1(n_1037),
.B2(n_1032),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1246),
.Y(n_1471)
);

AND2x2_ASAP7_75t_SL g1472 ( 
.A(n_1161),
.B(n_673),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1253),
.Y(n_1473)
);

INVx3_ASAP7_75t_L g1474 ( 
.A(n_1253),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1159),
.B(n_715),
.Y(n_1475)
);

AO22x2_ASAP7_75t_L g1476 ( 
.A1(n_1319),
.A2(n_988),
.B1(n_1002),
.B2(n_982),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1168),
.B(n_722),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1264),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1237),
.A2(n_1040),
.B1(n_1043),
.B2(n_1039),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1319),
.B(n_1031),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1194),
.B(n_679),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1168),
.B(n_723),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1264),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1254),
.A2(n_1053),
.B1(n_1072),
.B2(n_1047),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1194),
.Y(n_1485)
);

NAND3x1_ASAP7_75t_L g1486 ( 
.A(n_1209),
.B(n_1038),
.C(n_1034),
.Y(n_1486)
);

AO22x2_ASAP7_75t_L g1487 ( 
.A1(n_1209),
.A2(n_1048),
.B1(n_1049),
.B2(n_1041),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1162),
.B(n_680),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1235),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1169),
.B(n_1074),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1235),
.Y(n_1491)
);

AO22x2_ASAP7_75t_L g1492 ( 
.A1(n_1189),
.A2(n_1067),
.B1(n_1069),
.B2(n_1056),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_R g1493 ( 
.A1(n_1280),
.A2(n_1085),
.B1(n_1112),
.B2(n_1098),
.Y(n_1493)
);

AO22x2_ASAP7_75t_L g1494 ( 
.A1(n_1189),
.A2(n_1115),
.B1(n_1118),
.B2(n_1070),
.Y(n_1494)
);

AO22x2_ASAP7_75t_L g1495 ( 
.A1(n_1309),
.A2(n_1130),
.B1(n_1138),
.B2(n_1126),
.Y(n_1495)
);

AO22x2_ASAP7_75t_L g1496 ( 
.A1(n_1318),
.A2(n_1151),
.B1(n_701),
.B2(n_712),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1169),
.B(n_724),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1160),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1155),
.A2(n_1081),
.B1(n_1084),
.B2(n_1080),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1178),
.A2(n_1097),
.B1(n_1103),
.B2(n_1096),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1323),
.A2(n_1119),
.B1(n_1125),
.B2(n_1110),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1190),
.B(n_725),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1190),
.B(n_726),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1184),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1186),
.A2(n_1133),
.B1(n_1134),
.B2(n_1127),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1183),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1155),
.A2(n_1142),
.B1(n_1143),
.B2(n_1136),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1155),
.A2(n_1149),
.B1(n_1152),
.B2(n_1148),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1191),
.B(n_689),
.Y(n_1509)
);

AO22x2_ASAP7_75t_L g1510 ( 
.A1(n_1203),
.A2(n_739),
.B1(n_742),
.B2(n_719),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1191),
.B(n_728),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1198),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1198),
.B(n_747),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1212),
.B(n_730),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1212),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1157),
.A2(n_969),
.B1(n_1025),
.B2(n_959),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1221),
.B(n_734),
.Y(n_1517)
);

OA22x2_ASAP7_75t_L g1518 ( 
.A1(n_1157),
.A2(n_756),
.B1(n_764),
.B2(n_748),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1221),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1226),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1226),
.B(n_737),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1229),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1229),
.A2(n_791),
.B1(n_814),
.B2(n_770),
.Y(n_1523)
);

AO22x2_ASAP7_75t_L g1524 ( 
.A1(n_1157),
.A2(n_816),
.B1(n_825),
.B2(n_822),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1233),
.B(n_738),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1233),
.B(n_744),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1247),
.B(n_746),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1247),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1170),
.A2(n_1105),
.B1(n_1106),
.B2(n_1066),
.Y(n_1529)
);

AND2x2_ASAP7_75t_SL g1530 ( 
.A(n_1170),
.B(n_826),
.Y(n_1530)
);

NOR2xp33_ASAP7_75t_L g1531 ( 
.A(n_1245),
.B(n_830),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1245),
.B(n_832),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1170),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_753),
.B2(n_755),
.Y(n_1534)
);

AOI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1240),
.A2(n_759),
.B1(n_762),
.B2(n_750),
.Y(n_1535)
);

INVx2_ASAP7_75t_SL g1536 ( 
.A(n_1180),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1271),
.B(n_768),
.Y(n_1537)
);

OAI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1217),
.A2(n_1028),
.B1(n_1065),
.B2(n_833),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1153),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1192),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1281),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1153),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1321),
.B(n_854),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1222),
.B(n_873),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1306),
.B(n_896),
.Y(n_1545)
);

AO22x2_ASAP7_75t_L g1546 ( 
.A1(n_1156),
.A2(n_904),
.B1(n_908),
.B2(n_906),
.Y(n_1546)
);

AO22x2_ASAP7_75t_L g1547 ( 
.A1(n_1156),
.A2(n_909),
.B1(n_925),
.B2(n_918),
.Y(n_1547)
);

AOI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1240),
.A2(n_775),
.B1(n_780),
.B2(n_773),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1192),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1271),
.B(n_783),
.Y(n_1550)
);

AND2x4_ASAP7_75t_L g1551 ( 
.A(n_1306),
.B(n_949),
.Y(n_1551)
);

AOI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1240),
.A2(n_787),
.B1(n_797),
.B2(n_785),
.Y(n_1552)
);

AOI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1240),
.A2(n_806),
.B1(n_807),
.B2(n_798),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_R g1554 ( 
.A1(n_1214),
.A2(n_983),
.B1(n_987),
.B2(n_977),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1217),
.A2(n_993),
.B1(n_1015),
.B2(n_990),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1240),
.A2(n_811),
.B1(n_824),
.B2(n_813),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1153),
.Y(n_1557)
);

OAI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1217),
.A2(n_1026),
.B1(n_1029),
.B2(n_1021),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1214),
.B(n_41),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1271),
.B(n_827),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1222),
.B(n_1044),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1217),
.A2(n_1061),
.B1(n_1062),
.B2(n_1050),
.Y(n_1562)
);

OAI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1217),
.A2(n_1075),
.B1(n_1079),
.B2(n_1071),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1222),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1240),
.A2(n_828),
.B1(n_835),
.B2(n_831),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1240),
.A2(n_836),
.B1(n_842),
.B2(n_839),
.Y(n_1566)
);

OAI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1217),
.A2(n_1091),
.B1(n_1108),
.B2(n_1082),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1240),
.A2(n_860),
.B1(n_868),
.B2(n_864),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1217),
.A2(n_1122),
.B1(n_1147),
.B2(n_1116),
.Y(n_1569)
);

AO22x2_ASAP7_75t_L g1570 ( 
.A1(n_1156),
.A2(n_804),
.B1(n_45),
.B2(n_43),
.Y(n_1570)
);

OA22x2_ASAP7_75t_L g1571 ( 
.A1(n_1234),
.A2(n_872),
.B1(n_880),
.B2(n_870),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1217),
.A2(n_900),
.B1(n_913),
.B2(n_894),
.Y(n_1572)
);

OAI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1217),
.A2(n_922),
.B1(n_924),
.B2(n_921),
.Y(n_1573)
);

OAI22xp33_ASAP7_75t_SL g1574 ( 
.A1(n_1217),
.A2(n_929),
.B1(n_930),
.B2(n_927),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1271),
.B(n_931),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1153),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1240),
.A2(n_943),
.B1(n_951),
.B2(n_934),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1217),
.A2(n_956),
.B1(n_957),
.B2(n_955),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1302),
.A2(n_973),
.B1(n_985),
.B2(n_960),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1217),
.A2(n_998),
.B1(n_999),
.B2(n_991),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1240),
.A2(n_1006),
.B1(n_1008),
.B2(n_1005),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1272),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1222),
.B(n_1009),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1222),
.B(n_1150),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1240),
.A2(n_1012),
.B1(n_1013),
.B2(n_1011),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1271),
.B(n_1014),
.Y(n_1586)
);

AO22x2_ASAP7_75t_L g1587 ( 
.A1(n_1156),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1153),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1271),
.B(n_1024),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1271),
.B(n_1027),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1153),
.Y(n_1591)
);

NAND3x1_ASAP7_75t_L g1592 ( 
.A(n_1164),
.B(n_44),
.C(n_46),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1302),
.A2(n_1036),
.B1(n_1045),
.B2(n_1033),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1240),
.A2(n_1052),
.B1(n_1054),
.B2(n_1051),
.Y(n_1594)
);

OAI22xp33_ASAP7_75t_L g1595 ( 
.A1(n_1217),
.A2(n_1057),
.B1(n_1058),
.B2(n_1055),
.Y(n_1595)
);

AOI22xp5_ASAP7_75t_SL g1596 ( 
.A1(n_1302),
.A2(n_1073),
.B1(n_1076),
.B2(n_1063),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1240),
.A2(n_1086),
.B1(n_1087),
.B2(n_1077),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1302),
.A2(n_1095),
.B1(n_1099),
.B2(n_1092),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_L g1599 ( 
.A1(n_1240),
.A2(n_1109),
.B1(n_1113),
.B2(n_1104),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1192),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1302),
.A2(n_1123),
.B1(n_1124),
.B2(n_1114),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1153),
.Y(n_1602)
);

OAI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1217),
.A2(n_1129),
.B1(n_1131),
.B2(n_1128),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1192),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1192),
.Y(n_1605)
);

OAI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1217),
.A2(n_1144),
.B1(n_1145),
.B2(n_1135),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1222),
.B(n_888),
.Y(n_1607)
);

OAI22xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1217),
.A2(n_919),
.B1(n_1017),
.B2(n_888),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1240),
.A2(n_1017),
.B1(n_919),
.B2(n_888),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1217),
.A2(n_1017),
.B1(n_919),
.B2(n_52),
.Y(n_1610)
);

AO22x2_ASAP7_75t_L g1611 ( 
.A1(n_1156),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_R g1612 ( 
.A1(n_1214),
.A2(n_54),
.B1(n_50),
.B2(n_53),
.Y(n_1612)
);

AO22x2_ASAP7_75t_L g1613 ( 
.A1(n_1156),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1192),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1192),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1271),
.B(n_1017),
.Y(n_1616)
);

OA22x2_ASAP7_75t_L g1617 ( 
.A1(n_1234),
.A2(n_1017),
.B1(n_919),
.B2(n_57),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1240),
.A2(n_1017),
.B1(n_919),
.B2(n_58),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1302),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1153),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1192),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1222),
.B(n_919),
.Y(n_1622)
);

AOI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1240),
.A2(n_1017),
.B1(n_919),
.B2(n_61),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_SL g1624 ( 
.A(n_1180),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1222),
.B(n_340),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1271),
.B(n_347),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1302),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1271),
.B(n_348),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1153),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1166),
.B(n_59),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1192),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1302),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1153),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1222),
.B(n_64),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1240),
.A2(n_69),
.B1(n_66),
.B2(n_67),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1192),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1153),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1240),
.A2(n_71),
.B1(n_67),
.B2(n_70),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1272),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1153),
.Y(n_1640)
);

OAI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1217),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1240),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1271),
.B(n_352),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1153),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1271),
.B(n_353),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1271),
.B(n_355),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1192),
.Y(n_1647)
);

AOI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1240),
.A2(n_79),
.B1(n_74),
.B2(n_77),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1306),
.B(n_359),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1302),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_SL g1651 ( 
.A(n_1180),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1321),
.B(n_81),
.Y(n_1652)
);

AO22x2_ASAP7_75t_L g1653 ( 
.A1(n_1156),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1653)
);

AO22x2_ASAP7_75t_L g1654 ( 
.A1(n_1156),
.A2(n_85),
.B1(n_82),
.B2(n_83),
.Y(n_1654)
);

AO22x2_ASAP7_75t_L g1655 ( 
.A1(n_1156),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1217),
.A2(n_90),
.B1(n_87),
.B2(n_89),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1271),
.B(n_362),
.Y(n_1657)
);

AND2x2_ASAP7_75t_SL g1658 ( 
.A(n_1217),
.B(n_89),
.Y(n_1658)
);

AOI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1240),
.A2(n_94),
.B1(n_91),
.B2(n_93),
.Y(n_1659)
);

OAI22xp33_ASAP7_75t_SL g1660 ( 
.A1(n_1217),
.A2(n_95),
.B1(n_91),
.B2(n_93),
.Y(n_1660)
);

OAI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1217),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1504),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1663)
);

BUFx6f_ASAP7_75t_L g1664 ( 
.A(n_1378),
.Y(n_1664)
);

NOR2xp67_ASAP7_75t_L g1665 ( 
.A(n_1564),
.B(n_365),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1498),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1544),
.B(n_97),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1340),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1352),
.Y(n_1669)
);

INVxp33_ASAP7_75t_SL g1670 ( 
.A(n_1579),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1361),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1368),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1398),
.B(n_98),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1459),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1522),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1461),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1441),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1369),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1452),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1457),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1376),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1466),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1473),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1483),
.Y(n_1684)
);

CKINVDCx16_ASAP7_75t_R g1685 ( 
.A(n_1341),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1330),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1472),
.B(n_368),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1561),
.B(n_99),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1346),
.B(n_99),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1607),
.B(n_371),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1622),
.B(n_1421),
.Y(n_1691)
);

AND2x2_ASAP7_75t_SL g1692 ( 
.A(n_1658),
.B(n_100),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1416),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1422),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1371),
.B(n_101),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1400),
.B(n_1401),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1332),
.Y(n_1697)
);

CKINVDCx20_ASAP7_75t_R g1698 ( 
.A(n_1389),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1351),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1360),
.Y(n_1700)
);

CKINVDCx20_ASAP7_75t_R g1701 ( 
.A(n_1348),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1366),
.Y(n_1702)
);

XNOR2xp5_ASAP7_75t_L g1703 ( 
.A(n_1336),
.B(n_102),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1338),
.B(n_102),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1519),
.Y(n_1705)
);

BUFx6f_ASAP7_75t_L g1706 ( 
.A(n_1378),
.Y(n_1706)
);

XOR2xp5_ASAP7_75t_L g1707 ( 
.A(n_1356),
.B(n_372),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1342),
.B(n_103),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1377),
.B(n_103),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1419),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1453),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1458),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1380),
.B(n_104),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1460),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1462),
.Y(n_1715)
);

INVxp33_ASAP7_75t_L g1716 ( 
.A(n_1337),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1539),
.Y(n_1717)
);

XOR2xp5_ASAP7_75t_L g1718 ( 
.A(n_1350),
.B(n_373),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1437),
.Y(n_1719)
);

CKINVDCx16_ASAP7_75t_R g1720 ( 
.A(n_1327),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1464),
.Y(n_1721)
);

NOR2xp67_ASAP7_75t_L g1722 ( 
.A(n_1583),
.B(n_374),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1469),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1471),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1584),
.B(n_105),
.Y(n_1725)
);

CKINVDCx16_ASAP7_75t_R g1726 ( 
.A(n_1516),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1478),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1539),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1542),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1557),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1335),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1576),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1588),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1591),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1602),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1572),
.B(n_106),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1620),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1381),
.B(n_106),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1402),
.B(n_375),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1385),
.B(n_107),
.Y(n_1740)
);

INVxp33_ASAP7_75t_L g1741 ( 
.A(n_1375),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1629),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1451),
.B(n_379),
.Y(n_1743)
);

INVxp67_ASAP7_75t_SL g1744 ( 
.A(n_1520),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1412),
.B(n_109),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1388),
.B(n_109),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1633),
.Y(n_1747)
);

XNOR2xp5_ASAP7_75t_L g1748 ( 
.A(n_1529),
.B(n_110),
.Y(n_1748)
);

XOR2xp5_ASAP7_75t_L g1749 ( 
.A(n_1541),
.B(n_1397),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1637),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1640),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1439),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1540),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1644),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1549),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1600),
.Y(n_1756)
);

BUFx6f_ASAP7_75t_L g1757 ( 
.A(n_1644),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1329),
.B(n_112),
.Y(n_1758)
);

CKINVDCx16_ASAP7_75t_R g1759 ( 
.A(n_1333),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1436),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1418),
.B(n_112),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1604),
.Y(n_1762)
);

INVxp33_ASAP7_75t_L g1763 ( 
.A(n_1359),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1578),
.B(n_113),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1580),
.B(n_114),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1605),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1614),
.Y(n_1767)
);

CKINVDCx16_ASAP7_75t_R g1768 ( 
.A(n_1362),
.Y(n_1768)
);

XNOR2x2_ASAP7_75t_L g1769 ( 
.A(n_1587),
.B(n_114),
.Y(n_1769)
);

XNOR2xp5_ASAP7_75t_L g1770 ( 
.A(n_1570),
.B(n_115),
.Y(n_1770)
);

INVxp33_ASAP7_75t_L g1771 ( 
.A(n_1363),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1615),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1624),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1595),
.B(n_116),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1621),
.Y(n_1775)
);

NOR2xp33_ASAP7_75t_L g1776 ( 
.A(n_1603),
.B(n_117),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1606),
.B(n_117),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1475),
.B(n_1477),
.Y(n_1778)
);

INVx8_ASAP7_75t_L g1779 ( 
.A(n_1543),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1631),
.Y(n_1780)
);

XNOR2x2_ASAP7_75t_L g1781 ( 
.A(n_1587),
.B(n_118),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1636),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1647),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1538),
.B(n_118),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1485),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1456),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1651),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1427),
.B(n_119),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1468),
.Y(n_1789)
);

XOR2xp5_ASAP7_75t_L g1790 ( 
.A(n_1370),
.B(n_1358),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1409),
.B(n_380),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1474),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1489),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1367),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1444),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1482),
.B(n_381),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1450),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_L g1798 ( 
.A(n_1555),
.B(n_1558),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1506),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1534),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1405),
.A2(n_383),
.B(n_382),
.Y(n_1801)
);

XOR2xp5_ASAP7_75t_L g1802 ( 
.A(n_1596),
.B(n_384),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1562),
.B(n_119),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1447),
.Y(n_1804)
);

INVx2_ASAP7_75t_SL g1805 ( 
.A(n_1424),
.Y(n_1805)
);

INVx2_ASAP7_75t_SL g1806 ( 
.A(n_1537),
.Y(n_1806)
);

CKINVDCx20_ASAP7_75t_R g1807 ( 
.A(n_1454),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1491),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1582),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1639),
.Y(n_1810)
);

XNOR2x2_ASAP7_75t_L g1811 ( 
.A(n_1611),
.B(n_120),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1535),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1481),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1420),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1420),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1495),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1495),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1331),
.B(n_121),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1446),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1431),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1431),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1496),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1496),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1601),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1480),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1480),
.Y(n_1826)
);

NOR2xp33_ASAP7_75t_L g1827 ( 
.A(n_1563),
.B(n_121),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1509),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1513),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1347),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1355),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1355),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1536),
.B(n_122),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1374),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1497),
.B(n_387),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1374),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1393),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1386),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1393),
.Y(n_1839)
);

OAI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1533),
.A2(n_395),
.B(n_389),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1512),
.Y(n_1841)
);

CKINVDCx16_ASAP7_75t_R g1842 ( 
.A(n_1593),
.Y(n_1842)
);

XOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1571),
.B(n_396),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1326),
.B(n_122),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1530),
.Y(n_1845)
);

INVxp33_ASAP7_75t_L g1846 ( 
.A(n_1426),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1353),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1353),
.Y(n_1848)
);

INVxp33_ASAP7_75t_L g1849 ( 
.A(n_1433),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1411),
.Y(n_1850)
);

XOR2xp5_ASAP7_75t_L g1851 ( 
.A(n_1548),
.B(n_399),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1386),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1334),
.B(n_123),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1515),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1463),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1455),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1518),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1455),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1410),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1434),
.B(n_124),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1410),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1448),
.Y(n_1862)
);

INVxp67_ASAP7_75t_SL g1863 ( 
.A(n_1616),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1567),
.B(n_125),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1403),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1448),
.Y(n_1866)
);

XOR2xp5_ASAP7_75t_L g1867 ( 
.A(n_1552),
.B(n_400),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1383),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1357),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1492),
.Y(n_1870)
);

XNOR2x1_ASAP7_75t_L g1871 ( 
.A(n_1611),
.B(n_1613),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1492),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1494),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1569),
.B(n_125),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1494),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1488),
.Y(n_1876)
);

CKINVDCx20_ASAP7_75t_R g1877 ( 
.A(n_1553),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1465),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1556),
.B(n_126),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1465),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1565),
.B(n_126),
.Y(n_1881)
);

AND2x4_ASAP7_75t_L g1882 ( 
.A(n_1609),
.B(n_402),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1476),
.Y(n_1883)
);

INVx4_ASAP7_75t_L g1884 ( 
.A(n_1649),
.Y(n_1884)
);

NOR2xp33_ASAP7_75t_L g1885 ( 
.A(n_1566),
.B(n_127),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1476),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1487),
.Y(n_1887)
);

NOR2xp33_ASAP7_75t_L g1888 ( 
.A(n_1568),
.B(n_129),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_L g1889 ( 
.A(n_1502),
.B(n_404),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1577),
.B(n_130),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1487),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1559),
.B(n_131),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1503),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1511),
.Y(n_1894)
);

XOR2x2_ASAP7_75t_L g1895 ( 
.A(n_1364),
.B(n_131),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_L g1896 ( 
.A(n_1581),
.B(n_133),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1585),
.Y(n_1897)
);

CKINVDCx20_ASAP7_75t_R g1898 ( 
.A(n_1594),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1514),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1517),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1521),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1550),
.B(n_133),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1525),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1526),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1527),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1531),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1532),
.Y(n_1907)
);

XOR2x2_ASAP7_75t_L g1908 ( 
.A(n_1379),
.B(n_134),
.Y(n_1908)
);

OR2x6_ASAP7_75t_L g1909 ( 
.A(n_1652),
.B(n_134),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1528),
.Y(n_1910)
);

CKINVDCx5p33_ASAP7_75t_R g1911 ( 
.A(n_1598),
.Y(n_1911)
);

CKINVDCx20_ASAP7_75t_R g1912 ( 
.A(n_1597),
.Y(n_1912)
);

XOR2xp5_ASAP7_75t_L g1913 ( 
.A(n_1599),
.B(n_405),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1573),
.B(n_1574),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1438),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1407),
.B(n_407),
.Y(n_1916)
);

OR2x6_ASAP7_75t_L g1917 ( 
.A(n_1652),
.B(n_135),
.Y(n_1917)
);

INVx2_ASAP7_75t_SL g1918 ( 
.A(n_1560),
.Y(n_1918)
);

NOR2xp33_ASAP7_75t_L g1919 ( 
.A(n_1396),
.B(n_136),
.Y(n_1919)
);

NOR2xp33_ASAP7_75t_L g1920 ( 
.A(n_1349),
.B(n_138),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1384),
.B(n_139),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_SL g1922 ( 
.A(n_1339),
.B(n_140),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1438),
.Y(n_1923)
);

INVxp33_ASAP7_75t_L g1924 ( 
.A(n_1408),
.Y(n_1924)
);

INVx2_ASAP7_75t_SL g1925 ( 
.A(n_1575),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1445),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1445),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1586),
.B(n_408),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1589),
.B(n_140),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1430),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_L g1931 ( 
.A(n_1590),
.B(n_416),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1429),
.B(n_141),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1399),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1430),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1617),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1545),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1354),
.B(n_142),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1551),
.Y(n_1938)
);

XOR2xp5_ASAP7_75t_L g1939 ( 
.A(n_1345),
.B(n_417),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1415),
.B(n_143),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1618),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1623),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1546),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1486),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1417),
.B(n_1423),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1546),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1547),
.Y(n_1947)
);

CKINVDCx20_ASAP7_75t_R g1948 ( 
.A(n_1406),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1428),
.B(n_1432),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1382),
.B(n_143),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1547),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1372),
.B(n_144),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1626),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1510),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1510),
.Y(n_1955)
);

NOR2xp33_ASAP7_75t_L g1956 ( 
.A(n_1394),
.B(n_144),
.Y(n_1956)
);

INVx2_ASAP7_75t_SL g1957 ( 
.A(n_1343),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1343),
.B(n_145),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1524),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1395),
.B(n_146),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1500),
.B(n_1634),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1635),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1638),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1642),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1543),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1499),
.B(n_419),
.Y(n_1966)
);

CKINVDCx5p33_ASAP7_75t_R g1967 ( 
.A(n_1479),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1524),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1570),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1507),
.B(n_421),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1344),
.B(n_147),
.Y(n_1971)
);

INVx2_ASAP7_75t_SL g1972 ( 
.A(n_1392),
.Y(n_1972)
);

NOR2xp33_ASAP7_75t_L g1973 ( 
.A(n_1404),
.B(n_150),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1608),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1414),
.B(n_151),
.Y(n_1975)
);

BUFx3_ASAP7_75t_L g1976 ( 
.A(n_1628),
.Y(n_1976)
);

XNOR2x2_ASAP7_75t_L g1977 ( 
.A(n_1613),
.B(n_1653),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1643),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1645),
.Y(n_1979)
);

INVxp33_ASAP7_75t_SL g1980 ( 
.A(n_1484),
.Y(n_1980)
);

AOI21x1_ASAP7_75t_L g1981 ( 
.A1(n_1625),
.A2(n_424),
.B(n_422),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1646),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1657),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1508),
.B(n_425),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1671),
.Y(n_1985)
);

AND2x2_ASAP7_75t_SL g1986 ( 
.A(n_1692),
.B(n_1648),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1662),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1675),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1662),
.Y(n_1989)
);

INVx1_ASAP7_75t_SL g1990 ( 
.A(n_1716),
.Y(n_1990)
);

INVx2_ASAP7_75t_L g1991 ( 
.A(n_1672),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1666),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1681),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1693),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1863),
.B(n_1442),
.Y(n_1995)
);

INVx4_ASAP7_75t_L g1996 ( 
.A(n_1953),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1694),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1696),
.B(n_1653),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1819),
.B(n_1440),
.Y(n_1999)
);

NOR2xp33_ASAP7_75t_L g2000 ( 
.A(n_1924),
.B(n_1365),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1818),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1978),
.B(n_1979),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1663),
.B(n_1654),
.Y(n_2003)
);

NOR2xp67_ASAP7_75t_L g2004 ( 
.A(n_1884),
.B(n_1443),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1664),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1876),
.B(n_1654),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1753),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1797),
.B(n_1655),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1978),
.B(n_1467),
.Y(n_2009)
);

AND2x4_ASAP7_75t_SL g2010 ( 
.A(n_1698),
.B(n_1470),
.Y(n_2010)
);

HB1xp67_ASAP7_75t_L g2011 ( 
.A(n_1868),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1845),
.B(n_1387),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1830),
.B(n_1655),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1756),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1785),
.Y(n_2015)
);

HB1xp67_ASAP7_75t_L g2016 ( 
.A(n_1869),
.Y(n_2016)
);

BUFx6f_ASAP7_75t_L g2017 ( 
.A(n_1664),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1666),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1865),
.Y(n_2019)
);

INVx2_ASAP7_75t_L g2020 ( 
.A(n_1793),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1979),
.B(n_1610),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1668),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1974),
.A2(n_1501),
.B(n_1505),
.Y(n_2023)
);

BUFx6f_ASAP7_75t_L g2024 ( 
.A(n_1664),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1706),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1808),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1957),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1982),
.B(n_1373),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1906),
.B(n_1659),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1907),
.B(n_1328),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1706),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1982),
.B(n_1425),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1850),
.B(n_1490),
.Y(n_2033)
);

BUFx3_ASAP7_75t_L g2034 ( 
.A(n_1706),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1674),
.B(n_1632),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1833),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1668),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1676),
.B(n_1554),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_1806),
.B(n_151),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1678),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_1983),
.B(n_1691),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1845),
.B(n_1641),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1669),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1678),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1983),
.B(n_1523),
.Y(n_2045)
);

INVx2_ASAP7_75t_SL g2046 ( 
.A(n_1745),
.Y(n_2046)
);

INVx3_ASAP7_75t_L g2047 ( 
.A(n_1841),
.Y(n_2047)
);

INVx3_ASAP7_75t_L g2048 ( 
.A(n_1669),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1846),
.B(n_1435),
.Y(n_2049)
);

BUFx12f_ASAP7_75t_L g2050 ( 
.A(n_1773),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1918),
.B(n_153),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1859),
.B(n_426),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1925),
.B(n_153),
.Y(n_2053)
);

INVx3_ASAP7_75t_L g2054 ( 
.A(n_1739),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1953),
.B(n_1449),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_L g2056 ( 
.A(n_1953),
.B(n_1630),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1961),
.B(n_155),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1752),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1976),
.B(n_1656),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_1893),
.B(n_156),
.Y(n_2060)
);

OAI21xp5_ASAP7_75t_L g2061 ( 
.A1(n_1974),
.A2(n_1592),
.B(n_1660),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1755),
.Y(n_2062)
);

INVx4_ASAP7_75t_L g2063 ( 
.A(n_1845),
.Y(n_2063)
);

BUFx6f_ASAP7_75t_L g2064 ( 
.A(n_1717),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1894),
.B(n_156),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1882),
.B(n_1661),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1762),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1899),
.B(n_157),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_1717),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1900),
.B(n_157),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_1901),
.B(n_158),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1861),
.B(n_427),
.Y(n_2072)
);

NAND2x1p5_ASAP7_75t_L g2073 ( 
.A(n_1739),
.B(n_1493),
.Y(n_2073)
);

INVx1_ASAP7_75t_SL g2074 ( 
.A(n_1689),
.Y(n_2074)
);

AND2x2_ASAP7_75t_SL g2075 ( 
.A(n_1768),
.B(n_1612),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1688),
.B(n_1619),
.Y(n_2076)
);

BUFx3_ASAP7_75t_L g2077 ( 
.A(n_1717),
.Y(n_2077)
);

INVxp67_ASAP7_75t_L g2078 ( 
.A(n_1937),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1766),
.Y(n_2079)
);

AND2x4_ASAP7_75t_L g2080 ( 
.A(n_1857),
.B(n_428),
.Y(n_2080)
);

INVx2_ASAP7_75t_L g2081 ( 
.A(n_1767),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1903),
.B(n_159),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1904),
.B(n_159),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1882),
.B(n_433),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1772),
.Y(n_2085)
);

INVx2_ASAP7_75t_SL g2086 ( 
.A(n_1704),
.Y(n_2086)
);

AND2x6_ASAP7_75t_L g2087 ( 
.A(n_1968),
.B(n_1413),
.Y(n_2087)
);

INVx3_ASAP7_75t_L g2088 ( 
.A(n_1791),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_1966),
.B(n_1627),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1775),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1780),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1782),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1905),
.B(n_160),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1783),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1828),
.B(n_160),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_1829),
.B(n_161),
.Y(n_2096)
);

INVx3_ASAP7_75t_L g2097 ( 
.A(n_1791),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1677),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_1981),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1679),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1936),
.B(n_163),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_1860),
.Y(n_2102)
);

NOR2xp33_ASAP7_75t_L g2103 ( 
.A(n_1849),
.B(n_1650),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1760),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1966),
.B(n_164),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1984),
.B(n_165),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1916),
.A2(n_436),
.B(n_434),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1680),
.Y(n_2108)
);

AOI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_1798),
.A2(n_170),
.B1(n_165),
.B2(n_167),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1855),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1682),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_1938),
.B(n_170),
.Y(n_2112)
);

INVx1_ASAP7_75t_SL g2113 ( 
.A(n_1952),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1778),
.B(n_438),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1847),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_1813),
.B(n_441),
.Y(n_2116)
);

OR2x2_ASAP7_75t_SL g2117 ( 
.A(n_1685),
.B(n_173),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_1884),
.B(n_445),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1984),
.B(n_174),
.Y(n_2119)
);

INVxp67_ASAP7_75t_L g2120 ( 
.A(n_1950),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1854),
.B(n_447),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_1683),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1673),
.B(n_175),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1848),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1728),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1684),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1686),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1831),
.Y(n_2128)
);

INVx4_ASAP7_75t_L g2129 ( 
.A(n_1728),
.Y(n_2129)
);

CKINVDCx20_ASAP7_75t_R g2130 ( 
.A(n_1731),
.Y(n_2130)
);

INVxp67_ASAP7_75t_L g2131 ( 
.A(n_1920),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1832),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1697),
.Y(n_2133)
);

INVx4_ASAP7_75t_L g2134 ( 
.A(n_1728),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_1771),
.B(n_175),
.Y(n_2135)
);

INVxp67_ASAP7_75t_L g2136 ( 
.A(n_1919),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_1940),
.B(n_176),
.Y(n_2137)
);

AND2x4_ASAP7_75t_L g2138 ( 
.A(n_1856),
.B(n_450),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1805),
.B(n_176),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_1699),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1799),
.B(n_177),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1700),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1702),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1834),
.Y(n_2144)
);

OAI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1968),
.A2(n_452),
.B(n_451),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1862),
.B(n_455),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_1945),
.B(n_178),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1761),
.B(n_457),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1788),
.B(n_460),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1754),
.Y(n_2150)
);

BUFx3_ASAP7_75t_L g2151 ( 
.A(n_1754),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_1695),
.B(n_178),
.Y(n_2152)
);

HB1xp67_ASAP7_75t_L g2153 ( 
.A(n_1836),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1709),
.B(n_180),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_1941),
.B(n_181),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_1816),
.B(n_463),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1837),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1942),
.B(n_181),
.Y(n_2158)
);

HB1xp67_ASAP7_75t_L g2159 ( 
.A(n_1839),
.Y(n_2159)
);

NAND2x1p5_ASAP7_75t_L g2160 ( 
.A(n_1665),
.B(n_465),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1959),
.Y(n_2161)
);

OAI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_1824),
.A2(n_469),
.B(n_468),
.Y(n_2162)
);

AND2x6_ASAP7_75t_L g2163 ( 
.A(n_1935),
.B(n_470),
.Y(n_2163)
);

BUFx3_ASAP7_75t_L g2164 ( 
.A(n_1754),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_1710),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1711),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1822),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1725),
.B(n_475),
.Y(n_2168)
);

INVx2_ASAP7_75t_SL g2169 ( 
.A(n_1757),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1712),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1880),
.B(n_182),
.Y(n_2171)
);

BUFx5_ASAP7_75t_L g2172 ( 
.A(n_1823),
.Y(n_2172)
);

AND2x4_ASAP7_75t_L g2173 ( 
.A(n_1817),
.B(n_476),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1714),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_1949),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_1980),
.B(n_182),
.Y(n_2176)
);

INVxp67_ASAP7_75t_L g2177 ( 
.A(n_1932),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_1757),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1886),
.B(n_183),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1844),
.B(n_477),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1853),
.B(n_479),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1715),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1667),
.B(n_183),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_1962),
.B(n_184),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1721),
.Y(n_2185)
);

INVxp67_ASAP7_75t_SL g2186 ( 
.A(n_1757),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1723),
.Y(n_2187)
);

INVx3_ASAP7_75t_L g2188 ( 
.A(n_1724),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1727),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1729),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1730),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1732),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1733),
.Y(n_2193)
);

AND2x6_ASAP7_75t_L g2194 ( 
.A(n_1870),
.B(n_481),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1708),
.B(n_483),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1713),
.B(n_1740),
.Y(n_2196)
);

INVx2_ASAP7_75t_SL g2197 ( 
.A(n_1892),
.Y(n_2197)
);

BUFx3_ASAP7_75t_L g2198 ( 
.A(n_1814),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1969),
.Y(n_2199)
);

INVx1_ASAP7_75t_SL g2200 ( 
.A(n_1769),
.Y(n_2200)
);

OAI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_1687),
.A2(n_486),
.B(n_485),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1734),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_1944),
.Y(n_2203)
);

BUFx3_ASAP7_75t_L g2204 ( 
.A(n_1815),
.Y(n_2204)
);

NOR2xp33_ASAP7_75t_L g2205 ( 
.A(n_1967),
.B(n_185),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_1963),
.B(n_185),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1735),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1746),
.B(n_491),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1964),
.B(n_186),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_1887),
.B(n_1930),
.Y(n_2210)
);

INVx2_ASAP7_75t_L g2211 ( 
.A(n_1737),
.Y(n_2211)
);

HB1xp67_ASAP7_75t_L g2212 ( 
.A(n_1825),
.Y(n_2212)
);

BUFx3_ASAP7_75t_L g2213 ( 
.A(n_1820),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_1821),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_1902),
.B(n_492),
.Y(n_2215)
);

OAI21xp33_ASAP7_75t_L g2216 ( 
.A1(n_1736),
.A2(n_187),
.B(n_189),
.Y(n_2216)
);

NAND2x1p5_ASAP7_75t_L g2217 ( 
.A(n_1826),
.B(n_1972),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1934),
.B(n_189),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1742),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1726),
.B(n_190),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1747),
.Y(n_2221)
);

INVx4_ASAP7_75t_L g2222 ( 
.A(n_1910),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1787),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_1705),
.B(n_194),
.Y(n_2224)
);

INVx1_ASAP7_75t_SL g2225 ( 
.A(n_1781),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_1744),
.B(n_494),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1852),
.B(n_194),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1929),
.B(n_495),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1958),
.B(n_195),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1878),
.B(n_199),
.Y(n_2230)
);

INVx1_ASAP7_75t_SL g2231 ( 
.A(n_1811),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2027),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_1990),
.B(n_1720),
.Y(n_2233)
);

OR2x2_ASAP7_75t_L g2234 ( 
.A(n_1990),
.B(n_1872),
.Y(n_2234)
);

BUFx6f_ASAP7_75t_L g2235 ( 
.A(n_2017),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2048),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2136),
.B(n_1741),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_2203),
.Y(n_2238)
);

AND2x2_ASAP7_75t_L g2239 ( 
.A(n_2113),
.B(n_1883),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_L g2240 ( 
.A(n_2175),
.B(n_1763),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2054),
.B(n_1921),
.Y(n_2241)
);

OR2x2_ASAP7_75t_L g2242 ( 
.A(n_2113),
.B(n_1873),
.Y(n_2242)
);

NAND2x1_ASAP7_75t_L g2243 ( 
.A(n_1996),
.B(n_1750),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2048),
.Y(n_2244)
);

AND2x4_ASAP7_75t_L g2245 ( 
.A(n_1988),
.B(n_1838),
.Y(n_2245)
);

INVx1_ASAP7_75t_SL g2246 ( 
.A(n_2130),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2054),
.B(n_1875),
.Y(n_2247)
);

INVxp67_ASAP7_75t_L g2248 ( 
.A(n_2011),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1992),
.Y(n_2249)
);

OR2x6_ASAP7_75t_L g2250 ( 
.A(n_2063),
.B(n_1779),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2161),
.Y(n_2251)
);

NOR2xp33_ASAP7_75t_SL g2252 ( 
.A(n_2104),
.B(n_1670),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1996),
.B(n_1914),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2088),
.B(n_1891),
.Y(n_2254)
);

BUFx2_ASAP7_75t_L g2255 ( 
.A(n_2063),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_SL g2256 ( 
.A(n_2223),
.B(n_1842),
.Y(n_2256)
);

CKINVDCx6p67_ASAP7_75t_R g2257 ( 
.A(n_2050),
.Y(n_2257)
);

NOR2xp33_ASAP7_75t_L g2258 ( 
.A(n_2175),
.B(n_1701),
.Y(n_2258)
);

BUFx3_ASAP7_75t_L g2259 ( 
.A(n_2213),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2161),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1992),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2018),
.Y(n_2262)
);

AND2x6_ASAP7_75t_L g2263 ( 
.A(n_2138),
.B(n_1954),
.Y(n_2263)
);

BUFx2_ASAP7_75t_L g2264 ( 
.A(n_2199),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_2087),
.Y(n_2265)
);

NOR2x1_ASAP7_75t_L g2266 ( 
.A(n_2056),
.B(n_2041),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_2017),
.Y(n_2267)
);

HB1xp67_ASAP7_75t_L g2268 ( 
.A(n_2153),
.Y(n_2268)
);

BUFx4f_ASAP7_75t_L g2269 ( 
.A(n_2073),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2016),
.Y(n_2270)
);

BUFx2_ASAP7_75t_L g2271 ( 
.A(n_2087),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2088),
.B(n_2097),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2018),
.Y(n_2273)
);

BUFx2_ASAP7_75t_SL g2274 ( 
.A(n_2005),
.Y(n_2274)
);

AND2x4_ASAP7_75t_L g2275 ( 
.A(n_2198),
.B(n_1951),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2022),
.Y(n_2276)
);

NAND2x1p5_ASAP7_75t_L g2277 ( 
.A(n_2129),
.B(n_1915),
.Y(n_2277)
);

BUFx4f_ASAP7_75t_L g2278 ( 
.A(n_1999),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2022),
.Y(n_2279)
);

INVx5_ASAP7_75t_L g2280 ( 
.A(n_2017),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_2214),
.Y(n_2281)
);

NAND2x1p5_ASAP7_75t_L g2282 ( 
.A(n_2129),
.B(n_1923),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2097),
.B(n_1866),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2196),
.B(n_2002),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2074),
.B(n_1926),
.Y(n_2285)
);

AND2x6_ASAP7_75t_L g2286 ( 
.A(n_2138),
.B(n_1955),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2037),
.Y(n_2287)
);

NAND2x1p5_ASAP7_75t_L g2288 ( 
.A(n_2134),
.B(n_1927),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1987),
.B(n_1858),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2074),
.B(n_1738),
.Y(n_2290)
);

OR2x2_ASAP7_75t_L g2291 ( 
.A(n_2102),
.B(n_1759),
.Y(n_2291)
);

BUFx2_ASAP7_75t_L g2292 ( 
.A(n_2087),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_1987),
.B(n_1764),
.Y(n_2293)
);

INVxp67_ASAP7_75t_L g2294 ( 
.A(n_2197),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2037),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2043),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_1989),
.B(n_1765),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1989),
.B(n_1774),
.Y(n_2298)
);

BUFx4f_ASAP7_75t_L g2299 ( 
.A(n_1999),
.Y(n_2299)
);

HB1xp67_ASAP7_75t_L g2300 ( 
.A(n_2159),
.Y(n_2300)
);

NAND2x1p5_ASAP7_75t_L g2301 ( 
.A(n_2134),
.B(n_1751),
.Y(n_2301)
);

OR2x6_ASAP7_75t_L g2302 ( 
.A(n_2105),
.B(n_1779),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2043),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_2204),
.B(n_1943),
.Y(n_2304)
);

AND2x4_ASAP7_75t_L g2305 ( 
.A(n_2222),
.B(n_1946),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_2031),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_2222),
.B(n_1947),
.Y(n_2307)
);

INVx4_ASAP7_75t_L g2308 ( 
.A(n_2024),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2102),
.B(n_1871),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2212),
.B(n_1794),
.Y(n_2310)
);

INVx4_ASAP7_75t_L g2311 ( 
.A(n_2024),
.Y(n_2311)
);

INVx3_ASAP7_75t_L g2312 ( 
.A(n_2034),
.Y(n_2312)
);

CKINVDCx20_ASAP7_75t_R g2313 ( 
.A(n_2010),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2131),
.B(n_1879),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_2139),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2172),
.B(n_1776),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2172),
.B(n_1777),
.Y(n_2317)
);

BUFx12f_ASAP7_75t_L g2318 ( 
.A(n_2117),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2187),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2172),
.B(n_1722),
.Y(n_2320)
);

BUFx3_ASAP7_75t_L g2321 ( 
.A(n_2077),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2151),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2015),
.Y(n_2323)
);

NOR2xp33_ASAP7_75t_SL g2324 ( 
.A(n_2176),
.B(n_1911),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2177),
.B(n_1800),
.Y(n_2325)
);

NOR2xp33_ASAP7_75t_L g2326 ( 
.A(n_2078),
.B(n_1719),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2172),
.B(n_2019),
.Y(n_2327)
);

BUFx4f_ASAP7_75t_SL g2328 ( 
.A(n_2012),
.Y(n_2328)
);

AND2x6_ASAP7_75t_L g2329 ( 
.A(n_2146),
.B(n_1803),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2020),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_2187),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2026),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2120),
.B(n_1881),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_2087),
.Y(n_2334)
);

AND2x4_ASAP7_75t_L g2335 ( 
.A(n_2210),
.B(n_1795),
.Y(n_2335)
);

OR2x6_ASAP7_75t_SL g2336 ( 
.A(n_2066),
.B(n_1965),
.Y(n_2336)
);

OR2x6_ASAP7_75t_L g2337 ( 
.A(n_2106),
.B(n_1909),
.Y(n_2337)
);

BUFx6f_ASAP7_75t_L g2338 ( 
.A(n_2024),
.Y(n_2338)
);

CKINVDCx20_ASAP7_75t_R g2339 ( 
.A(n_2000),
.Y(n_2339)
);

INVx1_ASAP7_75t_L g2340 ( 
.A(n_2191),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_L g2341 ( 
.A(n_2172),
.B(n_1885),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2191),
.Y(n_2342)
);

AND2x4_ASAP7_75t_L g2343 ( 
.A(n_2164),
.B(n_1804),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2019),
.B(n_1888),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2033),
.B(n_1890),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2046),
.B(n_1896),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2110),
.B(n_1827),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2192),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2001),
.B(n_1809),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2036),
.B(n_1810),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2135),
.B(n_1971),
.Y(n_2351)
);

NAND2x1_ASAP7_75t_L g2352 ( 
.A(n_2163),
.B(n_1928),
.Y(n_2352)
);

BUFx2_ASAP7_75t_L g2353 ( 
.A(n_2220),
.Y(n_2353)
);

INVx3_ASAP7_75t_L g2354 ( 
.A(n_2025),
.Y(n_2354)
);

BUFx3_ASAP7_75t_L g2355 ( 
.A(n_2217),
.Y(n_2355)
);

AND2x4_ASAP7_75t_L g2356 ( 
.A(n_2127),
.B(n_1786),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_2110),
.B(n_1864),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2009),
.B(n_1874),
.Y(n_2358)
);

BUFx2_ASAP7_75t_L g2359 ( 
.A(n_2147),
.Y(n_2359)
);

NOR2xp67_ASAP7_75t_L g2360 ( 
.A(n_2086),
.B(n_2055),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1985),
.Y(n_2361)
);

BUFx2_ASAP7_75t_L g2362 ( 
.A(n_2025),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2192),
.Y(n_2363)
);

BUFx4f_ASAP7_75t_L g2364 ( 
.A(n_2156),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2029),
.B(n_1956),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_2183),
.B(n_1970),
.Y(n_2366)
);

AND2x4_ASAP7_75t_L g2367 ( 
.A(n_2133),
.B(n_1789),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2152),
.B(n_1960),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2219),
.Y(n_2369)
);

BUFx2_ASAP7_75t_L g2370 ( 
.A(n_2227),
.Y(n_2370)
);

BUFx8_ASAP7_75t_L g2371 ( 
.A(n_2038),
.Y(n_2371)
);

AND2x2_ASAP7_75t_L g2372 ( 
.A(n_2057),
.B(n_2030),
.Y(n_2372)
);

INVxp67_ASAP7_75t_L g2373 ( 
.A(n_2206),
.Y(n_2373)
);

BUFx4f_ASAP7_75t_L g2374 ( 
.A(n_2156),
.Y(n_2374)
);

OR2x6_ASAP7_75t_L g2375 ( 
.A(n_2119),
.B(n_1909),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2080),
.B(n_1758),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_2137),
.B(n_1703),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_2154),
.B(n_1973),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2035),
.B(n_1770),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2080),
.B(n_1975),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2025),
.Y(n_2381)
);

AND2x2_ASAP7_75t_L g2382 ( 
.A(n_2049),
.B(n_1748),
.Y(n_2382)
);

OR2x6_ASAP7_75t_L g2383 ( 
.A(n_2146),
.B(n_1917),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2219),
.Y(n_2384)
);

NAND2x1p5_ASAP7_75t_L g2385 ( 
.A(n_2064),
.B(n_1792),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_2064),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_1991),
.Y(n_2387)
);

CKINVDCx20_ASAP7_75t_R g2388 ( 
.A(n_2042),
.Y(n_2388)
);

INVx2_ASAP7_75t_L g2389 ( 
.A(n_1993),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2021),
.B(n_1931),
.Y(n_2390)
);

AND2x4_ASAP7_75t_L g2391 ( 
.A(n_2140),
.B(n_1807),
.Y(n_2391)
);

INVx2_ASAP7_75t_SL g2392 ( 
.A(n_2234),
.Y(n_2392)
);

NAND2x1p5_ASAP7_75t_L g2393 ( 
.A(n_2280),
.B(n_2064),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2261),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2249),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2264),
.Y(n_2396)
);

NAND2x1p5_ASAP7_75t_L g2397 ( 
.A(n_2280),
.B(n_2069),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2245),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2284),
.B(n_2059),
.Y(n_2399)
);

NAND2x1p5_ASAP7_75t_L g2400 ( 
.A(n_2255),
.B(n_2069),
.Y(n_2400)
);

INVx3_ASAP7_75t_SL g2401 ( 
.A(n_2257),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2262),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2273),
.Y(n_2403)
);

BUFx3_ASAP7_75t_L g2404 ( 
.A(n_2259),
.Y(n_2404)
);

INVx5_ASAP7_75t_L g2405 ( 
.A(n_2250),
.Y(n_2405)
);

NAND2x1p5_ASAP7_75t_L g2406 ( 
.A(n_2308),
.B(n_2069),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2276),
.Y(n_2407)
);

INVx5_ASAP7_75t_L g2408 ( 
.A(n_2250),
.Y(n_2408)
);

BUFx6f_ASAP7_75t_L g2409 ( 
.A(n_2235),
.Y(n_2409)
);

INVx3_ASAP7_75t_L g2410 ( 
.A(n_2236),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2279),
.Y(n_2411)
);

INVx4_ASAP7_75t_L g2412 ( 
.A(n_2235),
.Y(n_2412)
);

BUFx3_ASAP7_75t_L g2413 ( 
.A(n_2264),
.Y(n_2413)
);

INVx6_ASAP7_75t_SL g2414 ( 
.A(n_2383),
.Y(n_2414)
);

INVx1_ASAP7_75t_SL g2415 ( 
.A(n_2233),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_2306),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_2321),
.Y(n_2417)
);

BUFx3_ASAP7_75t_L g2418 ( 
.A(n_2391),
.Y(n_2418)
);

BUFx2_ASAP7_75t_L g2419 ( 
.A(n_2370),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2358),
.B(n_2141),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2345),
.B(n_1998),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2370),
.Y(n_2422)
);

BUFx6f_ASAP7_75t_L g2423 ( 
.A(n_2267),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_2365),
.B(n_2103),
.Y(n_2424)
);

BUFx6f_ASAP7_75t_L g2425 ( 
.A(n_2267),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_2244),
.Y(n_2426)
);

INVx2_ASAP7_75t_L g2427 ( 
.A(n_2303),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2287),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2295),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2278),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2338),
.Y(n_2431)
);

BUFx6f_ASAP7_75t_L g2432 ( 
.A(n_2338),
.Y(n_2432)
);

INVxp67_ASAP7_75t_SL g2433 ( 
.A(n_2327),
.Y(n_2433)
);

BUFx3_ASAP7_75t_L g2434 ( 
.A(n_2313),
.Y(n_2434)
);

AND2x2_ASAP7_75t_L g2435 ( 
.A(n_2372),
.B(n_2184),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2296),
.Y(n_2436)
);

BUFx12f_ASAP7_75t_L g2437 ( 
.A(n_2371),
.Y(n_2437)
);

BUFx3_ASAP7_75t_L g2438 ( 
.A(n_2355),
.Y(n_2438)
);

INVx4_ASAP7_75t_L g2439 ( 
.A(n_2381),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2319),
.Y(n_2440)
);

INVx1_ASAP7_75t_SL g2441 ( 
.A(n_2233),
.Y(n_2441)
);

INVx3_ASAP7_75t_SL g2442 ( 
.A(n_2246),
.Y(n_2442)
);

AND2x6_ASAP7_75t_L g2443 ( 
.A(n_2266),
.B(n_2052),
.Y(n_2443)
);

CKINVDCx5p33_ASAP7_75t_R g2444 ( 
.A(n_2339),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2344),
.B(n_2123),
.Y(n_2445)
);

INVx8_ASAP7_75t_L g2446 ( 
.A(n_2381),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2304),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_2331),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_2368),
.B(n_2200),
.Y(n_2449)
);

INVx1_ASAP7_75t_SL g2450 ( 
.A(n_2234),
.Y(n_2450)
);

NAND2x1p5_ASAP7_75t_L g2451 ( 
.A(n_2311),
.B(n_2125),
.Y(n_2451)
);

NAND2x1p5_ASAP7_75t_L g2452 ( 
.A(n_2312),
.B(n_2125),
.Y(n_2452)
);

HB1xp67_ASAP7_75t_L g2453 ( 
.A(n_2268),
.Y(n_2453)
);

BUFx3_ASAP7_75t_L g2454 ( 
.A(n_2232),
.Y(n_2454)
);

INVx2_ASAP7_75t_SL g2455 ( 
.A(n_2300),
.Y(n_2455)
);

BUFx6f_ASAP7_75t_L g2456 ( 
.A(n_2275),
.Y(n_2456)
);

AOI22xp33_ASAP7_75t_L g2457 ( 
.A1(n_2329),
.A2(n_1986),
.B1(n_2076),
.B2(n_2089),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_2322),
.Y(n_2458)
);

INVx3_ASAP7_75t_SL g2459 ( 
.A(n_2291),
.Y(n_2459)
);

BUFx5_ASAP7_75t_L g2460 ( 
.A(n_2340),
.Y(n_2460)
);

BUFx3_ASAP7_75t_L g2461 ( 
.A(n_2310),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2251),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2362),
.Y(n_2463)
);

INVx8_ASAP7_75t_L g2464 ( 
.A(n_2263),
.Y(n_2464)
);

INVxp67_ASAP7_75t_SL g2465 ( 
.A(n_2341),
.Y(n_2465)
);

INVx6_ASAP7_75t_L g2466 ( 
.A(n_2318),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_2378),
.B(n_2155),
.Y(n_2467)
);

INVx1_ASAP7_75t_SL g2468 ( 
.A(n_2291),
.Y(n_2468)
);

BUFx3_ASAP7_75t_L g2469 ( 
.A(n_2281),
.Y(n_2469)
);

CKINVDCx5p33_ASAP7_75t_R g2470 ( 
.A(n_2269),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2386),
.Y(n_2471)
);

BUFx6f_ASAP7_75t_L g2472 ( 
.A(n_2299),
.Y(n_2472)
);

INVx3_ASAP7_75t_L g2473 ( 
.A(n_2343),
.Y(n_2473)
);

INVx3_ASAP7_75t_L g2474 ( 
.A(n_2335),
.Y(n_2474)
);

INVx1_ASAP7_75t_SL g2475 ( 
.A(n_2353),
.Y(n_2475)
);

INVx6_ASAP7_75t_L g2476 ( 
.A(n_2383),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2342),
.Y(n_2477)
);

INVx2_ASAP7_75t_R g2478 ( 
.A(n_2348),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_2285),
.Y(n_2479)
);

INVx3_ASAP7_75t_SL g2480 ( 
.A(n_2309),
.Y(n_2480)
);

BUFx3_ASAP7_75t_L g2481 ( 
.A(n_2336),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2333),
.B(n_2209),
.Y(n_2482)
);

INVx2_ASAP7_75t_SL g2483 ( 
.A(n_2242),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2363),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2354),
.Y(n_2485)
);

BUFx6f_ASAP7_75t_L g2486 ( 
.A(n_2305),
.Y(n_2486)
);

INVx1_ASAP7_75t_SL g2487 ( 
.A(n_2309),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2293),
.B(n_2158),
.Y(n_2488)
);

NAND2x1p5_ASAP7_75t_L g2489 ( 
.A(n_2364),
.B(n_2125),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2260),
.Y(n_2490)
);

INVx5_ASAP7_75t_L g2491 ( 
.A(n_2263),
.Y(n_2491)
);

INVx8_ASAP7_75t_L g2492 ( 
.A(n_2263),
.Y(n_2492)
);

CKINVDCx20_ASAP7_75t_R g2493 ( 
.A(n_2388),
.Y(n_2493)
);

INVx1_ASAP7_75t_SL g2494 ( 
.A(n_2379),
.Y(n_2494)
);

BUFx3_ASAP7_75t_L g2495 ( 
.A(n_2349),
.Y(n_2495)
);

BUFx2_ASAP7_75t_L g2496 ( 
.A(n_2413),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2440),
.Y(n_2497)
);

AOI22xp33_ASAP7_75t_SL g2498 ( 
.A1(n_2424),
.A2(n_2324),
.B1(n_2382),
.B2(n_2377),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2440),
.Y(n_2499)
);

CKINVDCx11_ASAP7_75t_R g2500 ( 
.A(n_2401),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2448),
.Y(n_2501)
);

BUFx2_ASAP7_75t_L g2502 ( 
.A(n_2396),
.Y(n_2502)
);

AOI22xp33_ASAP7_75t_L g2503 ( 
.A1(n_2457),
.A2(n_2329),
.B1(n_2237),
.B2(n_2376),
.Y(n_2503)
);

OAI22xp33_ASAP7_75t_L g2504 ( 
.A1(n_2480),
.A2(n_2252),
.B1(n_2256),
.B2(n_2240),
.Y(n_2504)
);

OAI22xp33_ASAP7_75t_L g2505 ( 
.A1(n_2487),
.A2(n_2328),
.B1(n_2380),
.B2(n_2200),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2448),
.Y(n_2506)
);

BUFx12f_ASAP7_75t_L g2507 ( 
.A(n_2437),
.Y(n_2507)
);

BUFx12f_ASAP7_75t_L g2508 ( 
.A(n_2470),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2477),
.Y(n_2509)
);

AO22x1_ASAP7_75t_L g2510 ( 
.A1(n_2443),
.A2(n_2205),
.B1(n_2258),
.B2(n_2329),
.Y(n_2510)
);

INVx6_ASAP7_75t_L g2511 ( 
.A(n_2405),
.Y(n_2511)
);

OAI22xp5_ASAP7_75t_L g2512 ( 
.A1(n_2488),
.A2(n_2374),
.B1(n_2317),
.B2(n_2316),
.Y(n_2512)
);

CKINVDCx5p33_ASAP7_75t_R g2513 ( 
.A(n_2444),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2477),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_L g2515 ( 
.A1(n_2421),
.A2(n_1718),
.B1(n_2359),
.B2(n_1877),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2484),
.Y(n_2516)
);

BUFx6f_ASAP7_75t_L g2517 ( 
.A(n_2409),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2484),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_2399),
.B(n_2314),
.Y(n_2519)
);

AOI22xp33_ASAP7_75t_SL g2520 ( 
.A1(n_2430),
.A2(n_2075),
.B1(n_2325),
.B2(n_1948),
.Y(n_2520)
);

INVx4_ASAP7_75t_L g2521 ( 
.A(n_2446),
.Y(n_2521)
);

AOI22xp33_ASAP7_75t_L g2522 ( 
.A1(n_2482),
.A2(n_1897),
.B1(n_1898),
.B2(n_1812),
.Y(n_2522)
);

BUFx2_ASAP7_75t_SL g2523 ( 
.A(n_2404),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_2420),
.B(n_2297),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_SL g2525 ( 
.A1(n_2465),
.A2(n_2145),
.B(n_2162),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2442),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2435),
.B(n_2346),
.Y(n_2527)
);

BUFx2_ASAP7_75t_L g2528 ( 
.A(n_2419),
.Y(n_2528)
);

INVx6_ASAP7_75t_L g2529 ( 
.A(n_2405),
.Y(n_2529)
);

INVx3_ASAP7_75t_L g2530 ( 
.A(n_2464),
.Y(n_2530)
);

BUFx10_ASAP7_75t_L g2531 ( 
.A(n_2466),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_L g2532 ( 
.A1(n_2494),
.A2(n_1912),
.B1(n_2292),
.B2(n_2271),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2394),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2394),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2428),
.Y(n_2535)
);

INVx2_ASAP7_75t_L g2536 ( 
.A(n_2402),
.Y(n_2536)
);

OR2x2_ASAP7_75t_L g2537 ( 
.A(n_2449),
.B(n_2242),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2402),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2403),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_2419),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2403),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2415),
.A2(n_2334),
.B1(n_2265),
.B2(n_1707),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2407),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2407),
.Y(n_2544)
);

OR2x2_ASAP7_75t_L g2545 ( 
.A(n_2468),
.B(n_2298),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2411),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2467),
.B(n_2351),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2445),
.B(n_2373),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2411),
.Y(n_2549)
);

AOI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2441),
.A2(n_2265),
.B1(n_2326),
.B2(n_2225),
.Y(n_2550)
);

CKINVDCx5p33_ASAP7_75t_R g2551 ( 
.A(n_2434),
.Y(n_2551)
);

AOI22xp33_ASAP7_75t_SL g2552 ( 
.A1(n_2430),
.A2(n_1933),
.B1(n_2231),
.B2(n_2225),
.Y(n_2552)
);

BUFx2_ASAP7_75t_L g2553 ( 
.A(n_2422),
.Y(n_2553)
);

BUFx4f_ASAP7_75t_L g2554 ( 
.A(n_2472),
.Y(n_2554)
);

AOI22xp5_ASAP7_75t_SL g2555 ( 
.A1(n_2493),
.A2(n_1939),
.B1(n_1802),
.B2(n_2231),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2429),
.Y(n_2556)
);

BUFx3_ASAP7_75t_L g2557 ( 
.A(n_2438),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2429),
.Y(n_2558)
);

OAI22xp5_ASAP7_75t_SL g2559 ( 
.A1(n_2459),
.A2(n_2109),
.B1(n_1917),
.B2(n_2337),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2436),
.Y(n_2560)
);

OAI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_2433),
.A2(n_2366),
.B1(n_2347),
.B2(n_2357),
.Y(n_2561)
);

BUFx3_ASAP7_75t_L g2562 ( 
.A(n_2398),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_2479),
.A2(n_2216),
.B1(n_1867),
.B2(n_1913),
.Y(n_2563)
);

BUFx3_ASAP7_75t_L g2564 ( 
.A(n_2418),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2483),
.B(n_2239),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2436),
.Y(n_2566)
);

AOI22xp5_ASAP7_75t_L g2567 ( 
.A1(n_2443),
.A2(n_2216),
.B1(n_2290),
.B2(n_2241),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2462),
.Y(n_2568)
);

OAI21xp5_ASAP7_75t_SL g2569 ( 
.A1(n_2450),
.A2(n_2109),
.B(n_1851),
.Y(n_2569)
);

INVx2_ASAP7_75t_SL g2570 ( 
.A(n_2446),
.Y(n_2570)
);

INVx1_ASAP7_75t_L g2571 ( 
.A(n_2490),
.Y(n_2571)
);

INVx3_ASAP7_75t_L g2572 ( 
.A(n_2464),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2395),
.Y(n_2573)
);

INVx3_ASAP7_75t_L g2574 ( 
.A(n_2492),
.Y(n_2574)
);

AOI22xp33_ASAP7_75t_L g2575 ( 
.A1(n_2443),
.A2(n_2337),
.B1(n_2375),
.B2(n_2084),
.Y(n_2575)
);

CKINVDCx5p33_ASAP7_75t_R g2576 ( 
.A(n_2414),
.Y(n_2576)
);

INVx6_ASAP7_75t_L g2577 ( 
.A(n_2405),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_SL g2578 ( 
.A1(n_2555),
.A2(n_2481),
.B1(n_1977),
.B2(n_2163),
.Y(n_2578)
);

OAI21xp5_ASAP7_75t_SL g2579 ( 
.A1(n_2569),
.A2(n_1843),
.B(n_1922),
.Y(n_2579)
);

INVx2_ASAP7_75t_L g2580 ( 
.A(n_2536),
.Y(n_2580)
);

AOI22xp33_ASAP7_75t_L g2581 ( 
.A1(n_2559),
.A2(n_1895),
.B1(n_2253),
.B2(n_2107),
.Y(n_2581)
);

AOI22xp33_ASAP7_75t_SL g2582 ( 
.A1(n_2555),
.A2(n_2163),
.B1(n_2194),
.B2(n_2229),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2497),
.Y(n_2583)
);

OAI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2503),
.A2(n_2392),
.B1(n_2360),
.B2(n_2422),
.Y(n_2584)
);

OAI21xp33_ASAP7_75t_L g2585 ( 
.A1(n_2519),
.A2(n_1908),
.B(n_2028),
.Y(n_2585)
);

AOI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2498),
.A2(n_2472),
.B1(n_2302),
.B2(n_1790),
.Y(n_2586)
);

INVxp67_ASAP7_75t_L g2587 ( 
.A(n_2502),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2504),
.B(n_2460),
.Y(n_2588)
);

OAI22xp33_ASAP7_75t_L g2589 ( 
.A1(n_2569),
.A2(n_2375),
.B1(n_2302),
.B2(n_2475),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2499),
.Y(n_2590)
);

INVx5_ASAP7_75t_SL g2591 ( 
.A(n_2517),
.Y(n_2591)
);

AOI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2559),
.A2(n_2201),
.B1(n_2163),
.B2(n_2116),
.Y(n_2592)
);

BUFx2_ASAP7_75t_L g2593 ( 
.A(n_2496),
.Y(n_2593)
);

OAI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2550),
.A2(n_2315),
.B1(n_2384),
.B2(n_2369),
.Y(n_2594)
);

AOI22xp5_ASAP7_75t_L g2595 ( 
.A1(n_2522),
.A2(n_1749),
.B1(n_2474),
.B2(n_2473),
.Y(n_2595)
);

AND2x2_ASAP7_75t_L g2596 ( 
.A(n_2527),
.B(n_2003),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2524),
.B(n_2455),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2547),
.B(n_2006),
.Y(n_2598)
);

OAI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2563),
.A2(n_2552),
.B1(n_2532),
.B2(n_2542),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2501),
.Y(n_2600)
);

OAI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2575),
.A2(n_2238),
.B1(n_2454),
.B2(n_2282),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2515),
.A2(n_2288),
.B1(n_2277),
.B2(n_2476),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2548),
.B(n_2537),
.Y(n_2603)
);

AOI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_2520),
.A2(n_2116),
.B1(n_2168),
.B2(n_2194),
.Y(n_2604)
);

OAI222xp33_ASAP7_75t_L g2605 ( 
.A1(n_2567),
.A2(n_1784),
.B1(n_2390),
.B2(n_2032),
.C1(n_2427),
.C2(n_2289),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_SL g2606 ( 
.A1(n_2577),
.A2(n_2194),
.B1(n_2408),
.B2(n_2023),
.Y(n_2606)
);

NAND2xp5_ASAP7_75t_L g2607 ( 
.A(n_2545),
.B(n_2565),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2506),
.Y(n_2608)
);

INVx1_ASAP7_75t_SL g2609 ( 
.A(n_2528),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2538),
.Y(n_2610)
);

OAI22xp5_ASAP7_75t_L g2611 ( 
.A1(n_2505),
.A2(n_2476),
.B1(n_2491),
.B2(n_2294),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2540),
.B(n_2008),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2553),
.Y(n_2613)
);

AOI22xp33_ASAP7_75t_L g2614 ( 
.A1(n_2512),
.A2(n_2194),
.B1(n_2096),
.B2(n_2095),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2539),
.Y(n_2615)
);

AOI222xp33_ASAP7_75t_L g2616 ( 
.A1(n_2510),
.A2(n_2061),
.B1(n_2068),
.B2(n_2070),
.C1(n_2065),
.C2(n_2060),
.Y(n_2616)
);

HB1xp67_ASAP7_75t_L g2617 ( 
.A(n_2564),
.Y(n_2617)
);

AOI22xp33_ASAP7_75t_SL g2618 ( 
.A1(n_2577),
.A2(n_2408),
.B1(n_1840),
.B2(n_2466),
.Y(n_2618)
);

OAI22xp33_ASAP7_75t_L g2619 ( 
.A1(n_2567),
.A2(n_2408),
.B1(n_2491),
.B2(n_2456),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2509),
.Y(n_2620)
);

HB1xp67_ASAP7_75t_L g2621 ( 
.A(n_2562),
.Y(n_2621)
);

OAI222xp33_ASAP7_75t_L g2622 ( 
.A1(n_2561),
.A2(n_2283),
.B1(n_2453),
.B2(n_2254),
.C1(n_2247),
.C2(n_2270),
.Y(n_2622)
);

HB1xp67_ASAP7_75t_L g2623 ( 
.A(n_2517),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2566),
.Y(n_2624)
);

OAI21xp5_ASAP7_75t_SL g2625 ( 
.A1(n_2568),
.A2(n_2082),
.B(n_2071),
.Y(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2535),
.A2(n_2093),
.B1(n_2083),
.B2(n_2039),
.Y(n_2626)
);

INVx2_ASAP7_75t_SL g2627 ( 
.A(n_2554),
.Y(n_2627)
);

AOI22xp33_ASAP7_75t_L g2628 ( 
.A1(n_2573),
.A2(n_2053),
.B1(n_2051),
.B2(n_2286),
.Y(n_2628)
);

OAI22xp5_ASAP7_75t_SL g2629 ( 
.A1(n_2526),
.A2(n_2469),
.B1(n_2489),
.B2(n_2471),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_SL g2630 ( 
.A1(n_2511),
.A2(n_2286),
.B1(n_2492),
.B2(n_2460),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2571),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_2511),
.A2(n_2286),
.B1(n_2121),
.B2(n_2112),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2525),
.A2(n_2491),
.B1(n_2248),
.B2(n_2400),
.Y(n_2633)
);

AOI22xp33_ASAP7_75t_L g2634 ( 
.A1(n_2529),
.A2(n_2121),
.B1(n_2101),
.B2(n_2224),
.Y(n_2634)
);

INVx3_ASAP7_75t_L g2635 ( 
.A(n_2530),
.Y(n_2635)
);

OAI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2529),
.A2(n_2320),
.B1(n_2274),
.B2(n_2495),
.Y(n_2636)
);

CKINVDCx20_ASAP7_75t_R g2637 ( 
.A(n_2500),
.Y(n_2637)
);

AOI22xp33_ASAP7_75t_SL g2638 ( 
.A1(n_2523),
.A2(n_2460),
.B1(n_2461),
.B2(n_2456),
.Y(n_2638)
);

OAI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2514),
.A2(n_2452),
.B1(n_2397),
.B2(n_2393),
.Y(n_2639)
);

OAI21xp33_ASAP7_75t_L g2640 ( 
.A1(n_2516),
.A2(n_2045),
.B(n_2058),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2517),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2518),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2533),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2534),
.A2(n_2541),
.B1(n_2544),
.B2(n_2543),
.Y(n_2644)
);

OAI22xp5_ASAP7_75t_L g2645 ( 
.A1(n_2546),
.A2(n_2174),
.B1(n_2188),
.B2(n_1995),
.Y(n_2645)
);

NAND3xp33_ASAP7_75t_L g2646 ( 
.A(n_2549),
.B(n_1801),
.C(n_2148),
.Y(n_2646)
);

BUFx8_ASAP7_75t_L g2647 ( 
.A(n_2507),
.Y(n_2647)
);

NAND2xp5_ASAP7_75t_SL g2648 ( 
.A(n_2513),
.B(n_2460),
.Y(n_2648)
);

OAI21xp33_ASAP7_75t_L g2649 ( 
.A1(n_2556),
.A2(n_2067),
.B(n_2058),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2558),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2560),
.Y(n_2651)
);

INVx1_ASAP7_75t_SL g2652 ( 
.A(n_2557),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2530),
.A2(n_2188),
.B1(n_2174),
.B2(n_2149),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2551),
.A2(n_2447),
.B1(n_2486),
.B2(n_2367),
.Y(n_2654)
);

OR2x2_ASAP7_75t_L g2655 ( 
.A(n_2572),
.B(n_2463),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2572),
.Y(n_2656)
);

AOI22xp33_ASAP7_75t_SL g2657 ( 
.A1(n_2508),
.A2(n_2554),
.B1(n_2531),
.B2(n_2447),
.Y(n_2657)
);

INVxp67_ASAP7_75t_L g2658 ( 
.A(n_2570),
.Y(n_2658)
);

AOI22xp33_ASAP7_75t_SL g2659 ( 
.A1(n_2531),
.A2(n_2230),
.B1(n_2218),
.B2(n_2463),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2574),
.Y(n_2660)
);

AOI222xp33_ASAP7_75t_L g2661 ( 
.A1(n_2576),
.A2(n_2171),
.B1(n_2179),
.B2(n_2167),
.C1(n_2013),
.C2(n_2115),
.Y(n_2661)
);

AOI22xp33_ASAP7_75t_L g2662 ( 
.A1(n_2599),
.A2(n_2067),
.B1(n_2085),
.B2(n_2079),
.Y(n_2662)
);

AOI22xp33_ASAP7_75t_SL g2663 ( 
.A1(n_2602),
.A2(n_2574),
.B1(n_2160),
.B2(n_2228),
.Y(n_2663)
);

AOI22xp33_ASAP7_75t_L g2664 ( 
.A1(n_2581),
.A2(n_2079),
.B1(n_2090),
.B2(n_2085),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_L g2665 ( 
.A1(n_2578),
.A2(n_2094),
.B1(n_2090),
.B2(n_2478),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2585),
.A2(n_2094),
.B1(n_2173),
.B2(n_2081),
.Y(n_2666)
);

AOI22xp33_ASAP7_75t_L g2667 ( 
.A1(n_2616),
.A2(n_2215),
.B1(n_2114),
.B2(n_2181),
.Y(n_2667)
);

AOI22xp33_ASAP7_75t_L g2668 ( 
.A1(n_2592),
.A2(n_2180),
.B1(n_2208),
.B2(n_2195),
.Y(n_2668)
);

AOI22xp33_ASAP7_75t_SL g2669 ( 
.A1(n_2611),
.A2(n_2173),
.B1(n_2052),
.B2(n_2072),
.Y(n_2669)
);

OAI21xp33_ASAP7_75t_L g2670 ( 
.A1(n_2625),
.A2(n_2661),
.B(n_2626),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2659),
.A2(n_2301),
.B1(n_2414),
.B2(n_2385),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2603),
.B(n_2410),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_L g2673 ( 
.A1(n_2582),
.A2(n_2226),
.B1(n_2142),
.B2(n_2165),
.Y(n_2673)
);

AOI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_2588),
.A2(n_2226),
.B1(n_2143),
.B2(n_2170),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2604),
.A2(n_2166),
.B1(n_2185),
.B2(n_2182),
.Y(n_2675)
);

AOI22xp33_ASAP7_75t_SL g2676 ( 
.A1(n_2584),
.A2(n_2072),
.B1(n_2486),
.B2(n_2417),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2589),
.A2(n_2189),
.B1(n_2193),
.B2(n_2190),
.Y(n_2677)
);

AOI22xp33_ASAP7_75t_L g2678 ( 
.A1(n_2619),
.A2(n_2202),
.B1(n_2211),
.B2(n_2207),
.Y(n_2678)
);

OAI22xp5_ASAP7_75t_L g2679 ( 
.A1(n_2586),
.A2(n_2521),
.B1(n_2272),
.B2(n_2458),
.Y(n_2679)
);

OAI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_2634),
.A2(n_2521),
.B1(n_2410),
.B2(n_2426),
.Y(n_2680)
);

AOI22xp5_ASAP7_75t_L g2681 ( 
.A1(n_2579),
.A2(n_2356),
.B1(n_2004),
.B2(n_2221),
.Y(n_2681)
);

AOI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_2614),
.A2(n_2111),
.B1(n_2100),
.B2(n_2108),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2607),
.B(n_2426),
.Y(n_2683)
);

OAI21xp5_ASAP7_75t_L g2684 ( 
.A1(n_2625),
.A2(n_1690),
.B(n_2118),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2597),
.B(n_2323),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2631),
.Y(n_2686)
);

OAI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2632),
.A2(n_2485),
.B1(n_2412),
.B2(n_2439),
.Y(n_2687)
);

AOI22xp33_ASAP7_75t_L g2688 ( 
.A1(n_2598),
.A2(n_2111),
.B1(n_2122),
.B2(n_2098),
.Y(n_2688)
);

AOI222xp33_ASAP7_75t_L g2689 ( 
.A1(n_2579),
.A2(n_2167),
.B1(n_2091),
.B2(n_2062),
.C1(n_2092),
.C2(n_2124),
.Y(n_2689)
);

CKINVDCx5p33_ASAP7_75t_R g2690 ( 
.A(n_2637),
.Y(n_2690)
);

AOI22xp33_ASAP7_75t_L g2691 ( 
.A1(n_2606),
.A2(n_2126),
.B1(n_2047),
.B2(n_2330),
.Y(n_2691)
);

AOI22xp33_ASAP7_75t_L g2692 ( 
.A1(n_2618),
.A2(n_2047),
.B1(n_2361),
.B2(n_2332),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2596),
.B(n_2307),
.Y(n_2693)
);

AOI22xp33_ASAP7_75t_L g2694 ( 
.A1(n_2601),
.A2(n_2387),
.B1(n_2389),
.B2(n_2352),
.Y(n_2694)
);

BUFx2_ASAP7_75t_L g2695 ( 
.A(n_2593),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_L g2696 ( 
.A1(n_2640),
.A2(n_1796),
.B1(n_1835),
.B2(n_1743),
.Y(n_2696)
);

AOI22xp33_ASAP7_75t_L g2697 ( 
.A1(n_2628),
.A2(n_1889),
.B1(n_2044),
.B2(n_2040),
.Y(n_2697)
);

AOI22xp33_ASAP7_75t_L g2698 ( 
.A1(n_2633),
.A2(n_1994),
.B1(n_2007),
.B2(n_1997),
.Y(n_2698)
);

OAI222xp33_ASAP7_75t_L g2699 ( 
.A1(n_2587),
.A2(n_2115),
.B1(n_2124),
.B2(n_2157),
.C1(n_2128),
.C2(n_2132),
.Y(n_2699)
);

OAI222xp33_ASAP7_75t_L g2700 ( 
.A1(n_2609),
.A2(n_2128),
.B1(n_2132),
.B2(n_2144),
.C1(n_2157),
.C2(n_2406),
.Y(n_2700)
);

AOI222xp33_ASAP7_75t_L g2701 ( 
.A1(n_2605),
.A2(n_2144),
.B1(n_2350),
.B2(n_2014),
.C1(n_1994),
.C2(n_2169),
.Y(n_2701)
);

AOI22xp33_ASAP7_75t_SL g2702 ( 
.A1(n_2636),
.A2(n_2416),
.B1(n_2439),
.B2(n_2412),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_L g2703 ( 
.A(n_2613),
.B(n_2409),
.Y(n_2703)
);

OAI22xp5_ASAP7_75t_L g2704 ( 
.A1(n_2654),
.A2(n_2451),
.B1(n_2186),
.B2(n_2425),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2648),
.A2(n_2243),
.B1(n_2150),
.B2(n_2178),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2612),
.A2(n_2150),
.B1(n_2178),
.B2(n_2004),
.Y(n_2706)
);

AOI221xp5_ASAP7_75t_L g2707 ( 
.A1(n_2622),
.A2(n_2432),
.B1(n_2431),
.B2(n_2425),
.C(n_2423),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_SL g2708 ( 
.A1(n_2629),
.A2(n_2646),
.B1(n_2594),
.B2(n_2621),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2649),
.A2(n_2150),
.B1(n_2178),
.B2(n_2099),
.Y(n_2709)
);

AOI22xp33_ASAP7_75t_L g2710 ( 
.A1(n_2617),
.A2(n_2099),
.B1(n_2431),
.B2(n_2423),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2583),
.Y(n_2711)
);

AOI22xp33_ASAP7_75t_L g2712 ( 
.A1(n_2595),
.A2(n_2432),
.B1(n_203),
.B2(n_201),
.Y(n_2712)
);

AOI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2638),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2713)
);

OAI22xp5_ASAP7_75t_L g2714 ( 
.A1(n_2657),
.A2(n_207),
.B1(n_204),
.B2(n_206),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2590),
.Y(n_2715)
);

OAI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2630),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_2716)
);

AOI22xp33_ASAP7_75t_L g2717 ( 
.A1(n_2646),
.A2(n_211),
.B1(n_208),
.B2(n_210),
.Y(n_2717)
);

OAI22xp5_ASAP7_75t_L g2718 ( 
.A1(n_2658),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_2718)
);

OAI221xp5_ASAP7_75t_SL g2719 ( 
.A1(n_2652),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.C(n_216),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2708),
.B(n_2635),
.Y(n_2720)
);

NAND3xp33_ASAP7_75t_L g2721 ( 
.A(n_2717),
.B(n_2639),
.C(n_2644),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2711),
.B(n_2600),
.Y(n_2722)
);

NAND4xp25_ASAP7_75t_L g2723 ( 
.A(n_2719),
.B(n_2608),
.C(n_2642),
.D(n_2620),
.Y(n_2723)
);

AOI21xp5_ASAP7_75t_L g2724 ( 
.A1(n_2684),
.A2(n_2645),
.B(n_2653),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2672),
.B(n_2643),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2683),
.B(n_2650),
.Y(n_2726)
);

AND2x2_ASAP7_75t_SL g2727 ( 
.A(n_2717),
.B(n_2651),
.Y(n_2727)
);

NAND3xp33_ASAP7_75t_L g2728 ( 
.A(n_2689),
.B(n_2660),
.C(n_2656),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_2695),
.B(n_2623),
.Y(n_2729)
);

OAI21xp5_ASAP7_75t_SL g2730 ( 
.A1(n_2670),
.A2(n_2655),
.B(n_2627),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_2715),
.B(n_2641),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2662),
.A2(n_2635),
.B1(n_2647),
.B2(n_2610),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2712),
.A2(n_2647),
.B1(n_2624),
.B2(n_2615),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2686),
.B(n_2580),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2685),
.B(n_2591),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2693),
.B(n_2591),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2662),
.B(n_2591),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2703),
.B(n_214),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2665),
.B(n_2664),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2665),
.B(n_216),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2664),
.B(n_217),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2707),
.B(n_217),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2676),
.B(n_218),
.Y(n_2743)
);

OAI21xp5_ASAP7_75t_SL g2744 ( 
.A1(n_2714),
.A2(n_219),
.B(n_221),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2663),
.B(n_2666),
.Y(n_2745)
);

OAI22xp5_ASAP7_75t_L g2746 ( 
.A1(n_2713),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_2746)
);

OA21x2_ASAP7_75t_L g2747 ( 
.A1(n_2692),
.A2(n_2694),
.B(n_2696),
.Y(n_2747)
);

AOI22xp33_ASAP7_75t_L g2748 ( 
.A1(n_2669),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_L g2749 ( 
.A(n_2666),
.B(n_224),
.Y(n_2749)
);

NAND2xp33_ASAP7_75t_L g2750 ( 
.A(n_2681),
.B(n_225),
.Y(n_2750)
);

AND2x2_ASAP7_75t_L g2751 ( 
.A(n_2706),
.B(n_225),
.Y(n_2751)
);

NAND3xp33_ASAP7_75t_L g2752 ( 
.A(n_2716),
.B(n_226),
.C(n_230),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_SL g2753 ( 
.A(n_2671),
.B(n_497),
.Y(n_2753)
);

OAI221xp5_ASAP7_75t_L g2754 ( 
.A1(n_2667),
.A2(n_226),
.B1(n_231),
.B2(n_232),
.C(n_233),
.Y(n_2754)
);

OAI21xp5_ASAP7_75t_SL g2755 ( 
.A1(n_2718),
.A2(n_231),
.B(n_235),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2679),
.B(n_235),
.Y(n_2756)
);

OAI21xp33_ASAP7_75t_L g2757 ( 
.A1(n_2677),
.A2(n_2678),
.B(n_2674),
.Y(n_2757)
);

OAI21xp5_ASAP7_75t_SL g2758 ( 
.A1(n_2668),
.A2(n_237),
.B(n_239),
.Y(n_2758)
);

NAND3xp33_ASAP7_75t_L g2759 ( 
.A(n_2691),
.B(n_240),
.C(n_241),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2709),
.B(n_241),
.Y(n_2760)
);

OAI21xp5_ASAP7_75t_SL g2761 ( 
.A1(n_2702),
.A2(n_242),
.B(n_243),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2673),
.B(n_242),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_SL g2763 ( 
.A(n_2727),
.B(n_2720),
.Y(n_2763)
);

NAND3xp33_ASAP7_75t_L g2764 ( 
.A(n_2750),
.B(n_2758),
.C(n_2744),
.Y(n_2764)
);

OR2x2_ASAP7_75t_L g2765 ( 
.A(n_2722),
.B(n_2690),
.Y(n_2765)
);

NOR3xp33_ASAP7_75t_SL g2766 ( 
.A(n_2730),
.B(n_2700),
.C(n_2699),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2729),
.B(n_2705),
.Y(n_2767)
);

NAND3xp33_ASAP7_75t_L g2768 ( 
.A(n_2752),
.B(n_2698),
.C(n_2688),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_SL g2769 ( 
.A(n_2732),
.B(n_2680),
.Y(n_2769)
);

AOI22xp33_ASAP7_75t_L g2770 ( 
.A1(n_2754),
.A2(n_2675),
.B1(n_2687),
.B2(n_2682),
.Y(n_2770)
);

NAND3xp33_ASAP7_75t_L g2771 ( 
.A(n_2755),
.B(n_2701),
.C(n_2697),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2725),
.B(n_243),
.Y(n_2772)
);

OAI211xp5_ASAP7_75t_SL g2773 ( 
.A1(n_2761),
.A2(n_2710),
.B(n_2704),
.C(n_247),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2726),
.B(n_244),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_2735),
.B(n_498),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_SL g2776 ( 
.A1(n_2721),
.A2(n_2739),
.B1(n_2745),
.B2(n_2756),
.Y(n_2776)
);

OR2x2_ASAP7_75t_L g2777 ( 
.A(n_2722),
.B(n_245),
.Y(n_2777)
);

BUFx3_ASAP7_75t_L g2778 ( 
.A(n_2736),
.Y(n_2778)
);

NOR3xp33_ASAP7_75t_L g2779 ( 
.A(n_2723),
.B(n_245),
.C(n_247),
.Y(n_2779)
);

AOI22xp33_ASAP7_75t_L g2780 ( 
.A1(n_2753),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_2780)
);

AOI22xp33_ASAP7_75t_L g2781 ( 
.A1(n_2746),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_2781)
);

AND2x2_ASAP7_75t_L g2782 ( 
.A(n_2731),
.B(n_252),
.Y(n_2782)
);

NOR3xp33_ASAP7_75t_L g2783 ( 
.A(n_2746),
.B(n_252),
.C(n_253),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2738),
.B(n_2737),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_2734),
.B(n_253),
.Y(n_2785)
);

NAND4xp75_ASAP7_75t_L g2786 ( 
.A(n_2742),
.B(n_254),
.C(n_258),
.D(n_260),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2724),
.B(n_254),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2743),
.B(n_258),
.Y(n_2788)
);

OAI211xp5_ASAP7_75t_SL g2789 ( 
.A1(n_2741),
.A2(n_2740),
.B(n_2749),
.C(n_2748),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2728),
.B(n_499),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2778),
.B(n_2751),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2777),
.Y(n_2792)
);

NAND4xp75_ASAP7_75t_L g2793 ( 
.A(n_2787),
.B(n_2762),
.C(n_2760),
.D(n_2747),
.Y(n_2793)
);

NOR2x1_ASAP7_75t_L g2794 ( 
.A(n_2765),
.B(n_2747),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_2784),
.B(n_2760),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2776),
.B(n_2762),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2776),
.B(n_2757),
.Y(n_2797)
);

AND4x1_ASAP7_75t_L g2798 ( 
.A(n_2779),
.B(n_2759),
.C(n_2733),
.D(n_262),
.Y(n_2798)
);

AND2x2_ASAP7_75t_L g2799 ( 
.A(n_2767),
.B(n_260),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2782),
.B(n_261),
.Y(n_2800)
);

INVx4_ASAP7_75t_L g2801 ( 
.A(n_2786),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2772),
.Y(n_2802)
);

HB1xp67_ASAP7_75t_L g2803 ( 
.A(n_2785),
.Y(n_2803)
);

OAI22x1_ASAP7_75t_L g2804 ( 
.A1(n_2798),
.A2(n_2763),
.B1(n_2764),
.B2(n_2769),
.Y(n_2804)
);

HB1xp67_ASAP7_75t_L g2805 ( 
.A(n_2792),
.Y(n_2805)
);

OR2x2_ASAP7_75t_L g2806 ( 
.A(n_2795),
.B(n_2803),
.Y(n_2806)
);

INVxp67_ASAP7_75t_L g2807 ( 
.A(n_2794),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2802),
.Y(n_2808)
);

INVx2_ASAP7_75t_SL g2809 ( 
.A(n_2791),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2796),
.Y(n_2810)
);

XNOR2xp5_ASAP7_75t_L g2811 ( 
.A(n_2798),
.B(n_2788),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2793),
.Y(n_2812)
);

OA22x2_ASAP7_75t_L g2813 ( 
.A1(n_2804),
.A2(n_2801),
.B1(n_2797),
.B2(n_2799),
.Y(n_2813)
);

INVxp33_ASAP7_75t_L g2814 ( 
.A(n_2811),
.Y(n_2814)
);

AOI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2812),
.A2(n_2801),
.B1(n_2783),
.B2(n_2790),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2808),
.Y(n_2816)
);

INVx2_ASAP7_75t_SL g2817 ( 
.A(n_2805),
.Y(n_2817)
);

OAI22xp5_ASAP7_75t_L g2818 ( 
.A1(n_2810),
.A2(n_2771),
.B1(n_2766),
.B2(n_2781),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2806),
.Y(n_2819)
);

OA22x2_ASAP7_75t_L g2820 ( 
.A1(n_2807),
.A2(n_2774),
.B1(n_2775),
.B2(n_2800),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2816),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2819),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2817),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2820),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2818),
.Y(n_2825)
);

HB1xp67_ASAP7_75t_L g2826 ( 
.A(n_2813),
.Y(n_2826)
);

INVxp67_ASAP7_75t_L g2827 ( 
.A(n_2826),
.Y(n_2827)
);

INVx2_ASAP7_75t_L g2828 ( 
.A(n_2823),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2821),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2828),
.Y(n_2830)
);

OAI22xp5_ASAP7_75t_L g2831 ( 
.A1(n_2827),
.A2(n_2825),
.B1(n_2815),
.B2(n_2807),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2829),
.Y(n_2832)
);

O2A1O1Ixp33_ASAP7_75t_SL g2833 ( 
.A1(n_2827),
.A2(n_2814),
.B(n_2824),
.C(n_2822),
.Y(n_2833)
);

OA22x2_ASAP7_75t_L g2834 ( 
.A1(n_2831),
.A2(n_2809),
.B1(n_2773),
.B2(n_2789),
.Y(n_2834)
);

AOI221xp5_ASAP7_75t_L g2835 ( 
.A1(n_2833),
.A2(n_2773),
.B1(n_2789),
.B2(n_2780),
.C(n_2768),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2830),
.B(n_2770),
.Y(n_2836)
);

AOI22xp5_ASAP7_75t_L g2837 ( 
.A1(n_2832),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_2837)
);

AOI22xp5_ASAP7_75t_L g2838 ( 
.A1(n_2831),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_2838)
);

AOI221xp5_ASAP7_75t_L g2839 ( 
.A1(n_2833),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.C(n_270),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2836),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2839),
.A2(n_266),
.B1(n_268),
.B2(n_270),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2837),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2834),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2838),
.B(n_273),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2835),
.B(n_273),
.Y(n_2845)
);

AOI22xp5_ASAP7_75t_SL g2846 ( 
.A1(n_2845),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_2846)
);

AOI22x1_ASAP7_75t_L g2847 ( 
.A1(n_2843),
.A2(n_276),
.B1(n_278),
.B2(n_280),
.Y(n_2847)
);

AO22x2_ASAP7_75t_L g2848 ( 
.A1(n_2842),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_2848)
);

NOR2x1_ASAP7_75t_L g2849 ( 
.A(n_2844),
.B(n_281),
.Y(n_2849)
);

OAI22x1_ASAP7_75t_L g2850 ( 
.A1(n_2841),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2847),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_2848),
.Y(n_2852)
);

AND2x2_ASAP7_75t_SL g2853 ( 
.A(n_2846),
.B(n_2840),
.Y(n_2853)
);

HB1xp67_ASAP7_75t_L g2854 ( 
.A(n_2849),
.Y(n_2854)
);

INVx1_ASAP7_75t_L g2855 ( 
.A(n_2850),
.Y(n_2855)
);

AOI22xp33_ASAP7_75t_SL g2856 ( 
.A1(n_2853),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_2856)
);

AOI211xp5_ASAP7_75t_SL g2857 ( 
.A1(n_2854),
.A2(n_285),
.B(n_286),
.C(n_287),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2855),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2851),
.Y(n_2859)
);

INVxp67_ASAP7_75t_L g2860 ( 
.A(n_2852),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2858),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2860),
.Y(n_2862)
);

INVx1_ASAP7_75t_SL g2863 ( 
.A(n_2856),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2859),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2857),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2862),
.A2(n_286),
.B1(n_288),
.B2(n_289),
.Y(n_2866)
);

INVx2_ASAP7_75t_L g2867 ( 
.A(n_2866),
.Y(n_2867)
);

OAI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2867),
.A2(n_2865),
.B1(n_2863),
.B2(n_2861),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2868),
.Y(n_2869)
);

AOI221xp5_ASAP7_75t_L g2870 ( 
.A1(n_2869),
.A2(n_2864),
.B1(n_291),
.B2(n_292),
.C(n_293),
.Y(n_2870)
);

AOI211xp5_ASAP7_75t_L g2871 ( 
.A1(n_2870),
.A2(n_288),
.B(n_293),
.C(n_294),
.Y(n_2871)
);


endmodule