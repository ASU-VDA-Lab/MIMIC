module fake_jpeg_10774_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_13),
.B(n_0),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_41),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_28),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_42),
.B(n_71),
.C(n_8),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_43),
.B(n_56),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_18),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_58),
.Y(n_82)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_14),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_57),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_0),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_59),
.B(n_61),
.Y(n_85)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_0),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_66),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_64),
.Y(n_102)
);

INVx5_ASAP7_75t_SL g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_65),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_2),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_67),
.Y(n_103)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_19),
.B(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_72),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_6),
.B(n_7),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_24),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_75),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_6),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_24),
.B1(n_15),
.B2(n_37),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_79),
.A2(n_88),
.B1(n_92),
.B2(n_106),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_111),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_40),
.A2(n_54),
.B1(n_67),
.B2(n_47),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_35),
.B1(n_37),
.B2(n_23),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_90),
.A2(n_78),
.B1(n_77),
.B2(n_84),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_35),
.B1(n_23),
.B2(n_31),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_97),
.B(n_105),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_65),
.B(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_100),
.B(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_44),
.B(n_30),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_31),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_45),
.A2(n_26),
.B1(n_10),
.B2(n_11),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_69),
.A2(n_26),
.B1(n_11),
.B2(n_12),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_68),
.B1(n_12),
.B2(n_11),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_49),
.B(n_8),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_108),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_8),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_63),
.A2(n_52),
.B1(n_57),
.B2(n_55),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_88),
.B1(n_92),
.B2(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_117),
.A2(n_121),
.B1(n_124),
.B2(n_139),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_118),
.B(n_136),
.Y(n_180)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_53),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_125),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_72),
.B1(n_60),
.B2(n_41),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_85),
.B(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_26),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_141),
.Y(n_161)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_91),
.A2(n_95),
.B(n_86),
.C(n_98),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_137),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_114),
.Y(n_129)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_83),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_135),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_109),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_96),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_78),
.A2(n_103),
.B1(n_77),
.B2(n_84),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_143),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_149),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_150),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_99),
.B(n_76),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_93),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_122),
.Y(n_177)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_153),
.Y(n_172)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_133),
.B(n_123),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_117),
.B1(n_149),
.B2(n_118),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_133),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_169),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_121),
.C(n_136),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_173),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_143),
.B1(n_145),
.B2(n_128),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_132),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_144),
.B(n_134),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_146),
.Y(n_198)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_167),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_183),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_140),
.Y(n_183)
);

AND2x4_ASAP7_75t_SL g185 ( 
.A(n_170),
.B(n_176),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_185),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_165),
.B(n_151),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_191),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_168),
.A2(n_138),
.B(n_153),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_195),
.B(n_196),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_192),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_157),
.A2(n_139),
.B1(n_119),
.B2(n_152),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_160),
.B1(n_156),
.B2(n_180),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_135),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_170),
.B(n_157),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_162),
.C(n_166),
.Y(n_210)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_175),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_204),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_209),
.B1(n_214),
.B2(n_184),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_193),
.Y(n_207)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_207),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_156),
.B1(n_160),
.B2(n_161),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_213),
.C(n_189),
.Y(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_211),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_154),
.C(n_159),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_160),
.B1(n_171),
.B2(n_175),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_223),
.C(n_213),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_SL g216 ( 
.A1(n_201),
.A2(n_188),
.B(n_194),
.C(n_185),
.Y(n_216)
);

OAI31xp33_ASAP7_75t_L g227 ( 
.A1(n_216),
.A2(n_206),
.A3(n_212),
.B(n_214),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_203),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_183),
.C(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_203),
.Y(n_231)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_181),
.B(n_187),
.C(n_185),
.D(n_195),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_222),
.A2(n_225),
.B(n_202),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_181),
.C(n_192),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_184),
.B(n_185),
.Y(n_225)
);

AOI31xp67_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_229),
.A3(n_230),
.B(n_220),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_227),
.A2(n_228),
.B(n_216),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_202),
.B(n_206),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_219),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_219),
.B(n_204),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_232),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_227),
.Y(n_239)
);

AOI31xp67_ASAP7_75t_SL g241 ( 
.A1(n_234),
.A2(n_235),
.A3(n_185),
.B(n_198),
.Y(n_241)
);

AOI31xp67_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_225),
.A3(n_222),
.B(n_216),
.Y(n_235)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_236),
.A2(n_211),
.B(n_191),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_228),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_239),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_221),
.C(n_224),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_190),
.B1(n_200),
.B2(n_158),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_179),
.B(n_131),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_166),
.Y(n_247)
);

OAI221xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_211),
.B1(n_200),
.B2(n_199),
.C(n_171),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_240),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_248),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_250),
.A2(n_246),
.B(n_249),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_251),
.A2(n_179),
.B1(n_158),
.B2(n_174),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_174),
.Y(n_253)
);


endmodule