module fake_jpeg_18806_n_67 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_67);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_67;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_5),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_9),
.B(n_1),
.Y(n_24)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_22),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_35),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_26),
.A2(n_2),
.B(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_13),
.B1(n_18),
.B2(n_10),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_10),
.B(n_34),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_33),
.C(n_37),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_51),
.C(n_52),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_16),
.C(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_53),
.B(n_47),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_55),
.A2(n_43),
.B(n_49),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_50),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_49),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_55),
.A2(n_43),
.B(n_46),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_58),
.A2(n_60),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_59),
.B(n_54),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NOR3xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_40),
.C(n_41),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_40),
.C(n_41),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_63),
.A3(n_41),
.B1(n_21),
.B2(n_8),
.C1(n_7),
.C2(n_5),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_21),
.C(n_8),
.Y(n_67)
);


endmodule