module fake_ariane_2829_n_106 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_106);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_106;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp33_ASAP7_75t_SL g20 ( 
.A(n_18),
.Y(n_20)
);

INVxp67_ASAP7_75t_SL g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx2_ASAP7_75t_SL g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_28),
.Y(n_50)
);

NOR2xp67_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_17),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_20),
.B1(n_21),
.B2(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_55),
.Y(n_57)
);

NOR3xp33_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_39),
.C(n_23),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

OAI21x1_ASAP7_75t_L g61 ( 
.A1(n_51),
.A2(n_37),
.B(n_35),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_53),
.Y(n_63)
);

AOI21x1_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_37),
.B(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_62),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_65),
.A2(n_52),
.B1(n_42),
.B2(n_60),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

AO31x2_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_47),
.A3(n_38),
.B(n_30),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_36),
.B(n_60),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_49),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_63),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_63),
.B(n_73),
.C(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_71),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_75),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_71),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_71),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_84),
.Y(n_87)
);

OAI321xp33_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_38),
.A3(n_67),
.B1(n_62),
.B2(n_64),
.C(n_26),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_62),
.B1(n_71),
.B2(n_4),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_85),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_82),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_82),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_85),
.C(n_86),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_83),
.C(n_2),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_93),
.B(n_1),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_95),
.B(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_100),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_102),
.Y(n_103)
);

OAI322xp33_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_99),
.A3(n_97),
.B1(n_4),
.B2(n_5),
.C1(n_26),
.C2(n_9),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_60),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_13),
.B(n_15),
.Y(n_106)
);


endmodule