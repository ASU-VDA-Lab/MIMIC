module fake_jpeg_12423_n_620 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_620);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_620;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_SL g51 ( 
.A(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_13),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_61),
.Y(n_168)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_62),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_63),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_64),
.Y(n_182)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_20),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_67),
.B(n_74),
.Y(n_134)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_51),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g192 ( 
.A(n_69),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_70),
.Y(n_188)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g158 ( 
.A(n_72),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_73),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_39),
.B(n_11),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_10),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_78),
.B(n_89),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_79),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_33),
.B(n_18),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_96),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_85),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_54),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_86),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_87),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_10),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_93),
.B(n_94),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_42),
.B(n_10),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_33),
.B(n_9),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_103),
.Y(n_162)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_43),
.Y(n_104)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_28),
.Y(n_106)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_106),
.Y(n_208)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_42),
.B(n_9),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_123),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_28),
.Y(n_112)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_23),
.Y(n_113)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_37),
.Y(n_114)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_23),
.Y(n_115)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_115),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_59),
.Y(n_120)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_120),
.Y(n_174)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_27),
.Y(n_122)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_27),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_27),
.Y(n_124)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_43),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_125),
.A2(n_34),
.B(n_56),
.Y(n_163)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_126),
.B(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_34),
.B(n_12),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_37),
.B1(n_32),
.B2(n_29),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_140),
.A2(n_154),
.B1(n_161),
.B2(n_172),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g147 ( 
.A1(n_68),
.A2(n_29),
.B1(n_32),
.B2(n_44),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g261 ( 
.A1(n_147),
.A2(n_193),
.B(n_165),
.C(n_134),
.Y(n_261)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_67),
.B(n_25),
.CON(n_150),
.SN(n_150)
);

OAI21xp33_ASAP7_75t_L g274 ( 
.A1(n_150),
.A2(n_193),
.B(n_0),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_30),
.C(n_52),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_152),
.B(n_190),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_60),
.A2(n_56),
.B1(n_45),
.B2(n_44),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_87),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_156),
.B(n_175),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_61),
.A2(n_40),
.B1(n_57),
.B2(n_52),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_163),
.B(n_47),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_74),
.A2(n_45),
.B1(n_36),
.B2(n_57),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_167),
.A2(n_187),
.B1(n_88),
.B2(n_85),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_63),
.A2(n_40),
.B1(n_50),
.B2(n_24),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_78),
.B(n_36),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_94),
.B(n_50),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_177),
.B(n_184),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_110),
.B(n_25),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_178),
.B(n_183),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_121),
.B(n_46),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_105),
.B(n_46),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_64),
.A2(n_38),
.B1(n_30),
.B2(n_24),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_72),
.Y(n_190)
);

HAxp5_ASAP7_75t_SL g193 ( 
.A(n_104),
.B(n_49),
.CON(n_193),
.SN(n_193)
);

AO22x2_ASAP7_75t_L g194 ( 
.A1(n_70),
.A2(n_38),
.B1(n_22),
.B2(n_49),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_194),
.A2(n_124),
.B1(n_119),
.B2(n_116),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_99),
.A2(n_49),
.B1(n_47),
.B2(n_22),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_198),
.A2(n_122),
.B1(n_115),
.B2(n_113),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_100),
.A2(n_49),
.B1(n_47),
.B2(n_3),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_199),
.A2(n_13),
.B1(n_15),
.B2(n_5),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_SL g202 ( 
.A(n_69),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_112),
.B(n_109),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_204),
.B(n_6),
.Y(n_262)
);

BUFx16f_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_213),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_214),
.A2(n_242),
.B1(n_255),
.B2(n_258),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_143),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_216),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_143),
.Y(n_218)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_218),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_161),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_220),
.B(n_235),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_221),
.Y(n_325)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_222),
.Y(n_316)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_223),
.Y(n_317)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_224),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_147),
.A2(n_86),
.B1(n_75),
.B2(n_79),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_225),
.A2(n_248),
.B1(n_259),
.B2(n_158),
.Y(n_310)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_226),
.Y(n_299)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_151),
.Y(n_227)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_227),
.Y(n_328)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_228),
.Y(n_305)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_168),
.Y(n_229)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_229),
.Y(n_334)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_137),
.Y(n_230)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_230),
.Y(n_300)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_139),
.Y(n_231)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_231),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_148),
.B(n_49),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_232),
.Y(n_326)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_130),
.Y(n_233)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_233),
.Y(n_337)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_142),
.Y(n_236)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_236),
.Y(n_303)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_155),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_237),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_238),
.A2(n_260),
.B1(n_188),
.B2(n_200),
.Y(n_335)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_239),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_180),
.Y(n_240)
);

INVx8_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_241),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_146),
.A2(n_73),
.B1(n_98),
.B2(n_95),
.Y(n_242)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_180),
.Y(n_243)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_243),
.Y(n_320)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_186),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_246),
.Y(n_294)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_245),
.B(n_251),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_157),
.B(n_47),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_254),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_194),
.A2(n_111),
.B1(n_47),
.B2(n_91),
.Y(n_248)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

BUFx8_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

INVx4_ASAP7_75t_SL g291 ( 
.A(n_250),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_198),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_252),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_169),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_147),
.A2(n_8),
.B1(n_16),
.B2(n_3),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_140),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_256),
.B(n_262),
.Y(n_304)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_257),
.B(n_261),
.Y(n_315)
);

OAI22xp33_ASAP7_75t_L g258 ( 
.A1(n_194),
.A2(n_8),
.B1(n_15),
.B2(n_3),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_205),
.A2(n_6),
.B1(n_15),
.B2(n_3),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_176),
.A2(n_6),
.B1(n_13),
.B2(n_14),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_263),
.A2(n_264),
.B1(n_270),
.B2(n_271),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_150),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_141),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_265),
.B(n_266),
.Y(n_308)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_182),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_174),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_267),
.B(n_272),
.Y(n_314)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_268),
.B(n_269),
.Y(n_333)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_197),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_203),
.A2(n_0),
.B1(n_1),
.B2(n_201),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_188),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_133),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_159),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_275),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_274),
.A2(n_281),
.B1(n_158),
.B2(n_203),
.Y(n_319)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_181),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_145),
.B(n_0),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_276),
.B(n_129),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_197),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_279),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_164),
.A2(n_0),
.B1(n_1),
.B2(n_173),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_278),
.A2(n_209),
.B(n_165),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_153),
.B(n_0),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_208),
.B(n_1),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_280),
.B(n_209),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_128),
.A2(n_1),
.B1(n_131),
.B2(n_210),
.Y(n_281)
);

AND2x4_ASAP7_75t_SL g282 ( 
.A(n_162),
.B(n_144),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_136),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_282),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_287),
.B(n_298),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_289),
.B(n_310),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_296),
.B(n_339),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_282),
.Y(n_298)
);

CKINVDCx12_ASAP7_75t_R g301 ( 
.A(n_234),
.Y(n_301)
);

BUFx4f_ASAP7_75t_SL g369 ( 
.A(n_301),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_238),
.A2(n_210),
.B1(n_205),
.B2(n_189),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_311),
.A2(n_327),
.B1(n_335),
.B2(n_310),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_251),
.B(n_211),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_321),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_319),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_207),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_252),
.A2(n_133),
.B1(n_160),
.B2(n_132),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_322),
.A2(n_331),
.B1(n_215),
.B2(n_243),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_248),
.A2(n_189),
.B1(n_185),
.B2(n_191),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_214),
.A2(n_132),
.B1(n_129),
.B2(n_135),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_185),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_332),
.B(n_250),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_338),
.A2(n_278),
.B(n_260),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_191),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_340),
.B(n_218),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_292),
.A2(n_242),
.B1(n_281),
.B2(n_219),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_343),
.A2(n_355),
.B1(n_364),
.B2(n_372),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_351),
.B(n_352),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_308),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_345),
.B(n_349),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_288),
.B(n_212),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_346),
.B(n_378),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_288),
.B(n_253),
.C(n_222),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_361),
.C(n_374),
.Y(n_386)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_348),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_318),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_315),
.A2(n_274),
.B(n_261),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_315),
.A2(n_258),
.B(n_239),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_323),
.A2(n_200),
.B1(n_229),
.B2(n_266),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_353),
.A2(n_362),
.B1(n_366),
.B2(n_327),
.Y(n_396)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_315),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_370),
.Y(n_405)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_357),
.Y(n_399)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_306),
.Y(n_358)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_358),
.Y(n_409)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_359),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_288),
.B(n_224),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_323),
.A2(n_287),
.B1(n_298),
.B2(n_304),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_317),
.B(n_228),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_363),
.B(n_377),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_311),
.A2(n_275),
.B1(n_245),
.B2(n_249),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_312),
.A2(n_240),
.B1(n_271),
.B2(n_221),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_293),
.Y(n_368)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_303),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_371),
.B(n_381),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_286),
.A2(n_237),
.B1(n_241),
.B2(n_226),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_373),
.B(n_375),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_277),
.C(n_165),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_332),
.B(n_269),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_313),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_376),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_268),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_296),
.B(n_272),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_286),
.A2(n_233),
.B1(n_257),
.B2(n_216),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_379),
.A2(n_333),
.B(n_307),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_314),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_380),
.B(n_290),
.Y(n_410)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_382),
.B(n_291),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_324),
.B(n_215),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_301),
.Y(n_404)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_313),
.Y(n_384)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_384),
.Y(n_387)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_385),
.B(n_316),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_294),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_403),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_351),
.A2(n_338),
.B(n_285),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_392),
.A2(n_394),
.B(n_395),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_342),
.A2(n_289),
.B(n_295),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_354),
.A2(n_326),
.B(n_297),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_406),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_326),
.B1(n_320),
.B2(n_337),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_398),
.A2(n_412),
.B1(n_420),
.B2(n_384),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_355),
.A2(n_320),
.B1(n_302),
.B2(n_334),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_402),
.A2(n_370),
.B1(n_381),
.B2(n_371),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_342),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_404),
.B(n_377),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_373),
.B(n_302),
.Y(n_406)
);

AND2x2_ASAP7_75t_SL g407 ( 
.A(n_361),
.B(n_309),
.Y(n_407)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_407),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_410),
.B(n_418),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_367),
.A2(n_337),
.B1(n_334),
.B2(n_330),
.Y(n_412)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_362),
.B(n_378),
.C(n_350),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_413),
.A2(n_383),
.B(n_354),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_415),
.B(n_385),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_350),
.B(n_375),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_369),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_349),
.B(n_309),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_419),
.A2(n_366),
.B1(n_368),
.B2(n_344),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_367),
.A2(n_330),
.B1(n_325),
.B2(n_293),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_421),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_400),
.Y(n_460)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_389),
.Y(n_424)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_396),
.A2(n_345),
.B1(n_353),
.B2(n_364),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_425),
.A2(n_434),
.B1(n_439),
.B2(n_440),
.Y(n_479)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_428),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_431),
.A2(n_454),
.B(n_419),
.Y(n_475)
);

CKINVDCx14_ASAP7_75t_R g476 ( 
.A(n_432),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_433),
.A2(n_448),
.B1(n_399),
.B2(n_422),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_421),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_435),
.B(n_395),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_391),
.A2(n_380),
.B(n_374),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_437),
.Y(n_478)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_409),
.Y(n_438)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_438),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_360),
.B1(n_382),
.B2(n_352),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_393),
.A2(n_360),
.B1(n_363),
.B2(n_359),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_409),
.Y(n_441)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_391),
.A2(n_368),
.B1(n_348),
.B2(n_357),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_447),
.Y(n_463)
);

OAI21xp33_ASAP7_75t_L g443 ( 
.A1(n_404),
.A2(n_369),
.B(n_333),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_443),
.B(n_445),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_416),
.B(n_333),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_414),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_446),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_394),
.A2(n_293),
.B1(n_325),
.B2(n_307),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_393),
.A2(n_325),
.B1(n_307),
.B2(n_290),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_390),
.A2(n_305),
.B1(n_341),
.B2(n_316),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_449),
.A2(n_420),
.B1(n_399),
.B2(n_422),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_397),
.B(n_305),
.Y(n_452)
);

XOR2x1_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_453),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_397),
.B(n_328),
.Y(n_453)
);

OAI21x1_ASAP7_75t_R g454 ( 
.A1(n_414),
.A2(n_405),
.B(n_417),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_407),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_450),
.B(n_405),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_458),
.B(n_464),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_386),
.C(n_403),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_470),
.C(n_488),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_460),
.B(n_473),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_461),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_435),
.B(n_408),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_456),
.A2(n_392),
.B(n_407),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_469),
.A2(n_475),
.B(n_487),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_386),
.C(n_455),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_472),
.A2(n_480),
.B1(n_481),
.B2(n_482),
.Y(n_490)
);

XNOR2x1_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_400),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_474),
.B(n_433),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_427),
.A2(n_401),
.B1(n_413),
.B2(n_390),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_427),
.A2(n_413),
.B1(n_402),
.B2(n_408),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_426),
.B(n_388),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_483),
.B(n_484),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_426),
.B(n_341),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_456),
.A2(n_407),
.B(n_415),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_411),
.C(n_328),
.Y(n_488)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_485),
.Y(n_491)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_491),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_493),
.Y(n_538)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g495 ( 
.A1(n_475),
.A2(n_429),
.B(n_431),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_495),
.B(n_498),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_466),
.Y(n_496)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_496),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_481),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_464),
.B(n_452),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_500),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_479),
.A2(n_444),
.B1(n_428),
.B2(n_424),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_501),
.A2(n_463),
.B1(n_467),
.B2(n_478),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_458),
.B(n_432),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_504),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_465),
.A2(n_429),
.B(n_423),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_479),
.Y(n_505)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_459),
.B(n_429),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_512),
.Y(n_519)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_486),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_507),
.A2(n_509),
.B1(n_511),
.B2(n_515),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_470),
.B(n_445),
.C(n_439),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_508),
.B(n_460),
.C(n_474),
.Y(n_521)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_480),
.A2(n_425),
.B1(n_434),
.B2(n_444),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_510),
.A2(n_478),
.B1(n_463),
.B2(n_468),
.Y(n_518)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_465),
.A2(n_442),
.B(n_437),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_468),
.B(n_430),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_482),
.Y(n_524)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_462),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_488),
.B(n_453),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_516),
.B(n_517),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_518),
.A2(n_496),
.B1(n_515),
.B2(n_511),
.Y(n_553)
);

MAJx2_ASAP7_75t_L g560 ( 
.A(n_521),
.B(n_495),
.C(n_457),
.Y(n_560)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_524),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_506),
.B(n_473),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_525),
.B(n_527),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_514),
.B(n_471),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_502),
.B(n_487),
.C(n_469),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_528),
.B(n_535),
.C(n_539),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_502),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_529),
.B(n_532),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_531),
.A2(n_533),
.B1(n_540),
.B2(n_510),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_471),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_501),
.A2(n_476),
.B1(n_467),
.B2(n_477),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_508),
.B(n_466),
.C(n_447),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_504),
.B(n_438),
.C(n_446),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_498),
.A2(n_472),
.B1(n_457),
.B2(n_448),
.Y(n_540)
);

CKINVDCx14_ASAP7_75t_R g543 ( 
.A(n_536),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_552),
.Y(n_567)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_541),
.Y(n_544)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_544),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_534),
.B(n_489),
.Y(n_546)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_546),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_490),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_SL g576 ( 
.A(n_547),
.B(n_548),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_529),
.B(n_492),
.C(n_490),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_549),
.A2(n_559),
.B1(n_537),
.B2(n_524),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_528),
.B(n_525),
.C(n_539),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_551),
.C(n_519),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_521),
.B(n_492),
.C(n_512),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_533),
.Y(n_552)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_553),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_531),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_556),
.B(n_557),
.Y(n_578)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_538),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_530),
.B(n_513),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_558),
.Y(n_566)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_523),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_561),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_518),
.B(n_526),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_SL g563 ( 
.A(n_554),
.B(n_519),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_563),
.B(n_520),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_553),
.A2(n_522),
.B(n_497),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_565),
.A2(n_558),
.B(n_542),
.Y(n_587)
);

XOR2x1_ASAP7_75t_SL g568 ( 
.A(n_549),
.B(n_527),
.Y(n_568)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_568),
.B(n_570),
.Y(n_582)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_551),
.A2(n_497),
.B(n_540),
.Y(n_570)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_571),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_572),
.B(n_573),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_545),
.B(n_550),
.C(n_547),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_545),
.B(n_548),
.C(n_555),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_575),
.B(n_577),
.C(n_554),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_555),
.B(n_520),
.C(n_532),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_573),
.B(n_499),
.Y(n_580)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_580),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_569),
.B(n_557),
.Y(n_581)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_581),
.Y(n_596)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_565),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_583),
.A2(n_574),
.B1(n_566),
.B2(n_577),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_563),
.C(n_564),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g592 ( 
.A(n_585),
.B(n_588),
.Y(n_592)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_572),
.B(n_542),
.C(n_561),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_586),
.A2(n_587),
.B(n_590),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_562),
.A2(n_493),
.B1(n_509),
.B2(n_507),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_575),
.B(n_560),
.C(n_494),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_567),
.B(n_491),
.Y(n_591)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_591),
.B(n_570),
.Y(n_595)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_594),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_595),
.B(n_597),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_590),
.A2(n_568),
.B1(n_576),
.B2(n_564),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_598),
.B(n_600),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_578),
.B(n_571),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_599),
.A2(n_582),
.B(n_587),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_589),
.B(n_441),
.C(n_417),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_593),
.B(n_586),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_603),
.B(n_604),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g605 ( 
.A1(n_596),
.A2(n_579),
.B1(n_585),
.B2(n_584),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_605),
.B(n_607),
.C(n_595),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_601),
.B(n_588),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_609),
.A2(n_612),
.B(n_603),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_608),
.B(n_592),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_602),
.C(n_387),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_606),
.B(n_600),
.C(n_592),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_613),
.A2(n_614),
.B(n_610),
.Y(n_615)
);

AOI322xp5_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_454),
.A3(n_369),
.B1(n_336),
.B2(n_387),
.C1(n_449),
.C2(n_291),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_SL g617 ( 
.A1(n_616),
.A2(n_369),
.B(n_291),
.Y(n_617)
);

AOI321xp33_ASAP7_75t_L g618 ( 
.A1(n_617),
.A2(n_213),
.A3(n_329),
.B1(n_336),
.B2(n_454),
.C(n_369),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_618),
.B(n_213),
.Y(n_619)
);

OAI311xp33_ASAP7_75t_L g620 ( 
.A1(n_619),
.A2(n_329),
.A3(n_336),
.B1(n_454),
.C1(n_369),
.Y(n_620)
);


endmodule