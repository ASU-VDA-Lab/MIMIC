module fake_jpeg_17050_n_122 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_2),
.B(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_28),
.B(n_40),
.Y(n_52)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_33),
.B(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_18),
.A2(n_13),
.B1(n_20),
.B2(n_19),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_41),
.B1(n_19),
.B2(n_20),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_3),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_44),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_4),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_13),
.B1(n_23),
.B2(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_49),
.B1(n_50),
.B2(n_65),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_17),
.B1(n_4),
.B2(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_51),
.B(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_27),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_58),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_26),
.C(n_24),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_62),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_4),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_15),
.B1(n_25),
.B2(n_11),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_5),
.C(n_7),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_29),
.C(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_R g69 ( 
.A(n_52),
.B(n_43),
.Y(n_69)
);

NOR2xp67_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_57),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_76),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_72),
.B(n_80),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_58),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_52),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_87),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_62),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_61),
.B(n_47),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_90),
.B(n_95),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_77),
.C(n_82),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_75),
.A2(n_50),
.B1(n_56),
.B2(n_66),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_92),
.A2(n_81),
.B1(n_73),
.B2(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_106),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_72),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_100),
.B(n_102),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_73),
.C(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_103),
.B(n_104),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_74),
.C(n_85),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_64),
.B(n_90),
.Y(n_106)
);

AOI221xp5_ASAP7_75t_L g110 ( 
.A1(n_101),
.A2(n_90),
.B1(n_86),
.B2(n_88),
.C(n_93),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_110),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_98),
.C(n_103),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_115),
.C(n_108),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_104),
.C(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_116),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_119),
.Y(n_122)
);


endmodule