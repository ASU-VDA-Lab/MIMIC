module fake_jpeg_3039_n_563 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_563);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_563;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_SL g45 ( 
.A(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_57),
.Y(n_161)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_59),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_60),
.B(n_64),
.Y(n_130)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_62),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_20),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_68),
.B(n_71),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_69),
.Y(n_182)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_18),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_72),
.B(n_82),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_73),
.Y(n_212)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_14),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_76),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_55),
.B(n_17),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_78),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_14),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_120),
.Y(n_146)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_81),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g165 ( 
.A(n_84),
.Y(n_165)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_85),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_28),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_91),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_28),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_92),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_23),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_93),
.B(n_94),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_23),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_34),
.Y(n_95)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_97),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_30),
.Y(n_99)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_100),
.Y(n_205)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_102),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_103),
.Y(n_164)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_45),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_111),
.Y(n_178)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_106),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

CKINVDCx6p67_ASAP7_75t_R g189 ( 
.A(n_107),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_19),
.Y(n_110)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_45),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_112),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_19),
.Y(n_113)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_113),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_19),
.Y(n_114)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_115),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_30),
.B(n_17),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_116),
.B(n_0),
.Y(n_190)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_45),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_33),
.B(n_13),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_44),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_22),
.Y(n_127)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_22),
.Y(n_122)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_122),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_33),
.B(n_0),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_41),
.Y(n_163)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_36),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_124),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_125),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_127),
.B(n_188),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_54),
.B1(n_46),
.B2(n_50),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_132),
.A2(n_135),
.B1(n_139),
.B2(n_175),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_84),
.A2(n_87),
.B1(n_56),
.B2(n_88),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_54),
.B1(n_50),
.B2(n_22),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_52),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_140),
.B(n_158),
.Y(n_223)
);

INVx6_ASAP7_75t_SL g142 ( 
.A(n_107),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_142),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_38),
.B1(n_52),
.B2(n_37),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_144),
.A2(n_179),
.B(n_198),
.C(n_203),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_59),
.A2(n_37),
.B(n_21),
.C(n_38),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_145),
.A2(n_190),
.B(n_213),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_62),
.B(n_41),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_163),
.B(n_192),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_96),
.A2(n_21),
.B1(n_22),
.B2(n_51),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_171),
.A2(n_185),
.B1(n_179),
.B2(n_208),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_100),
.A2(n_51),
.B1(n_53),
.B2(n_36),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_51),
.B1(n_48),
.B2(n_35),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_73),
.A2(n_78),
.B1(n_81),
.B2(n_57),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_180),
.A2(n_181),
.B1(n_197),
.B2(n_201),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_63),
.A2(n_48),
.B1(n_35),
.B2(n_53),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_69),
.A2(n_53),
.B1(n_48),
.B2(n_35),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_187),
.Y(n_286)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_65),
.B(n_1),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_207),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_80),
.B(n_1),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_196),
.B(n_202),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_85),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_103),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_98),
.B(n_6),
.C(n_7),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g281 ( 
.A(n_199),
.B(n_176),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_110),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_102),
.B(n_7),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_67),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_67),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_204),
.A2(n_198),
.B1(n_203),
.B2(n_197),
.Y(n_294)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_66),
.A2(n_11),
.B1(n_12),
.B2(n_92),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_198),
.B1(n_203),
.B2(n_204),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_113),
.B(n_12),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_114),
.B(n_12),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_216),
.Y(n_243)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_119),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_140),
.B(n_108),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_219),
.B(n_230),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_177),
.A2(n_77),
.B1(n_106),
.B2(n_109),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_220),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_221),
.B(n_238),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_161),
.Y(n_224)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_224),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_184),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_184),
.Y(n_226)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_171),
.A2(n_107),
.B(n_77),
.C(n_12),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_227),
.A2(n_252),
.B(n_228),
.Y(n_308)
);

O2A1O1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_181),
.A2(n_197),
.B(n_185),
.C(n_180),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_228),
.A2(n_284),
.B(n_227),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_143),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_231),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_173),
.B(n_147),
.Y(n_232)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_232),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_234),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_235),
.B(n_252),
.Y(n_313)
);

BUFx12f_ASAP7_75t_L g236 ( 
.A(n_189),
.Y(n_236)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_236),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_154),
.Y(n_238)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_153),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_241),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_189),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_242),
.B(n_269),
.Y(n_303)
);

INVx13_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_244),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_133),
.Y(n_245)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_139),
.Y(n_246)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_174),
.B(n_141),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_247),
.B(n_248),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_138),
.B(n_146),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_134),
.B(n_169),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_249),
.B(n_255),
.Y(n_337)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_153),
.Y(n_250)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_135),
.A2(n_150),
.B1(n_186),
.B2(n_205),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_251),
.A2(n_285),
.B1(n_294),
.B2(n_296),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_SL g252 ( 
.A(n_164),
.B(n_170),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_150),
.Y(n_253)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_253),
.Y(n_318)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_155),
.B(n_211),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_172),
.B(n_218),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_256),
.B(n_257),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_178),
.B(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_191),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_258),
.B(n_262),
.Y(n_321)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_259),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_133),
.A2(n_167),
.B1(n_157),
.B2(n_152),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_260),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_162),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_261),
.B(n_266),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_126),
.B(n_167),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_165),
.Y(n_263)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_263),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_148),
.A2(n_159),
.B1(n_149),
.B2(n_168),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_237),
.B1(n_273),
.B2(n_282),
.Y(n_305)
);

OR2x2_ASAP7_75t_SL g265 ( 
.A(n_137),
.B(n_200),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g346 ( 
.A(n_265),
.B(n_276),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_156),
.B(n_149),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_128),
.Y(n_267)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_268),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_129),
.Y(n_269)
);

AND2x2_ASAP7_75t_SL g270 ( 
.A(n_151),
.B(n_136),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_270),
.B(n_275),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_148),
.B(n_159),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_271),
.B(n_279),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_136),
.B(n_194),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_274),
.B(n_292),
.Y(n_349)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_194),
.B(n_208),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_277),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_212),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_288),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_131),
.B(n_176),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_281),
.Y(n_326)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_131),
.Y(n_280)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_212),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_282),
.B(n_287),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_217),
.B(n_161),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_217),
.A2(n_175),
.B1(n_140),
.B2(n_105),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_166),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_166),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_182),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_289),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_182),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_290),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_161),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_293),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_172),
.B(n_141),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_153),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_161),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_297),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_175),
.A2(n_140),
.B1(n_105),
.B2(n_111),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_172),
.B(n_141),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_246),
.A2(n_261),
.B1(n_276),
.B2(n_281),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_302),
.A2(n_328),
.B1(n_347),
.B2(n_313),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_L g373 ( 
.A1(n_305),
.A2(n_345),
.B1(n_289),
.B2(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_308),
.Y(n_353)
);

AND2x4_ASAP7_75t_SL g309 ( 
.A(n_219),
.B(n_255),
.Y(n_309)
);

AND2x2_ASAP7_75t_SL g390 ( 
.A(n_309),
.B(n_350),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_313),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_271),
.A2(n_266),
.B1(n_223),
.B2(n_243),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_311),
.A2(n_254),
.B1(n_280),
.B2(n_250),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_248),
.A2(n_283),
.B1(n_272),
.B2(n_222),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_239),
.A2(n_284),
.B(n_265),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_334),
.A2(n_270),
.B(n_275),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_339),
.B(n_232),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_247),
.B(n_230),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_286),
.A2(n_231),
.B1(n_287),
.B2(n_263),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_239),
.A2(n_232),
.B1(n_275),
.B2(n_279),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_249),
.B(n_229),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_348),
.B(n_268),
.Y(n_368)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_351),
.Y(n_396)
);

AOI21xp33_ASAP7_75t_L g352 ( 
.A1(n_338),
.A2(n_239),
.B(n_240),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_352),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_307),
.A2(n_239),
.B1(n_236),
.B2(n_234),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_354),
.A2(n_361),
.B1(n_342),
.B2(n_325),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_355),
.B(n_366),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_320),
.B(n_337),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_356),
.B(n_358),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_332),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_377),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_320),
.B(n_286),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_359),
.A2(n_364),
.B(n_371),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g360 ( 
.A(n_304),
.Y(n_360)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_360),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g361 ( 
.A1(n_314),
.A2(n_253),
.B1(n_277),
.B2(n_245),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_306),
.B(n_233),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_372),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_326),
.B(n_270),
.C(n_293),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_363),
.B(n_374),
.C(n_382),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_346),
.A2(n_245),
.B(n_233),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_304),
.Y(n_365)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_373),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_368),
.B(n_370),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_305),
.A2(n_278),
.B1(n_290),
.B2(n_295),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_369),
.A2(n_378),
.B1(n_329),
.B2(n_325),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_337),
.B(n_241),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_338),
.A2(n_225),
.B(n_226),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_264),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_346),
.A2(n_259),
.B(n_244),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_309),
.B(n_236),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_375),
.B(n_379),
.Y(n_417)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_376),
.Y(n_427)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_331),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_334),
.A2(n_224),
.B1(n_236),
.B2(n_267),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_326),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_308),
.A2(n_347),
.B(n_310),
.Y(n_380)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_380),
.A2(n_386),
.B(n_303),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_343),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_383),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_299),
.B(n_311),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_384),
.B(n_385),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_299),
.B(n_316),
.C(n_350),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_321),
.A2(n_350),
.B(n_313),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g388 ( 
.A(n_342),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_388),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_306),
.B(n_349),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_389),
.B(n_390),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_309),
.B(n_321),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_391),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_349),
.B(n_301),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_392),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_353),
.A2(n_380),
.B1(n_372),
.B2(n_384),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_395),
.A2(n_398),
.B1(n_401),
.B2(n_405),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_353),
.A2(n_314),
.B1(n_324),
.B2(n_307),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_367),
.A2(n_391),
.B1(n_352),
.B2(n_356),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_367),
.A2(n_329),
.B1(n_319),
.B2(n_298),
.Y(n_405)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_378),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_411),
.A2(n_375),
.B1(n_374),
.B2(n_364),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_382),
.A2(n_322),
.B1(n_315),
.B2(n_327),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_426),
.B1(n_410),
.B2(n_413),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_369),
.A2(n_322),
.B1(n_300),
.B2(n_330),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_413),
.A2(n_418),
.B1(n_422),
.B2(n_423),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_386),
.A2(n_330),
.B1(n_344),
.B2(n_341),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_360),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_421),
.A2(n_408),
.B(n_407),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_371),
.A2(n_344),
.B1(n_341),
.B2(n_318),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_359),
.A2(n_318),
.B1(n_336),
.B2(n_323),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_390),
.A2(n_327),
.B1(n_323),
.B2(n_336),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_366),
.B1(n_376),
.B2(n_377),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_370),
.A2(n_312),
.B1(n_317),
.B2(n_333),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_434),
.B1(n_436),
.B2(n_449),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_379),
.C(n_363),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_433),
.C(n_453),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_358),
.Y(n_430)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_430),
.Y(n_475)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_431),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_390),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_435),
.A2(n_405),
.B(n_394),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_381),
.Y(n_437)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_SL g438 ( 
.A(n_420),
.B(n_385),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_355),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_441),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_420),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_440),
.B(n_418),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_383),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_442),
.A2(n_451),
.B1(n_421),
.B2(n_395),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_392),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_444),
.B(n_445),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_425),
.B(n_387),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_368),
.Y(n_446)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_409),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_447),
.Y(n_470)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_406),
.Y(n_448)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_365),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_450),
.Y(n_478)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_408),
.A2(n_362),
.B(n_390),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_406),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_452),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_415),
.B(n_389),
.C(n_360),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_427),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_404),
.B(n_357),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_399),
.B(n_351),
.Y(n_457)
);

OAI31xp33_ASAP7_75t_L g502 ( 
.A1(n_463),
.A2(n_474),
.A3(n_434),
.B(n_437),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_432),
.A2(n_416),
.B1(n_400),
.B2(n_394),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_464),
.A2(n_479),
.B1(n_481),
.B2(n_431),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_421),
.C(n_401),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_467),
.C(n_468),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_440),
.B(n_421),
.C(n_417),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_429),
.B(n_417),
.C(n_412),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_469),
.B(n_477),
.C(n_435),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_442),
.A2(n_394),
.B1(n_398),
.B2(n_400),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_472),
.A2(n_480),
.B1(n_482),
.B2(n_436),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_433),
.B(n_423),
.C(n_424),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_432),
.A2(n_394),
.B1(n_422),
.B2(n_426),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_443),
.A2(n_419),
.B1(n_397),
.B2(n_396),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_428),
.A2(n_397),
.B1(n_393),
.B2(n_388),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_443),
.A2(n_393),
.B1(n_335),
.B2(n_317),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_312),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_457),
.Y(n_498)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_478),
.Y(n_484)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_484),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_459),
.B(n_451),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_496),
.Y(n_508)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_461),
.Y(n_486)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_461),
.Y(n_488)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_488),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_489),
.A2(n_492),
.B1(n_500),
.B2(n_502),
.Y(n_515)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_458),
.Y(n_490)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_490),
.Y(n_519)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_478),
.Y(n_491)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_491),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_460),
.A2(n_479),
.B1(n_464),
.B2(n_472),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_476),
.Y(n_493)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_493),
.Y(n_511)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_465),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_494),
.B(n_499),
.Y(n_520)
);

INVx6_ASAP7_75t_L g495 ( 
.A(n_471),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_495),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_451),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_497),
.A2(n_463),
.B1(n_475),
.B2(n_481),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_498),
.B(n_501),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_462),
.B(n_447),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_470),
.A2(n_449),
.B1(n_441),
.B2(n_439),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_466),
.B(n_430),
.C(n_455),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_504),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_476),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_500),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_510),
.A2(n_480),
.B1(n_498),
.B2(n_469),
.Y(n_534)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_512),
.Y(n_530)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_502),
.A2(n_474),
.B(n_477),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_514),
.A2(n_489),
.B(n_492),
.Y(n_532)
);

BUFx24_ASAP7_75t_SL g516 ( 
.A(n_495),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_516),
.B(n_468),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_506),
.B(n_503),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_525),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_521),
.Y(n_523)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g524 ( 
.A(n_508),
.B(n_485),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_524),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_520),
.B(n_475),
.Y(n_526)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_526),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_513),
.B(n_496),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_527),
.B(n_528),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_519),
.B(n_487),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_507),
.B(n_484),
.Y(n_529)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_529),
.B(n_532),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_487),
.C(n_501),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_531),
.B(n_483),
.C(n_514),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_467),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_518),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_534),
.A2(n_510),
.B1(n_515),
.B2(n_517),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g548 ( 
.A(n_535),
.B(n_541),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_542),
.B(n_530),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_509),
.C(n_507),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_509),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_536),
.A2(n_523),
.B(n_531),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g553 ( 
.A1(n_545),
.A2(n_549),
.B(n_538),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_537),
.B(n_533),
.C(n_532),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_546),
.B(n_547),
.Y(n_552)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_543),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_539),
.A2(n_534),
.B(n_529),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_550),
.B(n_551),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_553),
.A2(n_538),
.B(n_541),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_548),
.B(n_544),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_555),
.B(n_551),
.Y(n_556)
);

A2O1A1Ixp33_ASAP7_75t_SL g558 ( 
.A1(n_556),
.A2(n_554),
.B(n_552),
.C(n_512),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_557),
.A2(n_540),
.B(n_491),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_558),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_559),
.B(n_540),
.C(n_511),
.Y(n_561)
);

NAND2x1_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_511),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_452),
.Y(n_563)
);


endmodule