module fake_jpeg_26135_n_43 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_43);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_43;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_32;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_25),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_24),
.B(n_27),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_10),
.B1(n_14),
.B2(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_20),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_24),
.B(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_21),
.C(n_18),
.Y(n_29)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_32),
.B1(n_5),
.B2(n_12),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_11),
.B1(n_13),
.B2(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_38),
.A2(n_33),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_36),
.Y(n_41)
);

BUFx24_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_39),
.B1(n_16),
.B2(n_1),
.Y(n_43)
);


endmodule