module fake_jpeg_7066_n_41 (n_3, n_2, n_1, n_0, n_4, n_5, n_41);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_41;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_3),
.B(n_2),
.Y(n_6)
);

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_5),
.B(n_1),
.Y(n_8)
);

INVx4_ASAP7_75t_SL g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_4),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_20),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_0),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_15),
.A2(n_16),
.B(n_17),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g17 ( 
.A1(n_11),
.A2(n_2),
.B1(n_4),
.B2(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_11),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_15),
.B(n_16),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_8),
.B1(n_10),
.B2(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_16),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_20),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_32),
.B(n_33),
.Y(n_36)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_30),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

AND2x2_ASAP7_75t_SL g38 ( 
.A(n_35),
.B(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_35),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_36),
.B(n_39),
.Y(n_41)
);


endmodule