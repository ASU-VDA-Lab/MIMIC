module fake_aes_2737_n_22 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_22;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_6), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_9), .B(n_7), .Y(n_14) );
OR2x6_ASAP7_75t_SL g15 ( .A(n_13), .B(n_0), .Y(n_15) );
BUFx2_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_15), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_17), .B(n_13), .Y(n_18) );
NOR3xp33_ASAP7_75t_L g19 ( .A(n_18), .B(n_11), .C(n_10), .Y(n_19) );
AOI211xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_12), .B(n_14), .C(n_3), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_1), .B1(n_4), .B2(n_5), .Y(n_22) );
endmodule