module fake_aes_11222_n_667 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_667);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_667;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g89 ( .A(n_63), .Y(n_89) );
INVx2_ASAP7_75t_SL g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_52), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_13), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_49), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_77), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_73), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_78), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_61), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_56), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_31), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_38), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_59), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_87), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_45), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_3), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_9), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_88), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_32), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_69), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_37), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_65), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_24), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_26), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_47), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_60), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_19), .Y(n_117) );
INVxp67_ASAP7_75t_L g118 ( .A(n_17), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_21), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_57), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_9), .Y(n_121) );
INVxp67_ASAP7_75t_L g122 ( .A(n_51), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_50), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_68), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_4), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_3), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_43), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_39), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_105), .B(n_0), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_90), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_105), .Y(n_134) );
OAI21x1_ASAP7_75t_L g135 ( .A1(n_98), .A2(n_36), .B(n_84), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_90), .B(n_1), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_105), .B(n_1), .Y(n_137) );
HB1xp67_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
INVx2_ASAP7_75t_SL g139 ( .A(n_89), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_98), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_106), .B(n_2), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_102), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_102), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_106), .B(n_2), .Y(n_144) );
NOR2xp33_ASAP7_75t_SL g145 ( .A(n_108), .B(n_40), .Y(n_145) );
INVx4_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g148 ( .A(n_121), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_91), .B(n_94), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_102), .B(n_5), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_92), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_99), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_114), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_114), .B(n_6), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_119), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_94), .Y(n_158) );
INVx4_ASAP7_75t_SL g159 ( .A(n_151), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
BUFx2_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_146), .B(n_117), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_146), .B(n_116), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_150), .B(n_96), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_151), .Y(n_170) );
NAND2xp33_ASAP7_75t_SL g171 ( .A(n_146), .B(n_111), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g172 ( .A1(n_151), .A2(n_127), .B1(n_129), .B2(n_128), .Y(n_172) );
INVxp67_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_149), .B(n_96), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_139), .B(n_93), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_139), .B(n_95), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_139), .B(n_97), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_150), .B(n_122), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_156), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_147), .B(n_130), .Y(n_183) );
BUFx2_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
INVx4_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
INVx1_ASAP7_75t_SL g186 ( .A(n_148), .Y(n_186) );
INVx5_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_140), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx4_ASAP7_75t_SL g190 ( .A(n_156), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_143), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_166), .B(n_131), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_169), .B(n_147), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_163), .B(n_145), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_161), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_169), .B(n_158), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g198 ( .A1(n_173), .A2(n_152), .B1(n_145), .B2(n_136), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
OR2x6_ASAP7_75t_L g200 ( .A(n_163), .B(n_137), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_169), .B(n_158), .Y(n_201) );
NAND2xp33_ASAP7_75t_L g202 ( .A(n_182), .B(n_101), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_181), .A2(n_156), .B1(n_137), .B2(n_136), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_169), .B(n_156), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_178), .Y(n_206) );
INVx1_ASAP7_75t_SL g207 ( .A(n_186), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g208 ( .A1(n_170), .A2(n_137), .B(n_155), .C(n_135), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_159), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_183), .B(n_132), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_185), .A2(n_137), .B1(n_155), .B2(n_132), .Y(n_211) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_160), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_164), .B(n_141), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_175), .B(n_141), .Y(n_215) );
AOI22xp33_ASAP7_75t_L g216 ( .A1(n_185), .A2(n_155), .B1(n_144), .B2(n_157), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_178), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_179), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_167), .Y(n_219) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_162), .B(n_135), .Y(n_220) );
AND3x1_ASAP7_75t_L g221 ( .A(n_172), .B(n_152), .C(n_176), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_159), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_159), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_185), .A2(n_144), .B1(n_157), .B2(n_153), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_157), .B1(n_154), .B2(n_153), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_167), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_179), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_171), .A2(n_113), .B1(n_101), .B2(n_103), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_168), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_184), .A2(n_123), .B1(n_103), .B2(n_104), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_180), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_168), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_162), .B(n_100), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_174), .B(n_134), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_162), .B(n_109), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_162), .B(n_134), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_184), .B(n_142), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_207), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_227), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_202), .A2(n_165), .B(n_182), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_179), .B1(n_170), .B2(n_188), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_198), .A2(n_170), .B(n_191), .C(n_189), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_215), .B(n_159), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_200), .A2(n_191), .B1(n_189), .B2(n_188), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_212), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_220), .A2(n_135), .B(n_192), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_231), .B(n_190), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_210), .B(n_190), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_202), .A2(n_177), .B(n_192), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_203), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_193), .B(n_190), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_236), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_227), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_208), .A2(n_177), .B(n_104), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_193), .B(n_190), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_214), .A2(n_124), .B(n_110), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_200), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_213), .Y(n_259) );
O2A1O1Ixp5_ASAP7_75t_L g260 ( .A1(n_195), .A2(n_119), .B(n_110), .C(n_112), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_213), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_205), .A2(n_201), .B(n_194), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_219), .Y(n_263) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_227), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_219), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_227), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_197), .A2(n_125), .B(n_112), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_233), .A2(n_128), .B(n_115), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_200), .A2(n_142), .B1(n_115), .B2(n_120), .Y(n_269) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_227), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_234), .B(n_107), .Y(n_271) );
INVx1_ASAP7_75t_SL g272 ( .A(n_234), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_230), .B(n_129), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_209), .B(n_187), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_235), .A2(n_125), .B(n_123), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_211), .B(n_124), .Y(n_276) );
OAI21xp5_ASAP7_75t_L g277 ( .A1(n_220), .A2(n_226), .B(n_232), .Y(n_277) );
INVx4_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_226), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_221), .B(n_7), .Y(n_280) );
BUFx6f_ASAP7_75t_L g281 ( .A(n_209), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_250), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
NOR2x1_ASAP7_75t_R g284 ( .A(n_258), .B(n_218), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_250), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_238), .Y(n_286) );
O2A1O1Ixp33_ASAP7_75t_L g287 ( .A1(n_280), .A2(n_237), .B(n_216), .C(n_229), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_245), .A2(n_228), .B1(n_204), .B2(n_229), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_272), .A2(n_232), .B1(n_224), .B2(n_223), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_271), .B(n_222), .Y(n_290) );
BUFx4f_ASAP7_75t_SL g291 ( .A(n_245), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_246), .A2(n_220), .B(n_225), .Y(n_292) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_262), .A2(n_120), .B(n_143), .C(n_153), .Y(n_293) );
NOR2xp67_ASAP7_75t_L g294 ( .A(n_258), .B(n_8), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_246), .A2(n_217), .B(n_206), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_252), .B(n_153), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_273), .B(n_153), .Y(n_297) );
AO31x2_ASAP7_75t_L g298 ( .A1(n_254), .A2(n_217), .A3(n_206), .B(n_199), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_256), .B(n_143), .Y(n_299) );
O2A1O1Ixp5_ASAP7_75t_L g300 ( .A1(n_277), .A2(n_199), .B(n_196), .C(n_154), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_256), .B(n_153), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_261), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_269), .Y(n_303) );
CKINVDCx8_ASAP7_75t_R g304 ( .A(n_255), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_242), .A2(n_154), .B(n_196), .C(n_187), .Y(n_305) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_276), .A2(n_154), .B1(n_187), .B2(n_11), .C(n_12), .Y(n_306) );
OAI21xp5_ASAP7_75t_L g307 ( .A1(n_243), .A2(n_187), .B(n_154), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_259), .B(n_154), .Y(n_308) );
OAI221xp5_ASAP7_75t_L g309 ( .A1(n_251), .A2(n_187), .B1(n_10), .B2(n_11), .C(n_12), .Y(n_309) );
NAND3xp33_ASAP7_75t_L g310 ( .A(n_260), .B(n_187), .C(n_10), .Y(n_310) );
AOI222xp33_ASAP7_75t_L g311 ( .A1(n_263), .A2(n_8), .B1(n_13), .B2(n_14), .C1(n_15), .C2(n_16), .Y(n_311) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_244), .A2(n_14), .B1(n_15), .B2(n_16), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_259), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_264), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_255), .B(n_17), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_240), .A2(n_53), .B(n_83), .Y(n_316) );
INVxp33_ASAP7_75t_SL g317 ( .A(n_241), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_317), .A2(n_255), .B1(n_279), .B2(n_248), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_305), .A2(n_265), .B(n_275), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_305), .A2(n_268), .B(n_249), .Y(n_320) );
OA21x2_ASAP7_75t_L g321 ( .A1(n_300), .A2(n_265), .B(n_267), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_291), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_286), .B(n_283), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_282), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_302), .B(n_248), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_293), .A2(n_257), .B(n_274), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_282), .Y(n_327) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_295), .A2(n_274), .B(n_247), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_285), .B(n_253), .Y(n_329) );
OAI22xp5_ASAP7_75t_SL g330 ( .A1(n_303), .A2(n_278), .B1(n_253), .B2(n_239), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_285), .B(n_253), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_313), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_315), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_313), .B(n_278), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_296), .A2(n_239), .B(n_270), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_288), .B(n_239), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_314), .Y(n_337) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_293), .A2(n_270), .B(n_266), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_317), .B(n_278), .Y(n_339) );
AO31x2_ASAP7_75t_L g340 ( .A1(n_308), .A2(n_270), .A3(n_266), .B(n_264), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_314), .Y(n_341) );
BUFx4f_ASAP7_75t_SL g342 ( .A(n_315), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_295), .A2(n_270), .B(n_266), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_297), .A2(n_266), .B(n_264), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_287), .B(n_264), .Y(n_346) );
OA21x2_ASAP7_75t_L g347 ( .A1(n_292), .A2(n_281), .B(n_54), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_342), .A2(n_303), .B1(n_315), .B2(n_304), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_327), .B(n_299), .Y(n_349) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_343), .A2(n_307), .B(n_292), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_323), .B(n_284), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_327), .B(n_301), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_332), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_332), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_343), .A2(n_306), .B(n_312), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_346), .A2(n_316), .B(n_310), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_333), .B(n_314), .Y(n_357) );
INVx3_ASAP7_75t_L g358 ( .A(n_324), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_333), .A2(n_294), .B(n_309), .C(n_290), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g360 ( .A1(n_339), .A2(n_304), .B1(n_289), .B2(n_314), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_344), .B(n_298), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_318), .A2(n_311), .B1(n_301), .B2(n_281), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_324), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_339), .B(n_281), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_324), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_344), .B(n_334), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g367 ( .A1(n_319), .A2(n_298), .B(n_281), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_329), .Y(n_369) );
OA21x2_ASAP7_75t_L g370 ( .A1(n_346), .A2(n_298), .B(n_48), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_329), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_322), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_331), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_336), .B(n_298), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
INVx3_ASAP7_75t_L g377 ( .A(n_368), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_361), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_361), .B(n_338), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_368), .Y(n_380) );
AND2x2_ASAP7_75t_SL g381 ( .A(n_370), .B(n_347), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_368), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_361), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_358), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_361), .B(n_338), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_348), .A2(n_336), .B1(n_325), .B2(n_319), .C(n_326), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_376), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_363), .B(n_338), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_363), .B(n_338), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_365), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_369), .B(n_325), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_354), .B(n_340), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_366), .B(n_340), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_376), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_358), .B(n_340), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_376), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_376), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_358), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_350), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_374), .B(n_340), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_350), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_369), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_367), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_374), .B(n_328), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_366), .B(n_328), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_407), .B(n_375), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_392), .B(n_348), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_392), .B(n_372), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_391), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_388), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_407), .B(n_375), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_397), .B(n_350), .Y(n_418) );
OR2x2_ASAP7_75t_L g419 ( .A(n_397), .B(n_373), .Y(n_419) );
NOR2xp33_ASAP7_75t_R g420 ( .A(n_403), .B(n_351), .Y(n_420) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_395), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_391), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_388), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_393), .B(n_373), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_393), .Y(n_426) );
AND2x4_ASAP7_75t_SL g427 ( .A(n_396), .B(n_364), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_394), .B(n_371), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_396), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_411), .B(n_350), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_394), .B(n_371), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_405), .B(n_349), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_396), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_405), .B(n_349), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_395), .B(n_360), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g437 ( .A1(n_378), .A2(n_360), .B1(n_362), .B2(n_364), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_405), .B(n_352), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_411), .B(n_352), .Y(n_439) );
NOR4xp25_ASAP7_75t_SL g440 ( .A(n_386), .B(n_359), .C(n_330), .D(n_355), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_411), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_409), .B(n_364), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_380), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_410), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_378), .B(n_364), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_409), .B(n_355), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_380), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_382), .B(n_334), .Y(n_448) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_383), .B(n_330), .Y(n_449) );
NOR2x1_ASAP7_75t_L g450 ( .A(n_387), .B(n_357), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_377), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_382), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_383), .B(n_367), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_379), .B(n_370), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_379), .B(n_370), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_389), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_389), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_409), .B(n_355), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_379), .B(n_370), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_390), .B(n_355), .Y(n_460) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_377), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_399), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_416), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_418), .B(n_385), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_441), .B(n_398), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_418), .B(n_385), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_413), .B(n_390), .Y(n_468) );
OAI332xp33_ASAP7_75t_L g469 ( .A1(n_413), .A2(n_386), .A3(n_400), .B1(n_398), .B2(n_404), .B3(n_406), .C1(n_19), .C2(n_18), .Y(n_469) );
OAI21xp33_ASAP7_75t_L g470 ( .A1(n_460), .A2(n_400), .B(n_408), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_430), .B(n_399), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_421), .B(n_387), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_456), .B(n_402), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_422), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_457), .B(n_402), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_430), .B(n_399), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_432), .B(n_408), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_426), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_420), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_422), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_420), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_462), .B(n_377), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_425), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_428), .Y(n_487) );
NOR2x1_ASAP7_75t_L g488 ( .A(n_450), .B(n_414), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_435), .B(n_377), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_453), .B(n_406), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_414), .B(n_403), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_439), .B(n_384), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_423), .Y(n_493) );
INVx2_ASAP7_75t_SL g494 ( .A(n_427), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_423), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_438), .B(n_406), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_458), .B(n_404), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_453), .B(n_404), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_419), .B(n_384), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_412), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_458), .B(n_401), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_417), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_453), .B(n_384), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_434), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_446), .B(n_401), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_429), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_447), .B(n_401), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_452), .B(n_403), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_436), .B(n_403), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_454), .B(n_381), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_429), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_454), .B(n_381), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_449), .B(n_381), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_455), .B(n_356), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_448), .Y(n_516) );
INVxp67_ASAP7_75t_SL g517 ( .A(n_461), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_442), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_433), .B(n_357), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_449), .B(n_18), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_445), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_445), .Y(n_522) );
OAI31xp33_ASAP7_75t_L g523 ( .A1(n_482), .A2(n_427), .A3(n_436), .B(n_433), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_494), .B(n_444), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_478), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_486), .B(n_455), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_463), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_474), .Y(n_528) );
NOR2xp67_ASAP7_75t_L g529 ( .A(n_494), .B(n_459), .Y(n_529) );
OAI22xp33_ASAP7_75t_L g530 ( .A1(n_484), .A2(n_451), .B1(n_459), .B2(n_347), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_471), .B(n_451), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_481), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_516), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_467), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_487), .B(n_437), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_518), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_471), .B(n_440), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_479), .B(n_357), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_498), .B(n_356), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_521), .Y(n_540) );
OA21x2_ASAP7_75t_L g541 ( .A1(n_470), .A2(n_337), .B(n_341), .Y(n_541) );
NAND2x1p5_ASAP7_75t_L g542 ( .A(n_519), .B(n_347), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_468), .B(n_357), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_472), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_501), .B(n_356), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_472), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_522), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_503), .B(n_356), .Y(n_548) );
NOR2xp33_ASAP7_75t_SL g549 ( .A(n_488), .B(n_357), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_465), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_485), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_479), .B(n_347), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_497), .B(n_320), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_465), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_504), .B(n_341), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_514), .A2(n_320), .B1(n_326), .B2(n_337), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_505), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_464), .B(n_328), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_517), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_480), .B(n_320), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_464), .B(n_328), .Y(n_561) );
INVx1_ASAP7_75t_SL g562 ( .A(n_492), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_466), .B(n_341), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_506), .Y(n_564) );
INVx2_ASAP7_75t_SL g565 ( .A(n_519), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_496), .B(n_320), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_506), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_466), .B(n_337), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_500), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_485), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_489), .B(n_321), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_511), .B(n_321), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_497), .B(n_321), .Y(n_573) );
OAI32xp33_ASAP7_75t_L g574 ( .A1(n_520), .A2(n_20), .A3(n_22), .B1(n_23), .B2(n_25), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_502), .B(n_321), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_559), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_525), .Y(n_577) );
AOI221xp5_ASAP7_75t_SL g578 ( .A1(n_533), .A2(n_491), .B1(n_513), .B2(n_511), .C(n_515), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_544), .B(n_475), .Y(n_579) );
OAI22xp33_ASAP7_75t_L g580 ( .A1(n_549), .A2(n_477), .B1(n_475), .B2(n_491), .Y(n_580) );
OAI31xp33_ASAP7_75t_L g581 ( .A1(n_537), .A2(n_513), .A3(n_504), .B(n_515), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_557), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_527), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_528), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_559), .B(n_509), .C(n_508), .Y(n_585) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_546), .Y(n_586) );
AOI221xp5_ASAP7_75t_SL g587 ( .A1(n_535), .A2(n_569), .B1(n_562), .B2(n_570), .C(n_526), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_535), .B(n_502), .Y(n_588) );
INVx3_ASAP7_75t_SL g589 ( .A(n_524), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_524), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_564), .B(n_490), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_550), .B(n_477), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_536), .A2(n_469), .B1(n_490), .B2(n_499), .C(n_504), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_529), .A2(n_523), .B(n_530), .Y(n_595) );
NAND2xp33_ASAP7_75t_L g596 ( .A(n_565), .B(n_510), .Y(n_596) );
XNOR2xp5_ASAP7_75t_L g597 ( .A(n_563), .B(n_519), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_532), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_543), .A2(n_490), .B1(n_499), .B2(n_510), .Y(n_599) );
NAND2xp33_ASAP7_75t_SL g600 ( .A(n_538), .B(n_512), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_534), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
OAI21xp5_ASAP7_75t_L g603 ( .A1(n_530), .A2(n_499), .B(n_507), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_567), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_526), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_551), .B(n_531), .Y(n_606) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_539), .Y(n_607) );
OAI21xp5_ASAP7_75t_L g608 ( .A1(n_539), .A2(n_507), .B(n_495), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_540), .B(n_495), .Y(n_609) );
NAND4xp75_ASAP7_75t_L g610 ( .A(n_543), .B(n_493), .C(n_483), .D(n_476), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_547), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_576), .A2(n_574), .B(n_545), .C(n_548), .Y(n_612) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_578), .A2(n_558), .A3(n_561), .B1(n_572), .B2(n_553), .C1(n_548), .C2(n_545), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_605), .B(n_560), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_587), .B(n_568), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_594), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_600), .A2(n_553), .B1(n_555), .B2(n_573), .Y(n_617) );
OAI31xp33_ASAP7_75t_L g618 ( .A1(n_600), .A2(n_552), .A3(n_542), .B(n_566), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_595), .A2(n_573), .B(n_575), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_609), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_599), .A2(n_555), .B1(n_575), .B2(n_556), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_582), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_589), .B(n_571), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_596), .A2(n_541), .B1(n_542), .B2(n_493), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_581), .B(n_541), .C(n_483), .Y(n_625) );
AOI21xp5_ASAP7_75t_L g626 ( .A1(n_596), .A2(n_541), .B(n_476), .Y(n_626) );
NOR3xp33_ASAP7_75t_L g627 ( .A(n_603), .B(n_473), .C(n_467), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_607), .A2(n_473), .B1(n_335), .B2(n_345), .C(n_30), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_589), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_588), .B(n_33), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_580), .B(n_34), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_583), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_577), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_617), .A2(n_590), .B1(n_597), .B2(n_610), .Y(n_634) );
A2O1A1Ixp33_ASAP7_75t_L g635 ( .A1(n_613), .A2(n_593), .B(n_585), .C(n_591), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_620), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_619), .A2(n_602), .B1(n_584), .B2(n_598), .C(n_604), .Y(n_637) );
NAND4xp75_ASAP7_75t_L g638 ( .A(n_631), .B(n_591), .C(n_592), .D(n_608), .Y(n_638) );
O2A1O1Ixp5_ASAP7_75t_L g639 ( .A1(n_615), .A2(n_611), .B(n_594), .C(n_601), .Y(n_639) );
NOR4xp25_ASAP7_75t_L g640 ( .A(n_612), .B(n_579), .C(n_601), .D(n_606), .Y(n_640) );
NOR2xp33_ASAP7_75t_R g641 ( .A(n_630), .B(n_597), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_623), .A2(n_586), .B1(n_579), .B2(n_606), .Y(n_642) );
NAND2xp33_ASAP7_75t_SL g643 ( .A(n_629), .B(n_610), .Y(n_643) );
OAI21xp33_ASAP7_75t_L g644 ( .A1(n_621), .A2(n_41), .B(n_42), .Y(n_644) );
BUFx3_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g646 ( .A1(n_629), .A2(n_44), .B(n_46), .Y(n_646) );
NOR4xp75_ASAP7_75t_L g647 ( .A(n_638), .B(n_614), .C(n_618), .D(n_625), .Y(n_647) );
XNOR2x2_ASAP7_75t_L g648 ( .A(n_634), .B(n_624), .Y(n_648) );
AOI21xp5_ASAP7_75t_L g649 ( .A1(n_643), .A2(n_626), .B(n_633), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_645), .B(n_632), .Y(n_650) );
NOR5xp2_ASAP7_75t_L g651 ( .A(n_635), .B(n_627), .C(n_628), .D(n_616), .E(n_66), .Y(n_651) );
AOI211xp5_ASAP7_75t_L g652 ( .A1(n_640), .A2(n_55), .B(n_58), .C(n_64), .Y(n_652) );
OAI21xp5_ASAP7_75t_L g653 ( .A1(n_639), .A2(n_67), .B(n_70), .Y(n_653) );
NAND4xp75_ASAP7_75t_L g654 ( .A(n_649), .B(n_639), .C(n_646), .D(n_637), .Y(n_654) );
NOR2xp67_ASAP7_75t_SL g655 ( .A(n_653), .B(n_636), .Y(n_655) );
BUFx2_ASAP7_75t_L g656 ( .A(n_648), .Y(n_656) );
NOR2xp67_ASAP7_75t_L g657 ( .A(n_650), .B(n_642), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_656), .Y(n_658) );
AND2x4_ASAP7_75t_SL g659 ( .A(n_657), .B(n_647), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_654), .A2(n_652), .B1(n_644), .B2(n_651), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_658), .B(n_655), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_659), .Y(n_662) );
AOI22x1_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_661), .B1(n_660), .B2(n_641), .Y(n_663) );
OAI21xp5_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_71), .B(n_72), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g665 ( .A1(n_664), .A2(n_74), .B(n_75), .Y(n_665) );
NAND3x2_ASAP7_75t_L g666 ( .A(n_665), .B(n_76), .C(n_79), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_666), .A2(n_80), .B1(n_81), .B2(n_85), .Y(n_667) );
endmodule