module real_aes_18119_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1441;
wire n_1382;
wire n_875;
wire n_951;
wire n_1225;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_1380;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_1011;
wire n_286;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1403;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_1463;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1455;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_1097;
wire n_703;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVx1_ASAP7_75t_L g746 ( .A(n_0), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_1), .A2(n_4), .B1(n_1156), .B2(n_1159), .Y(n_1155) );
AOI221x1_ASAP7_75t_SL g757 ( .A1(n_2), .A2(n_240), .B1(n_758), .B2(n_759), .C(n_760), .Y(n_757) );
AOI21xp33_ASAP7_75t_L g825 ( .A1(n_2), .A2(n_451), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g687 ( .A(n_3), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g724 ( .A1(n_3), .A2(n_725), .B(n_726), .C(n_733), .Y(n_724) );
CKINVDCx5p33_ASAP7_75t_R g1388 ( .A(n_5), .Y(n_1388) );
CKINVDCx5p33_ASAP7_75t_R g954 ( .A(n_6), .Y(n_954) );
INVx1_ASAP7_75t_L g552 ( .A(n_7), .Y(n_552) );
INVx1_ASAP7_75t_L g647 ( .A(n_8), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_8), .A2(n_107), .B1(n_677), .B2(n_679), .Y(n_676) );
INVx1_ASAP7_75t_L g314 ( .A(n_9), .Y(n_314) );
OAI22xp33_ASAP7_75t_L g441 ( .A1(n_9), .A2(n_114), .B1(n_442), .B2(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g995 ( .A(n_10), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g1008 ( .A1(n_10), .A2(n_243), .B1(n_448), .B2(n_603), .Y(n_1008) );
OAI221xp5_ASAP7_75t_L g996 ( .A1(n_11), .A2(n_198), .B1(n_322), .B2(n_326), .C(n_997), .Y(n_996) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_11), .A2(n_198), .B1(n_1011), .B2(n_1012), .Y(n_1010) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_12), .A2(n_236), .B1(n_292), .B2(n_301), .C(n_730), .Y(n_989) );
AOI222xp33_ASAP7_75t_L g1018 ( .A1(n_12), .A2(n_64), .B1(n_133), .B2(n_405), .C1(n_574), .C2(n_577), .Y(n_1018) );
INVx1_ASAP7_75t_L g1074 ( .A(n_13), .Y(n_1074) );
INVx1_ASAP7_75t_L g263 ( .A(n_14), .Y(n_263) );
AND2x2_ASAP7_75t_L g288 ( .A(n_14), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g312 ( .A(n_14), .B(n_212), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_14), .B(n_273), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g1101 ( .A1(n_15), .A2(n_105), .B1(n_301), .B2(n_626), .C(n_628), .Y(n_1101) );
INVx1_ASAP7_75t_L g1123 ( .A(n_15), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_16), .A2(n_241), .B1(n_322), .B2(n_326), .C(n_332), .Y(n_321) );
INVx1_ASAP7_75t_L g431 ( .A(n_16), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g476 ( .A1(n_17), .A2(n_477), .B(n_481), .C(n_488), .Y(n_476) );
INVx1_ASAP7_75t_L g509 ( .A(n_17), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_18), .A2(n_167), .B1(n_413), .B2(n_842), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_18), .A2(n_91), .B1(n_653), .B2(n_732), .C(n_975), .Y(n_974) );
CKINVDCx5p33_ASAP7_75t_R g1350 ( .A(n_19), .Y(n_1350) );
INVx1_ASAP7_75t_L g944 ( .A(n_20), .Y(n_944) );
INVx2_ASAP7_75t_L g1152 ( .A(n_21), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_21), .B(n_100), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_21), .B(n_1158), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_22), .A2(n_145), .B1(n_463), .B2(n_467), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_22), .A2(n_145), .B1(n_514), .B2(n_516), .Y(n_513) );
INVx1_ASAP7_75t_L g1038 ( .A(n_23), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_24), .A2(n_127), .B1(n_374), .B2(n_782), .Y(n_781) );
OAI221xp5_ASAP7_75t_L g789 ( .A1(n_24), .A2(n_218), .B1(n_790), .B2(n_792), .C(n_794), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g1177 ( .A1(n_25), .A2(n_217), .B1(n_1156), .B2(n_1159), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_26), .Y(n_1358) );
OAI22xp33_ASAP7_75t_L g473 ( .A1(n_27), .A2(n_39), .B1(n_265), .B2(n_474), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_27), .A2(n_39), .B1(n_493), .B2(n_496), .Y(n_492) );
INVx1_ASAP7_75t_L g1042 ( .A(n_28), .Y(n_1042) );
OAI22xp33_ASAP7_75t_L g1379 ( .A1(n_29), .A2(n_242), .B1(n_265), .B2(n_1380), .Y(n_1379) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_29), .A2(n_242), .B1(n_493), .B2(n_1394), .Y(n_1393) );
INVxp67_ASAP7_75t_SL g1439 ( .A(n_30), .Y(n_1439) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_30), .A2(n_67), .B1(n_285), .B2(n_631), .Y(n_1453) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_31), .A2(n_190), .B1(n_404), .B2(n_707), .Y(n_942) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_31), .A2(n_60), .B1(n_906), .B2(n_960), .C(n_962), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g1102 ( .A1(n_32), .A2(n_77), .B1(n_631), .B2(n_632), .Y(n_1102) );
INVx1_ASAP7_75t_L g1127 ( .A(n_32), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1363 ( .A(n_33), .Y(n_1363) );
INVx1_ASAP7_75t_L g1425 ( .A(n_34), .Y(n_1425) );
INVx1_ASAP7_75t_L g595 ( .A(n_35), .Y(n_595) );
INVx1_ASAP7_75t_L g883 ( .A(n_36), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_36), .A2(n_244), .B1(n_1149), .B2(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g548 ( .A(n_37), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_38), .A2(n_219), .B1(n_715), .B2(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g727 ( .A(n_38), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_40), .A2(n_209), .B1(n_653), .B2(n_991), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_40), .A2(n_105), .B1(n_669), .B2(n_917), .Y(n_1128) );
INVx1_ASAP7_75t_L g1037 ( .A(n_41), .Y(n_1037) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_42), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_43), .A2(n_79), .B1(n_672), .B2(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g873 ( .A(n_43), .Y(n_873) );
AOI22xp5_ASAP7_75t_L g1170 ( .A1(n_44), .A2(n_228), .B1(n_1156), .B2(n_1159), .Y(n_1170) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_45), .A2(n_125), .B1(n_292), .B2(n_295), .C(n_301), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_45), .A2(n_82), .B1(n_404), .B2(n_428), .Y(n_427) );
AO22x1_ASAP7_75t_L g1174 ( .A1(n_46), .A2(n_58), .B1(n_1149), .B2(n_1153), .Y(n_1174) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_47), .A2(n_110), .B1(n_706), .B2(n_707), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_47), .A2(n_219), .B1(n_285), .B2(n_732), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_48), .A2(n_156), .B1(n_304), .B2(n_309), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_48), .A2(n_99), .B1(n_418), .B2(n_421), .Y(n_417) );
INVx1_ASAP7_75t_L g1441 ( .A(n_49), .Y(n_1441) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_49), .A2(n_123), .B1(n_991), .B2(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g544 ( .A(n_50), .Y(n_544) );
INVx1_ASAP7_75t_L g360 ( .A(n_51), .Y(n_360) );
INVx1_ASAP7_75t_L g390 ( .A(n_51), .Y(n_390) );
INVx1_ASAP7_75t_L g713 ( .A(n_52), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_52), .A2(n_226), .B1(n_285), .B2(n_732), .Y(n_731) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_53), .A2(n_593), .B1(n_680), .B2(n_681), .Y(n_592) );
INVxp67_ASAP7_75t_L g681 ( .A(n_53), .Y(n_681) );
INVxp67_ASAP7_75t_SL g999 ( .A(n_54), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_54), .A2(n_236), .B1(n_797), .B2(n_839), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_55), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_56), .Y(n_619) );
INVx1_ASAP7_75t_L g1111 ( .A(n_57), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_58), .A2(n_683), .B1(n_684), .B2(n_740), .Y(n_682) );
INVxp67_ASAP7_75t_L g740 ( .A(n_58), .Y(n_740) );
INVx1_ASAP7_75t_L g256 ( .A(n_59), .Y(n_256) );
AOI22xp33_ASAP7_75t_SL g951 ( .A1(n_60), .A2(n_175), .B1(n_405), .B2(n_839), .Y(n_951) );
INVx2_ASAP7_75t_L g366 ( .A(n_61), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_62), .Y(n_1360) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_63), .A2(n_135), .B1(n_516), .B2(n_1077), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1088 ( .A1(n_63), .A2(n_135), .B1(n_1089), .B2(n_1090), .Y(n_1088) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_64), .A2(n_143), .B1(n_991), .B2(n_992), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g1428 ( .A1(n_65), .A2(n_142), .B1(n_474), .B2(n_1429), .Y(n_1428) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_65), .A2(n_142), .B1(n_1068), .B2(n_1394), .Y(n_1458) );
INVx1_ASAP7_75t_L g1424 ( .A(n_66), .Y(n_1424) );
INVxp67_ASAP7_75t_SL g1447 ( .A(n_67), .Y(n_1447) );
OAI22xp5_ASAP7_75t_L g372 ( .A1(n_68), .A2(n_206), .B1(n_373), .B2(n_384), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_69), .A2(n_247), .B1(n_652), .B2(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g667 ( .A(n_69), .Y(n_667) );
INVx1_ASAP7_75t_L g560 ( .A(n_70), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_71), .A2(n_172), .B1(n_1149), .B2(n_1153), .Y(n_1171) );
INVx1_ASAP7_75t_L g371 ( .A(n_72), .Y(n_371) );
AO221x2_ASAP7_75t_L g1241 ( .A1(n_73), .A2(n_207), .B1(n_1156), .B2(n_1159), .C(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1404 ( .A(n_73), .Y(n_1404) );
AOI22xp5_ASAP7_75t_L g1411 ( .A1(n_73), .A2(n_1412), .B1(n_1459), .B2(n_1462), .Y(n_1411) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_74), .A2(n_121), .B1(n_1068), .B2(n_1070), .Y(n_1067) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_74), .A2(n_121), .B1(n_474), .B2(n_1081), .Y(n_1080) );
AOI221xp5_ASAP7_75t_L g1105 ( .A1(n_75), .A2(n_102), .B1(n_628), .B2(n_901), .C(n_1001), .Y(n_1105) );
INVxp67_ASAP7_75t_SL g1115 ( .A(n_75), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1381 ( .A1(n_76), .A2(n_238), .B1(n_463), .B2(n_467), .Y(n_1381) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_76), .A2(n_238), .B1(n_1402), .B2(n_1403), .Y(n_1401) );
INVxp67_ASAP7_75t_SL g1117 ( .A(n_77), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_78), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_78), .A2(n_201), .B1(n_327), .B2(n_370), .C(n_738), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g852 ( .A1(n_79), .A2(n_115), .B1(n_653), .B2(n_853), .C(n_855), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_80), .A2(n_107), .B1(n_631), .B2(n_632), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_80), .A2(n_182), .B1(n_669), .B2(n_672), .Y(n_668) );
INVx1_ASAP7_75t_L g487 ( .A(n_81), .Y(n_487) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_81), .A2(n_500), .B(n_502), .C(n_504), .Y(n_499) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_82), .Y(n_340) );
INVx1_ASAP7_75t_L g948 ( .A(n_83), .Y(n_948) );
XOR2x2_ASAP7_75t_L g456 ( .A(n_84), .B(n_457), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_85), .A2(n_161), .B1(n_534), .B2(n_762), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g935 ( .A(n_85), .B(n_514), .Y(n_935) );
INVx1_ASAP7_75t_L g1028 ( .A(n_86), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_87), .Y(n_849) );
OAI221xp5_ASAP7_75t_SL g613 ( .A1(n_88), .A2(n_89), .B1(n_614), .B2(n_616), .C(n_618), .Y(n_613) );
INVx1_ASAP7_75t_L g640 ( .A(n_88), .Y(n_640) );
INVx1_ASAP7_75t_L g656 ( .A(n_89), .Y(n_656) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_90), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g941 ( .A1(n_91), .A2(n_116), .B1(n_418), .B2(n_421), .Y(n_941) );
OA222x2_ASAP7_75t_L g748 ( .A1(n_92), .A2(n_191), .B1(n_218), .B2(n_749), .C1(n_751), .C2(n_755), .Y(n_748) );
INVx1_ASAP7_75t_L g806 ( .A(n_92), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_93), .A2(n_1414), .B1(n_1415), .B2(n_1416), .Y(n_1413) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_93), .Y(n_1414) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_94), .Y(n_258) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_94), .B(n_256), .Y(n_1150) );
OAI211xp5_ASAP7_75t_SL g986 ( .A1(n_95), .A2(n_987), .B(n_988), .C(n_993), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g1006 ( .A1(n_95), .A2(n_199), .B1(n_384), .B2(n_1007), .Y(n_1006) );
XNOR2xp5_ASAP7_75t_L g984 ( .A(n_96), .B(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1137 ( .A(n_97), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g846 ( .A(n_98), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_99), .A2(n_144), .B1(n_297), .B2(n_342), .C(n_344), .Y(n_341) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_100), .B(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1158 ( .A(n_100), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g897 ( .A1(n_101), .A2(n_180), .B1(n_285), .B2(n_732), .Y(n_897) );
INVxp67_ASAP7_75t_SL g915 ( .A(n_101), .Y(n_915) );
INVx1_ASAP7_75t_L g1125 ( .A(n_102), .Y(n_1125) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_103), .A2(n_108), .B1(n_409), .B2(n_807), .Y(n_840) );
INVx1_ASAP7_75t_L g876 ( .A(n_103), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g998 ( .A(n_104), .Y(n_998) );
INVx1_ASAP7_75t_L g835 ( .A(n_106), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g866 ( .A1(n_106), .A2(n_223), .B1(n_335), .B2(n_338), .Y(n_866) );
INVx1_ASAP7_75t_L g858 ( .A(n_108), .Y(n_858) );
INVx1_ASAP7_75t_L g604 ( .A(n_109), .Y(n_604) );
AOI21xp33_ASAP7_75t_L g729 ( .A1(n_110), .A2(n_650), .B(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_111), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g394 ( .A(n_111), .Y(n_394) );
INVx1_ASAP7_75t_L g426 ( .A(n_111), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_112), .A2(n_204), .B1(n_1149), .B2(n_1153), .Y(n_1148) );
INVx1_ASAP7_75t_L g1045 ( .A(n_113), .Y(n_1045) );
INVx1_ASAP7_75t_L g317 ( .A(n_114), .Y(n_317) );
AOI22xp33_ASAP7_75t_SL g844 ( .A1(n_115), .A2(n_146), .B1(n_428), .B2(n_839), .Y(n_844) );
INVx1_ASAP7_75t_L g964 ( .A(n_116), .Y(n_964) );
INVx1_ASAP7_75t_L g1426 ( .A(n_117), .Y(n_1426) );
INVxp67_ASAP7_75t_SL g947 ( .A(n_118), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g967 ( .A1(n_118), .A2(n_224), .B1(n_335), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_119), .A2(n_239), .B1(n_304), .B2(n_309), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_119), .A2(n_221), .B1(n_415), .B2(n_677), .Y(n_827) );
INVx1_ASAP7_75t_L g1075 ( .A(n_120), .Y(n_1075) );
OAI211xp5_ASAP7_75t_L g1082 ( .A1(n_120), .A2(n_488), .B(n_1083), .C(n_1084), .Y(n_1082) );
NOR2xp33_ASAP7_75t_L g1108 ( .A(n_122), .B(n_327), .Y(n_1108) );
INVxp67_ASAP7_75t_SL g1133 ( .A(n_122), .Y(n_1133) );
INVxp67_ASAP7_75t_SL g1434 ( .A(n_123), .Y(n_1434) );
INVx1_ASAP7_75t_L g698 ( .A(n_124), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_124), .A2(n_157), .B1(n_722), .B2(n_723), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_125), .A2(n_162), .B1(n_402), .B2(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g905 ( .A(n_126), .Y(n_905) );
INVx1_ASAP7_75t_L g808 ( .A(n_127), .Y(n_808) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_128), .Y(n_712) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_129), .Y(n_773) );
INVx1_ASAP7_75t_L g559 ( .A(n_130), .Y(n_559) );
INVx1_ASAP7_75t_L g955 ( .A(n_131), .Y(n_955) );
INVx1_ASAP7_75t_L g702 ( .A(n_132), .Y(n_702) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_132), .A2(n_297), .B(n_344), .Y(n_734) );
AOI221xp5_ASAP7_75t_L g1000 ( .A1(n_133), .A2(n_205), .B1(n_901), .B2(n_1001), .C(n_1002), .Y(n_1000) );
INVx1_ASAP7_75t_L g1049 ( .A(n_134), .Y(n_1049) );
INVx1_ASAP7_75t_L g1107 ( .A(n_136), .Y(n_1107) );
INVx1_ASAP7_75t_L g1110 ( .A(n_137), .Y(n_1110) );
OAI322xp33_ASAP7_75t_L g1113 ( .A1(n_137), .A2(n_586), .A3(n_606), .B1(n_708), .B2(n_1114), .C1(n_1118), .C2(n_1124), .Y(n_1113) );
AO22x1_ASAP7_75t_L g1175 ( .A1(n_138), .A2(n_215), .B1(n_1156), .B2(n_1159), .Y(n_1175) );
BUFx3_ASAP7_75t_L g359 ( .A(n_139), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_140), .A2(n_248), .B1(n_732), .B2(n_903), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_140), .A2(n_181), .B1(n_796), .B2(n_917), .Y(n_916) );
INVx1_ASAP7_75t_L g1098 ( .A(n_141), .Y(n_1098) );
INVx1_ASAP7_75t_L g1025 ( .A(n_143), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_144), .A2(n_156), .B1(n_409), .B2(n_413), .Y(n_408) );
AOI211xp5_ASAP7_75t_SL g870 ( .A1(n_146), .A2(n_871), .B(n_872), .C(n_875), .Y(n_870) );
CKINVDCx5p33_ASAP7_75t_R g946 ( .A(n_147), .Y(n_946) );
INVx1_ASAP7_75t_L g978 ( .A(n_148), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_149), .A2(n_165), .B1(n_1156), .B2(n_1159), .Y(n_1202) );
BUFx6f_ASAP7_75t_L g270 ( .A(n_150), .Y(n_270) );
INVx1_ASAP7_75t_L g1435 ( .A(n_151), .Y(n_1435) );
INVx1_ASAP7_75t_L g598 ( .A(n_152), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_153), .A2(n_183), .B1(n_421), .B2(n_842), .Y(n_841) );
INVx1_ASAP7_75t_L g857 ( .A(n_153), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g907 ( .A1(n_154), .A2(n_184), .B1(n_908), .B2(n_909), .C(n_910), .Y(n_907) );
INVx1_ASAP7_75t_L g927 ( .A(n_154), .Y(n_927) );
OAI22xp33_ASAP7_75t_SL g893 ( .A1(n_155), .A2(n_197), .B1(n_772), .B2(n_874), .Y(n_893) );
INVx1_ASAP7_75t_L g930 ( .A(n_155), .Y(n_930) );
INVx1_ASAP7_75t_L g697 ( .A(n_157), .Y(n_697) );
INVx1_ASAP7_75t_L g895 ( .A(n_158), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_158), .A2(n_248), .B1(n_796), .B2(n_922), .Y(n_921) );
AOI21xp5_ASAP7_75t_SL g900 ( .A1(n_159), .A2(n_649), .B(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g914 ( .A(n_159), .Y(n_914) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_160), .Y(n_899) );
INVx1_ASAP7_75t_L g929 ( .A(n_161), .Y(n_929) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_162), .Y(n_336) );
INVx1_ASAP7_75t_L g1445 ( .A(n_163), .Y(n_1445) );
INVx1_ASAP7_75t_L g531 ( .A(n_164), .Y(n_531) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_166), .Y(n_1130) );
INVx1_ASAP7_75t_L g963 ( .A(n_167), .Y(n_963) );
INVx1_ASAP7_75t_L g1420 ( .A(n_168), .Y(n_1420) );
INVx1_ASAP7_75t_L g1391 ( .A(n_169), .Y(n_1391) );
OAI211xp5_ASAP7_75t_L g1395 ( .A1(n_169), .A2(n_502), .B(n_1396), .C(n_1399), .Y(n_1395) );
INVx1_ASAP7_75t_L g1422 ( .A(n_170), .Y(n_1422) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_171), .Y(n_832) );
XOR2x2_ASAP7_75t_L g279 ( .A(n_173), .B(n_280), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g1178 ( .A1(n_173), .A2(n_229), .B1(n_1149), .B2(n_1153), .Y(n_1178) );
INVx1_ASAP7_75t_L g484 ( .A(n_174), .Y(n_484) );
INVx1_ASAP7_75t_L g976 ( .A(n_175), .Y(n_976) );
INVx1_ASAP7_75t_L g1103 ( .A(n_176), .Y(n_1103) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_177), .Y(n_1351) );
XOR2xp5_ASAP7_75t_L g1032 ( .A(n_178), .B(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1040 ( .A(n_179), .Y(n_1040) );
INVxp67_ASAP7_75t_L g920 ( .A(n_180), .Y(n_920) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_181), .A2(n_649), .B(n_650), .Y(n_896) );
AOI21xp33_ASAP7_75t_L g648 ( .A1(n_182), .A2(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g879 ( .A(n_183), .Y(n_879) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_184), .Y(n_932) );
INVx1_ASAP7_75t_L g1442 ( .A(n_185), .Y(n_1442) );
INVx1_ASAP7_75t_L g535 ( .A(n_186), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_187), .A2(n_225), .B1(n_1149), .B2(n_1153), .Y(n_1201) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_188), .Y(n_269) );
OAI211xp5_ASAP7_75t_L g1382 ( .A1(n_189), .A2(n_488), .B(n_1383), .C(n_1386), .Y(n_1382) );
INVx1_ASAP7_75t_L g1400 ( .A(n_189), .Y(n_1400) );
INVx1_ASAP7_75t_L g977 ( .A(n_190), .Y(n_977) );
INVx1_ASAP7_75t_L g795 ( .A(n_191), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g1365 ( .A(n_192), .Y(n_1365) );
INVx1_ASAP7_75t_L g693 ( .A(n_193), .Y(n_693) );
INVx1_ASAP7_75t_L g1437 ( .A(n_194), .Y(n_1437) );
CKINVDCx5p33_ASAP7_75t_R g786 ( .A(n_195), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_196), .A2(n_208), .B1(n_626), .B2(n_628), .C(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g663 ( .A(n_196), .Y(n_663) );
INVx1_ASAP7_75t_L g934 ( .A(n_197), .Y(n_934) );
AO22x1_ASAP7_75t_L g1191 ( .A1(n_200), .A2(n_216), .B1(n_1149), .B2(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g691 ( .A(n_201), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_202), .Y(n_1356) );
CKINVDCx16_ASAP7_75t_R g1243 ( .A(n_203), .Y(n_1243) );
INVxp67_ASAP7_75t_SL g1024 ( .A(n_205), .Y(n_1024) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_206), .A2(n_283), .B(n_290), .C(n_313), .Y(n_282) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_208), .A2(n_247), .B1(n_574), .B2(n_675), .Y(n_674) );
INVxp67_ASAP7_75t_SL g1119 ( .A(n_209), .Y(n_1119) );
AOI22xp5_ASAP7_75t_L g1164 ( .A1(n_210), .A2(n_235), .B1(n_1156), .B2(n_1159), .Y(n_1164) );
CKINVDCx5p33_ASAP7_75t_R g621 ( .A(n_211), .Y(n_621) );
BUFx3_ASAP7_75t_L g273 ( .A(n_212), .Y(n_273) );
INVx1_ASAP7_75t_L g289 ( .A(n_212), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g1354 ( .A(n_213), .Y(n_1354) );
CKINVDCx20_ASAP7_75t_R g1245 ( .A(n_214), .Y(n_1245) );
INVx1_ASAP7_75t_L g546 ( .A(n_220), .Y(n_546) );
INVx1_ASAP7_75t_L g761 ( .A(n_221), .Y(n_761) );
CKINVDCx5p33_ASAP7_75t_R g769 ( .A(n_222), .Y(n_769) );
INVx1_ASAP7_75t_L g881 ( .A(n_223), .Y(n_881) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_224), .Y(n_957) );
INVx1_ASAP7_75t_L g704 ( .A(n_226), .Y(n_704) );
INVx2_ASAP7_75t_L g351 ( .A(n_227), .Y(n_351) );
INVx1_ASAP7_75t_L g364 ( .A(n_227), .Y(n_364) );
INVx1_ASAP7_75t_L g369 ( .A(n_227), .Y(n_369) );
AO22x1_ASAP7_75t_L g1193 ( .A1(n_230), .A2(n_246), .B1(n_1156), .B2(n_1159), .Y(n_1193) );
CKINVDCx5p33_ASAP7_75t_R g787 ( .A(n_231), .Y(n_787) );
INVx1_ASAP7_75t_L g1052 ( .A(n_232), .Y(n_1052) );
INVx1_ASAP7_75t_L g886 ( .A(n_233), .Y(n_886) );
OAI211xp5_ASAP7_75t_L g1071 ( .A1(n_234), .A2(n_500), .B(n_1072), .C(n_1073), .Y(n_1071) );
INVx1_ASAP7_75t_L g1087 ( .A(n_234), .Y(n_1087) );
INVx1_ASAP7_75t_L g1047 ( .A(n_237), .Y(n_1047) );
INVx1_ASAP7_75t_L g821 ( .A(n_239), .Y(n_821) );
INVx1_ASAP7_75t_L g820 ( .A(n_240), .Y(n_820) );
INVx1_ASAP7_75t_L g436 ( .A(n_241), .Y(n_436) );
INVx1_ASAP7_75t_L g994 ( .A(n_243), .Y(n_994) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_245), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_274), .B(n_1140), .Y(n_249) );
BUFx4f_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_259), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g1410 ( .A(n_253), .B(n_262), .Y(n_1410) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1461 ( .A(n_255), .B(n_258), .Y(n_1461) );
INVx1_ASAP7_75t_L g1466 ( .A(n_255), .Y(n_1466) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g1468 ( .A(n_258), .B(n_1466), .Y(n_1468) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x4_ASAP7_75t_L g459 ( .A(n_262), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g302 ( .A(n_263), .B(n_273), .Y(n_302) );
AND2x4_ASAP7_75t_L g345 ( .A(n_263), .B(n_272), .Y(n_345) );
INVx1_ASAP7_75t_L g1081 ( .A(n_264), .Y(n_1081) );
AND2x4_ASAP7_75t_SL g1409 ( .A(n_264), .B(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1429 ( .A(n_264), .Y(n_1429) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_271), .Y(n_265) );
OR2x6_ASAP7_75t_L g465 ( .A(n_266), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g335 ( .A(n_267), .Y(n_335) );
BUFx4f_ASAP7_75t_L g878 ( .A(n_267), .Y(n_878) );
INVx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
INVx2_ASAP7_75t_L g287 ( .A(n_269), .Y(n_287) );
AND2x2_ASAP7_75t_L g294 ( .A(n_269), .B(n_270), .Y(n_294) );
AND2x2_ASAP7_75t_L g299 ( .A(n_269), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g307 ( .A(n_269), .Y(n_307) );
INVx1_ASAP7_75t_L g377 ( .A(n_269), .Y(n_377) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_269), .B(n_270), .Y(n_480) );
AND2x2_ASAP7_75t_L g286 ( .A(n_270), .B(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g300 ( .A(n_270), .Y(n_300) );
INVx1_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
BUFx2_ASAP7_75t_L g330 ( .A(n_270), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_270), .B(n_287), .Y(n_339) );
OR2x2_ASAP7_75t_L g543 ( .A(n_270), .B(n_307), .Y(n_543) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g490 ( .A(n_272), .Y(n_490) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g472 ( .A(n_273), .Y(n_472) );
AND2x4_ASAP7_75t_L g486 ( .A(n_273), .B(n_376), .Y(n_486) );
XNOR2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_982), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_741), .B1(n_980), .B2(n_981), .Y(n_275) );
INVx2_ASAP7_75t_SL g980 ( .A(n_276), .Y(n_980) );
AO22x1_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B1(n_590), .B2(n_591), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
XNOR2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_456), .Y(n_278) );
NAND3xp33_ASAP7_75t_L g280 ( .A(n_281), .B(n_352), .C(n_396), .Y(n_280) );
OAI21xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_321), .B(n_346), .Y(n_281) );
INVx2_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g987 ( .A(n_284), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_284), .A2(n_319), .B1(n_1110), .B2(n_1111), .Y(n_1109) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
INVx1_ASAP7_75t_L g961 ( .A(n_285), .Y(n_961) );
BUFx2_ASAP7_75t_L g992 ( .A(n_285), .Y(n_992) );
HB1xp67_ASAP7_75t_L g1451 ( .A(n_285), .Y(n_1451) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
BUFx3_ASAP7_75t_L g632 ( .A(n_286), .Y(n_632) );
BUFx3_ASAP7_75t_L g653 ( .A(n_286), .Y(n_653) );
AND2x2_ASAP7_75t_L g316 ( .A(n_288), .B(n_306), .Y(n_316) );
AND2x4_ASAP7_75t_L g319 ( .A(n_288), .B(n_320), .Y(n_319) );
AND2x4_ASAP7_75t_SL g325 ( .A(n_288), .B(n_293), .Y(n_325) );
AND2x2_ASAP7_75t_L g611 ( .A(n_288), .B(n_320), .Y(n_611) );
AND2x2_ASAP7_75t_L g655 ( .A(n_288), .B(n_309), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_288), .B(n_369), .Y(n_754) );
BUFx2_ASAP7_75t_L g862 ( .A(n_288), .Y(n_862) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_289), .Y(n_466) );
AOI21xp5_ASAP7_75t_SL g290 ( .A1(n_291), .A2(n_303), .B(n_311), .Y(n_290) );
AOI222xp33_ASAP7_75t_L g1423 ( .A1(n_292), .A2(n_482), .B1(n_1424), .B2(n_1425), .C1(n_1426), .C2(n_1427), .Y(n_1423) );
BUFx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x6_ASAP7_75t_L g311 ( .A(n_293), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g343 ( .A(n_293), .Y(n_343) );
AND2x2_ASAP7_75t_L g489 ( .A(n_293), .B(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g628 ( .A(n_293), .Y(n_628) );
BUFx3_ASAP7_75t_L g871 ( .A(n_293), .Y(n_871) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_293), .Y(n_1002) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g643 ( .A(n_294), .Y(n_643) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g758 ( .A(n_296), .Y(n_758) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g730 ( .A(n_298), .Y(n_730) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_299), .Y(n_320) );
AND2x4_ASAP7_75t_L g475 ( .A(n_299), .B(n_466), .Y(n_475) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_299), .Y(n_1001) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_302), .B(n_556), .Y(n_555) );
INVx4_ASAP7_75t_L g650 ( .A(n_302), .Y(n_650) );
AND2x4_ASAP7_75t_L g776 ( .A(n_302), .B(n_556), .Y(n_776) );
OAI21xp33_ASAP7_75t_L g872 ( .A1(n_302), .A2(n_873), .B(n_874), .Y(n_872) );
OAI221xp5_ASAP7_75t_L g975 ( .A1(n_302), .A2(n_479), .B1(n_874), .B2(n_976), .C(n_977), .Y(n_975) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g631 ( .A(n_305), .Y(n_631) );
INVx2_ASAP7_75t_SL g635 ( .A(n_305), .Y(n_635) );
INVx1_ASAP7_75t_L g652 ( .A(n_305), .Y(n_652) );
INVx3_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_306), .B(n_312), .Y(n_370) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_306), .Y(n_732) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_307), .Y(n_638) );
AND2x4_ASAP7_75t_L g752 ( .A(n_309), .B(n_753), .Y(n_752) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g903 ( .A(n_310), .Y(n_903) );
AOI211xp5_ASAP7_75t_SL g736 ( .A1(n_311), .A2(n_657), .B(n_693), .C(n_737), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g988 ( .A1(n_311), .A2(n_989), .B(n_990), .Y(n_988) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_311), .A2(n_657), .B1(n_1101), .B2(n_1102), .C(n_1103), .Y(n_1100) );
INVx1_ASAP7_75t_L g331 ( .A(n_312), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_312), .B(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_312), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_312), .B(n_351), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_317), .B2(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g722 ( .A(n_315), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_315), .A2(n_319), .B1(n_994), .B2(n_995), .Y(n_993) );
AOI221xp5_ASAP7_75t_SL g1104 ( .A1(n_315), .A2(n_1105), .B1(n_1106), .B2(n_1107), .C(n_1108), .Y(n_1104) );
BUFx6f_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g601 ( .A(n_316), .B(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g725 ( .A(n_319), .Y(n_725) );
INVx1_ASAP7_75t_L g627 ( .A(n_320), .Y(n_627) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_320), .Y(n_649) );
INVx2_ASAP7_75t_L g865 ( .A(n_320), .Y(n_865) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx4_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g657 ( .A(n_325), .Y(n_657) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NOR2x1_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g639 ( .A(n_329), .Y(n_639) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g483 ( .A(n_330), .B(n_472), .Y(n_483) );
INVx1_ASAP7_75t_L g784 ( .A(n_330), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_330), .A2(n_637), .B1(n_832), .B2(n_849), .Y(n_869) );
BUFx2_ASAP7_75t_L g972 ( .A(n_330), .Y(n_972) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_330), .B(n_472), .Y(n_1387) );
INVx1_ASAP7_75t_L g973 ( .A(n_331), .Y(n_973) );
OAI221xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_336), .B1(n_337), .B2(n_340), .C(n_341), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g997 ( .A1(n_333), .A2(n_536), .B1(n_998), .B2(n_999), .C(n_1000), .Y(n_997) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
BUFx3_ASAP7_75t_L g534 ( .A(n_335), .Y(n_534) );
BUFx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g471 ( .A(n_338), .B(n_472), .Y(n_471) );
INVx8_ASAP7_75t_L g539 ( .A(n_338), .Y(n_539) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g629 ( .A(n_345), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g855 ( .A1(n_345), .A2(n_856), .B1(n_857), .B2(n_858), .C(n_859), .Y(n_855) );
INVx1_ASAP7_75t_L g901 ( .A(n_345), .Y(n_901) );
OAI221xp5_ASAP7_75t_L g962 ( .A1(n_345), .A2(n_541), .B1(n_856), .B2(n_963), .C(n_964), .Y(n_962) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_347), .A2(n_720), .B(n_736), .Y(n_719) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI31xp33_ASAP7_75t_L g851 ( .A1(n_349), .A2(n_852), .A3(n_860), .B(n_870), .Y(n_851) );
HB1xp67_ASAP7_75t_L g889 ( .A(n_349), .Y(n_889) );
OAI31xp33_ASAP7_75t_L g958 ( .A1(n_349), .A2(n_959), .A3(n_965), .B(n_974), .Y(n_958) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_349), .Y(n_1112) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AND3x4_ASAP7_75t_L g399 ( .A(n_350), .B(n_394), .C(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g424 ( .A(n_351), .Y(n_424) );
AOI21xp33_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_371), .B(n_372), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g1027 ( .A1(n_353), .A2(n_1028), .B(n_1029), .Y(n_1027) );
AOI21xp5_ASAP7_75t_L g1129 ( .A1(n_353), .A2(n_1130), .B(n_1131), .Y(n_1129) );
INVx8_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_367), .Y(n_354) );
INVx1_ASAP7_75t_L g620 ( .A(n_355), .Y(n_620) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_361), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_357), .Y(n_577) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx2_ASAP7_75t_L g518 ( .A(n_358), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_359), .Y(n_383) );
INVx2_ASAP7_75t_L g387 ( .A(n_359), .Y(n_387) );
AND2x4_ASAP7_75t_L g406 ( .A(n_359), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g445 ( .A(n_359), .B(n_389), .Y(n_445) );
INVx1_ASAP7_75t_L g382 ( .A(n_360), .Y(n_382) );
INVx2_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
OR2x2_ASAP7_75t_L g379 ( .A(n_361), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g447 ( .A(n_361), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_361), .Y(n_450) );
OR2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_365), .Y(n_361) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_362), .Y(n_524) );
INVx1_ASAP7_75t_L g557 ( .A(n_362), .Y(n_557) );
OR2x2_ASAP7_75t_L g563 ( .A(n_362), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g378 ( .A(n_363), .Y(n_378) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g811 ( .A(n_365), .Y(n_811) );
INVx3_ASAP7_75t_L g392 ( .A(n_366), .Y(n_392) );
BUFx3_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
NAND2xp33_ASAP7_75t_SL g564 ( .A(n_366), .B(n_394), .Y(n_564) );
INVx1_ASAP7_75t_L g750 ( .A(n_367), .Y(n_750) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
AND2x4_ASAP7_75t_L g435 ( .A(n_368), .B(n_391), .Y(n_435) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g589 ( .A(n_369), .Y(n_589) );
INVx2_ASAP7_75t_L g1097 ( .A(n_373), .Y(n_1097) );
AND2x4_ASAP7_75t_L g373 ( .A(n_374), .B(n_379), .Y(n_373) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_374), .B(n_379), .Y(n_1007) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_378), .Y(n_374) );
INVx1_ASAP7_75t_L g739 ( .A(n_375), .Y(n_739) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVxp67_ASAP7_75t_L g395 ( .A(n_378), .Y(n_395) );
INVx1_ASAP7_75t_L g460 ( .A(n_378), .Y(n_460) );
INVx1_ASAP7_75t_L g602 ( .A(n_378), .Y(n_602) );
INVx2_ASAP7_75t_L g622 ( .A(n_379), .Y(n_622) );
INVx4_ASAP7_75t_L g501 ( .A(n_380), .Y(n_501) );
INVx3_ASAP7_75t_L g824 ( .A(n_380), .Y(n_824) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_380), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g1364 ( .A(n_380), .Y(n_1364) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g571 ( .A(n_381), .Y(n_571) );
BUFx2_ASAP7_75t_L g1398 ( .A(n_381), .Y(n_1398) );
NAND2x1p5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
BUFx2_ASAP7_75t_L g512 ( .A(n_382), .Y(n_512) );
AND2x4_ASAP7_75t_L g415 ( .A(n_383), .B(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g434 ( .A(n_383), .Y(n_434) );
BUFx2_ASAP7_75t_L g508 ( .A(n_383), .Y(n_508) );
INVx3_ASAP7_75t_L g596 ( .A(n_384), .Y(n_596) );
INVx5_ASAP7_75t_L g882 ( .A(n_384), .Y(n_882) );
OR2x6_ASAP7_75t_L g384 ( .A(n_385), .B(n_395), .Y(n_384) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_386), .B(n_391), .Y(n_385) );
BUFx3_ASAP7_75t_L g404 ( .A(n_386), .Y(n_404) );
BUFx3_ASAP7_75t_L g671 ( .A(n_386), .Y(n_671) );
INVx8_ASAP7_75t_L g678 ( .A(n_386), .Y(n_678) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_386), .Y(n_802) );
AND2x4_ASAP7_75t_L g386 ( .A(n_387), .B(n_388), .Y(n_386) );
AND2x4_ASAP7_75t_L g411 ( .A(n_387), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVxp67_ASAP7_75t_L g412 ( .A(n_390), .Y(n_412) );
AND2x6_ASAP7_75t_L g791 ( .A(n_391), .B(n_433), .Y(n_791) );
AND2x2_ASAP7_75t_L g793 ( .A(n_391), .B(n_440), .Y(n_793) );
INVx1_ASAP7_75t_L g799 ( .A(n_391), .Y(n_799) );
AND2x4_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_392), .B(n_426), .Y(n_425) );
OR2x4_ASAP7_75t_L g495 ( .A(n_392), .B(n_445), .Y(n_495) );
INVx1_ASAP7_75t_L g498 ( .A(n_392), .Y(n_498) );
AND2x4_ASAP7_75t_L g503 ( .A(n_392), .B(n_406), .Y(n_503) );
OR2x6_ASAP7_75t_L g517 ( .A(n_392), .B(n_518), .Y(n_517) );
NAND3x1_ASAP7_75t_L g588 ( .A(n_392), .B(n_426), .C(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_394), .Y(n_522) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_441), .C(n_452), .Y(n_396) );
NAND2xp5_ASAP7_75t_SL g397 ( .A(n_398), .B(n_430), .Y(n_397) );
AOI33xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .A3(n_408), .B1(n_417), .B2(n_422), .B3(n_427), .Y(n_398) );
AOI33xp33_ASAP7_75t_L g837 ( .A1(n_399), .A2(n_422), .A3(n_838), .B1(n_840), .B2(n_841), .B3(n_844), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g940 ( .A(n_399), .B(n_941), .C(n_942), .Y(n_940) );
INVx3_ASAP7_75t_L g507 ( .A(n_400), .Y(n_507) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g706 ( .A(n_404), .Y(n_706) );
INVx1_ASAP7_75t_L g716 ( .A(n_404), .Y(n_716) );
BUFx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g429 ( .A(n_406), .Y(n_429) );
BUFx2_ASAP7_75t_L g455 ( .A(n_406), .Y(n_455) );
BUFx2_ASAP7_75t_L g672 ( .A(n_406), .Y(n_672) );
BUFx2_ASAP7_75t_L g695 ( .A(n_406), .Y(n_695) );
BUFx3_ASAP7_75t_L g797 ( .A(n_406), .Y(n_797) );
BUFx2_ASAP7_75t_L g922 ( .A(n_406), .Y(n_922) );
INVx1_ASAP7_75t_L g416 ( .A(n_407), .Y(n_416) );
INVx1_ASAP7_75t_L g1355 ( .A(n_409), .Y(n_1355) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g497 ( .A(n_410), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g662 ( .A(n_410), .Y(n_662) );
BUFx6f_ASAP7_75t_L g819 ( .A(n_410), .Y(n_819) );
INVx2_ASAP7_75t_L g1438 ( .A(n_410), .Y(n_1438) );
INVx1_ASAP7_75t_L g1446 ( .A(n_410), .Y(n_1446) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_411), .Y(n_420) );
BUFx8_ASAP7_75t_L g451 ( .A(n_411), .Y(n_451) );
INVx2_ASAP7_75t_L g575 ( .A(n_411), .Y(n_575) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx5_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx3_ASAP7_75t_L g421 ( .A(n_415), .Y(n_421) );
BUFx12f_ASAP7_75t_L g675 ( .A(n_415), .Y(n_675) );
BUFx3_ASAP7_75t_L g807 ( .A(n_415), .Y(n_807) );
INVx1_ASAP7_75t_L g440 ( .A(n_416), .Y(n_440) );
INVx8_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g1116 ( .A(n_419), .Y(n_1116) );
INVx5_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_420), .Y(n_580) );
INVx3_ASAP7_75t_L g804 ( .A(n_420), .Y(n_804) );
INVx2_ASAP7_75t_SL g843 ( .A(n_420), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_420), .A2(n_839), .B1(n_929), .B2(n_930), .Y(n_928) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_422), .B(n_950), .C(n_951), .Y(n_949) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OR2x6_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
AND2x4_ASAP7_75t_L g528 ( .A(n_424), .B(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g659 ( .A(n_424), .Y(n_659) );
INVx3_ASAP7_75t_L g816 ( .A(n_425), .Y(n_816) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g679 ( .A(n_429), .Y(n_679) );
INVx1_ASAP7_75t_L g707 ( .A(n_429), .Y(n_707) );
INVx2_ASAP7_75t_L g917 ( .A(n_429), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B1(n_436), .B2(n_437), .Y(n_430) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
AND2x4_ASAP7_75t_SL g615 ( .A(n_433), .B(n_435), .Y(n_615) );
NAND2x1_ASAP7_75t_L g1011 ( .A(n_433), .B(n_435), .Y(n_1011) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g437 ( .A(n_435), .B(n_438), .Y(n_437) );
AND2x4_ASAP7_75t_L g454 ( .A(n_435), .B(n_455), .Y(n_454) );
AND2x4_ASAP7_75t_SL g617 ( .A(n_435), .B(n_438), .Y(n_617) );
INVx1_ASAP7_75t_L g1012 ( .A(n_437), .Y(n_1012) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_437), .A2(n_454), .B1(n_615), .B2(n_1103), .C(n_1133), .Y(n_1132) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx2_ASAP7_75t_SL g584 ( .A(n_443), .Y(n_584) );
OR2x6_ASAP7_75t_L g603 ( .A(n_443), .B(n_446), .Y(n_603) );
OAI22xp33_ASAP7_75t_L g1036 ( .A1(n_443), .A2(n_823), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_443), .A2(n_1049), .B1(n_1050), .B2(n_1052), .Y(n_1048) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x4_ASAP7_75t_L g515 ( .A(n_445), .B(n_498), .Y(n_515) );
BUFx4f_ASAP7_75t_L g568 ( .A(n_445), .Y(n_568) );
BUFx3_ASAP7_75t_L g815 ( .A(n_445), .Y(n_815) );
BUFx3_ASAP7_75t_L g1122 ( .A(n_445), .Y(n_1122) );
INVxp67_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g607 ( .A(n_447), .B(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_449), .B(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_449), .B(n_944), .Y(n_943) );
AND2x4_ASAP7_75t_L g449 ( .A(n_450), .B(n_451), .Y(n_449) );
AND2x4_ASAP7_75t_L g833 ( .A(n_450), .B(n_834), .Y(n_833) );
AND2x4_ASAP7_75t_L g1136 ( .A(n_450), .B(n_834), .Y(n_1136) );
INVx2_ASAP7_75t_SL g1046 ( .A(n_451), .Y(n_1046) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
OAI211xp5_ASAP7_75t_SL g660 ( .A1(n_453), .A2(n_562), .B(n_661), .C(n_673), .Y(n_660) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_454), .A2(n_615), .B1(n_617), .B2(n_849), .C(n_850), .Y(n_848) );
AOI221xp5_ASAP7_75t_L g953 ( .A1(n_454), .A2(n_615), .B1(n_617), .B2(n_954), .C(n_955), .Y(n_953) );
HB1xp67_ASAP7_75t_L g1029 ( .A(n_454), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_461), .B1(n_491), .B2(n_519), .C(n_525), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx3_ASAP7_75t_L g1093 ( .A(n_459), .Y(n_1093) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_459), .Y(n_1430) );
NOR3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .C(n_476), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
HB1xp67_ASAP7_75t_L g1089 ( .A(n_465), .Y(n_1089) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_471), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_472), .B(n_732), .Y(n_1421) );
INVx3_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g1380 ( .A(n_475), .Y(n_1380) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g856 ( .A(n_478), .Y(n_856) );
INVx2_ASAP7_75t_L g1062 ( .A(n_478), .Y(n_1062) );
INVx4_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx4f_ASAP7_75t_L g545 ( .A(n_479), .Y(n_545) );
BUFx4f_ASAP7_75t_L g772 ( .A(n_479), .Y(n_772) );
OR2x6_ASAP7_75t_L g777 ( .A(n_479), .B(n_778), .Y(n_777) );
BUFx6f_ASAP7_75t_L g910 ( .A(n_479), .Y(n_910) );
BUFx4f_ASAP7_75t_L g1083 ( .A(n_479), .Y(n_1083) );
BUFx4f_ASAP7_75t_L g1385 ( .A(n_479), .Y(n_1385) );
BUFx6f_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx3_ASAP7_75t_L g551 ( .A(n_480), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B1(n_485), .B2(n_487), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g1084 ( .A1(n_482), .A2(n_1074), .B1(n_1085), .B2(n_1087), .Y(n_1084) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_484), .A2(n_505), .B1(n_509), .B2(n_510), .Y(n_504) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g1086 ( .A(n_486), .Y(n_1086) );
INVx2_ASAP7_75t_L g1390 ( .A(n_486), .Y(n_1390) );
NAND3xp33_ASAP7_75t_L g1418 ( .A(n_488), .B(n_1419), .C(n_1423), .Y(n_1418) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR3xp33_ASAP7_75t_L g491 ( .A(n_492), .B(n_499), .C(n_513), .Y(n_491) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_494), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g1069 ( .A(n_495), .Y(n_1069) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_497), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g1070 ( .A(n_497), .Y(n_1070) );
INVx2_ASAP7_75t_L g1394 ( .A(n_497), .Y(n_1394) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g814 ( .A(n_501), .Y(n_814) );
NAND4xp25_ASAP7_75t_L g685 ( .A(n_502), .B(n_686), .C(n_690), .D(n_696), .Y(n_685) );
NAND3xp33_ASAP7_75t_L g1455 ( .A(n_502), .B(n_1456), .C(n_1457), .Y(n_1455) );
CKINVDCx8_ASAP7_75t_R g502 ( .A(n_503), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g924 ( .A1(n_503), .A2(n_925), .A3(n_935), .B(n_936), .Y(n_924) );
CKINVDCx8_ASAP7_75t_R g1072 ( .A(n_503), .Y(n_1072) );
BUFx3_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx3_ASAP7_75t_L g692 ( .A(n_506), .Y(n_692) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
AND2x4_ASAP7_75t_L g511 ( .A(n_507), .B(n_512), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g925 ( .A1(n_507), .A2(n_926), .B(n_928), .C(n_931), .Y(n_925) );
AND2x4_ASAP7_75t_L g933 ( .A(n_507), .B(n_508), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g690 ( .A1(n_510), .A2(n_691), .B1(n_692), .B2(n_693), .C1(n_694), .C2(n_695), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_510), .A2(n_692), .B1(n_1388), .B2(n_1400), .Y(n_1399) );
AOI222xp33_ASAP7_75t_L g1456 ( .A1(n_510), .A2(n_692), .B1(n_717), .B2(n_1424), .C1(n_1425), .C2(n_1426), .Y(n_1456) );
BUFx6f_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g931 ( .A1(n_511), .A2(n_932), .B1(n_933), .B2(n_934), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_511), .A2(n_933), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_SL g699 ( .A(n_515), .Y(n_699) );
BUFx2_ASAP7_75t_L g1402 ( .A(n_515), .Y(n_1402) );
BUFx3_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g689 ( .A(n_517), .Y(n_689) );
INVx1_ASAP7_75t_L g666 ( .A(n_518), .Y(n_666) );
BUFx3_ASAP7_75t_L g1361 ( .A(n_518), .Y(n_1361) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_520), .A2(n_685), .B(n_700), .C(n_719), .Y(n_684) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_523), .Y(n_520) );
AND2x2_ASAP7_75t_L g936 ( .A(n_521), .B(n_523), .Y(n_936) );
AND2x2_ASAP7_75t_SL g1078 ( .A(n_521), .B(n_523), .Y(n_1078) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_561), .Y(n_525) );
OAI33xp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_530), .A3(n_540), .B1(n_547), .B2(n_553), .B3(n_558), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g766 ( .A(n_528), .Y(n_766) );
INVx2_ASAP7_75t_L g1055 ( .A(n_528), .Y(n_1055) );
INVx1_ASAP7_75t_L g1367 ( .A(n_528), .Y(n_1367) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B1(n_535), .B2(n_536), .Y(n_530) );
OAI22xp33_ASAP7_75t_L g565 ( .A1(n_531), .A2(n_548), .B1(n_566), .B2(n_569), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_532), .A2(n_536), .B1(n_559), .B2(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_534), .A2(n_761), .B1(n_762), .B2(n_764), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_535), .A2(n_552), .B1(n_583), .B2(n_585), .Y(n_582) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_538), .A2(n_876), .B1(n_877), .B2(n_879), .Y(n_875) );
INVx4_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g763 ( .A(n_539), .Y(n_763) );
INVx2_ASAP7_75t_L g968 ( .A(n_539), .Y(n_968) );
INVx1_ASAP7_75t_L g1060 ( .A(n_539), .Y(n_1060) );
BUFx6f_ASAP7_75t_L g1371 ( .A(n_539), .Y(n_1371) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B1(n_545), .B2(n_546), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_541), .A2(n_548), .B1(n_549), .B2(n_552), .Y(n_547) );
OAI22xp33_ASAP7_75t_SL g1063 ( .A1(n_541), .A2(n_1038), .B1(n_1052), .B2(n_1064), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_541), .A2(n_1083), .B1(n_1354), .B2(n_1358), .Y(n_1372) );
INVx1_ASAP7_75t_L g1375 ( .A(n_541), .Y(n_1375) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g859 ( .A(n_542), .Y(n_859) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g771 ( .A(n_543), .Y(n_771) );
BUFx3_ASAP7_75t_L g874 ( .A(n_543), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_544), .A2(n_559), .B1(n_573), .B2(n_576), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_546), .A2(n_560), .B1(n_579), .B2(n_581), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_549), .A2(n_647), .B(n_648), .C(n_651), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g1373 ( .A1(n_549), .A2(n_1351), .B1(n_1365), .B2(n_1374), .Y(n_1373) );
INVx5_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g728 ( .A(n_551), .Y(n_728) );
OR2x2_ASAP7_75t_L g755 ( .A(n_551), .B(n_754), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_551), .B(n_869), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_551), .B(n_971), .Y(n_970) );
OAI33xp33_ASAP7_75t_L g1053 ( .A1(n_553), .A2(n_1054), .A3(n_1056), .B1(n_1061), .B2(n_1063), .B3(n_1065), .Y(n_1053) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
OAI33xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .A3(n_572), .B1(n_578), .B2(n_582), .B3(n_586), .Y(n_561) );
BUFx4f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx4f_ASAP7_75t_L g709 ( .A(n_563), .Y(n_709) );
BUFx2_ASAP7_75t_L g1014 ( .A(n_563), .Y(n_1014) );
BUFx8_ASAP7_75t_L g1348 ( .A(n_563), .Y(n_1348) );
BUFx2_ASAP7_75t_L g826 ( .A(n_564), .Y(n_826) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g1352 ( .A(n_570), .Y(n_1352) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_571), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_573), .A2(n_702), .B1(n_703), .B2(n_704), .C(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g1023 ( .A(n_574), .Y(n_1023) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx3_ASAP7_75t_L g608 ( .A(n_575), .Y(n_608) );
BUFx2_ASAP7_75t_L g711 ( .A(n_575), .Y(n_711) );
BUFx2_ASAP7_75t_L g1041 ( .A(n_575), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g1022 ( .A1(n_576), .A2(n_1023), .B1(n_1024), .B2(n_1025), .C(n_1026), .Y(n_1022) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_576), .A2(n_1045), .B1(n_1046), .B2(n_1047), .Y(n_1044) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx3_ASAP7_75t_L g581 ( .A(n_577), .Y(n_581) );
CKINVDCx8_ASAP7_75t_R g703 ( .A(n_577), .Y(n_703) );
INVx3_ASAP7_75t_L g1043 ( .A(n_577), .Y(n_1043) );
INVx1_ASAP7_75t_L g1126 ( .A(n_577), .Y(n_1126) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_581), .A2(n_711), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_710) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_585), .A2(n_1119), .B1(n_1120), .B2(n_1123), .Y(n_1118) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_586), .A2(n_701), .B1(n_708), .B2(n_710), .Y(n_700) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g673 ( .A(n_587), .B(n_674), .C(n_676), .Y(n_673) );
INVx2_ASAP7_75t_L g923 ( .A(n_587), .Y(n_923) );
CKINVDCx5p33_ASAP7_75t_R g1443 ( .A(n_587), .Y(n_1443) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx3_ASAP7_75t_L g1021 ( .A(n_588), .Y(n_1021) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
XOR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_682), .Y(n_591) );
INVx1_ASAP7_75t_L g680 ( .A(n_593), .Y(n_680) );
NAND3xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .C(n_612), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_595), .A2(n_655), .B1(n_656), .B2(n_657), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_604), .B2(n_605), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_603), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_601), .A2(n_610), .B1(n_786), .B2(n_787), .Y(n_785) );
AND2x4_ASAP7_75t_L g610 ( .A(n_602), .B(n_611), .Y(n_610) );
NAND2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_609), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx2_ASAP7_75t_L g919 ( .A(n_608), .Y(n_919) );
INVx2_ASAP7_75t_L g1359 ( .A(n_608), .Y(n_1359) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g612 ( .A(n_613), .B(n_623), .C(n_660), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_619), .B(n_635), .Y(n_634) );
AOI222xp33_ASAP7_75t_L g831 ( .A1(n_620), .A2(n_622), .B1(n_832), .B2(n_833), .C1(n_835), .C2(n_836), .Y(n_831) );
AOI222xp33_ASAP7_75t_L g945 ( .A1(n_620), .A2(n_622), .B1(n_833), .B2(n_946), .C1(n_947), .C2(n_948), .Y(n_945) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_621), .A2(n_637), .B1(n_639), .B2(n_640), .C(n_641), .Y(n_636) );
AOI31xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_646), .A3(n_654), .B(n_658), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_630), .B(n_633), .Y(n_624) );
INVx2_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
BUFx2_ASAP7_75t_L g759 ( .A(n_628), .Y(n_759) );
AOI221xp5_ASAP7_75t_L g863 ( .A1(n_628), .A2(n_846), .B1(n_850), .B2(n_864), .C(n_866), .Y(n_863) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_628), .A2(n_864), .B1(n_944), .B2(n_955), .C(n_967), .Y(n_966) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .B(n_644), .Y(n_633) );
INVx1_ASAP7_75t_L g909 ( .A(n_637), .Y(n_909) );
AOI22xp5_ASAP7_75t_L g971 ( .A1(n_637), .A2(n_946), .B1(n_954), .B2(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g908 ( .A(n_639), .Y(n_908) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g867 ( .A1(n_645), .A2(n_732), .B(n_836), .C(n_868), .Y(n_867) );
A2O1A1Ixp33_ASAP7_75t_SL g904 ( .A1(n_645), .A2(n_905), .B(n_906), .C(n_907), .Y(n_904) );
INVx2_ASAP7_75t_L g723 ( .A(n_655), .Y(n_723) );
OAI31xp67_ASAP7_75t_L g788 ( .A1(n_658), .A2(n_789), .A3(n_800), .B(n_812), .Y(n_788) );
INVx1_ASAP7_75t_L g1003 ( .A(n_658), .Y(n_1003) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_663), .B1(n_664), .B2(n_667), .C(n_668), .Y(n_661) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g1017 ( .A(n_671), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_672), .A2(n_806), .B1(n_807), .B2(n_808), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_675), .A2(n_797), .B1(n_905), .B2(n_927), .Y(n_926) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g796 ( .A(n_678), .Y(n_796) );
INVx2_ASAP7_75t_L g834 ( .A(n_678), .Y(n_834) );
INVx8_ASAP7_75t_L g839 ( .A(n_678), .Y(n_839) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g1403 ( .A(n_689), .Y(n_1403) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_689), .A2(n_699), .B1(n_1420), .B2(n_1422), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_694), .B(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g718 ( .A(n_695), .Y(n_718) );
INVx2_ASAP7_75t_L g1077 ( .A(n_699), .Y(n_1077) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_703), .A2(n_818), .B1(n_820), .B2(n_821), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g912 ( .A1(n_703), .A2(n_913), .B1(n_914), .B2(n_915), .C(n_916), .Y(n_912) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_703), .A2(n_899), .B1(n_919), .B2(n_920), .C(n_921), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_703), .A2(n_1115), .B1(n_1116), .B2(n_1117), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1353 ( .A1(n_703), .A2(n_1354), .B1(n_1355), .B2(n_1356), .Y(n_1353) );
OAI22xp33_ASAP7_75t_L g911 ( .A1(n_708), .A2(n_912), .B1(n_918), .B2(n_923), .Y(n_911) );
OAI33xp33_ASAP7_75t_L g1035 ( .A1(n_708), .A2(n_1019), .A3(n_1036), .B1(n_1039), .B2(n_1044), .B3(n_1048), .Y(n_1035) );
OAI33xp33_ASAP7_75t_L g1432 ( .A1(n_708), .A2(n_1433), .A3(n_1436), .B1(n_1440), .B2(n_1443), .B3(n_1444), .Y(n_1432) );
BUFx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI211xp5_ASAP7_75t_SL g733 ( .A1(n_712), .A2(n_728), .B(n_734), .C(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g720 ( .A(n_721), .B(n_724), .Y(n_720) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B(n_729), .C(n_731), .Y(n_726) );
INVx3_ASAP7_75t_L g854 ( .A(n_732), .Y(n_854) );
BUFx6f_ASAP7_75t_L g906 ( .A(n_732), .Y(n_906) );
A2O1A1Ixp33_ASAP7_75t_L g969 ( .A1(n_732), .A2(n_948), .B(n_970), .C(n_973), .Y(n_969) );
INVx3_ASAP7_75t_SL g981 ( .A(n_741), .Y(n_981) );
BUFx3_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OA22x2_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_744), .B1(n_884), .B2(n_979), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
XOR2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_828), .Y(n_744) );
XNOR2x1_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
NAND4xp75_ASAP7_75t_L g747 ( .A(n_748), .B(n_756), .C(n_785), .D(n_788), .Y(n_747) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AOI211x1_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_765), .B(n_767), .C(n_781), .Y(n_756) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g813 ( .A1(n_764), .A2(n_773), .B1(n_814), .B2(n_815), .C(n_816), .Y(n_813) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI21xp5_ASAP7_75t_L g767 ( .A1(n_768), .A2(n_775), .B(n_777), .Y(n_767) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_770), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_768) );
OAI211xp5_ASAP7_75t_L g822 ( .A1(n_769), .A2(n_823), .B(n_825), .C(n_827), .Y(n_822) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
OAI211xp5_ASAP7_75t_SL g894 ( .A1(n_772), .A2(n_895), .B(n_896), .C(n_897), .Y(n_894) );
OAI211xp5_ASAP7_75t_SL g898 ( .A1(n_772), .A2(n_899), .B(n_900), .C(n_902), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g1448 ( .A1(n_775), .A2(n_1054), .B1(n_1449), .B2(n_1452), .Y(n_1448) );
CKINVDCx5p33_ASAP7_75t_R g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g1376 ( .A(n_776), .Y(n_1376) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NAND2x2_ASAP7_75t_L g782 ( .A(n_779), .B(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_786), .A2(n_787), .B1(n_802), .B2(n_803), .Y(n_801) );
INVx4_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
A2O1A1Ixp33_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_796), .B(n_797), .C(n_798), .Y(n_794) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AOI21xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_805), .B(n_809), .Y(n_800) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OAI21xp5_ASAP7_75t_SL g812 ( .A1(n_813), .A2(n_817), .B(n_822), .Y(n_812) );
OAI22xp33_ASAP7_75t_L g1349 ( .A1(n_815), .A2(n_1350), .B1(n_1351), .B2(n_1352), .Y(n_1349) );
OAI22xp33_ASAP7_75t_L g1362 ( .A1(n_815), .A2(n_1363), .B1(n_1364), .B2(n_1365), .Y(n_1362) );
OAI22xp33_ASAP7_75t_L g1433 ( .A1(n_815), .A2(n_1352), .B1(n_1434), .B2(n_1435), .Y(n_1433) );
OAI22xp33_ASAP7_75t_L g1440 ( .A1(n_815), .A2(n_1050), .B1(n_1441), .B2(n_1442), .Y(n_1440) );
OAI221xp5_ASAP7_75t_L g1124 ( .A1(n_818), .A2(n_1125), .B1(n_1126), .B2(n_1127), .C(n_1128), .Y(n_1124) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx2_ASAP7_75t_SL g913 ( .A(n_819), .Y(n_913) );
INVx2_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
XNOR2x1_ASAP7_75t_L g828 ( .A(n_829), .B(n_883), .Y(n_828) );
OR2x2_ASAP7_75t_L g829 ( .A(n_830), .B(n_847), .Y(n_829) );
NAND3xp33_ASAP7_75t_L g830 ( .A(n_831), .B(n_837), .C(n_845), .Y(n_830) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NAND3xp33_ASAP7_75t_SL g847 ( .A(n_848), .B(n_851), .C(n_880), .Y(n_847) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx2_ASAP7_75t_SL g991 ( .A(n_854), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_859), .A2(n_1040), .B1(n_1045), .B2(n_1062), .Y(n_1061) );
OAI221xp5_ASAP7_75t_SL g1449 ( .A1(n_859), .A2(n_1083), .B1(n_1437), .B2(n_1445), .C(n_1450), .Y(n_1449) );
OAI221xp5_ASAP7_75t_SL g1452 ( .A1(n_859), .A2(n_1083), .B1(n_1435), .B2(n_1442), .C(n_1453), .Y(n_1452) );
OAI21xp33_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_863), .B(n_867), .Y(n_860) );
OAI21xp5_ASAP7_75t_SL g965 ( .A1(n_861), .A2(n_966), .B(n_969), .Y(n_965) );
INVxp67_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g891 ( .A1(n_862), .A2(n_892), .B(n_893), .Y(n_891) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx4_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
BUFx6f_ASAP7_75t_L g1058 ( .A(n_878), .Y(n_1058) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_882), .B(n_957), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g1134 ( .A(n_882), .B(n_1111), .Y(n_1134) );
XNOR2xp5_ASAP7_75t_L g884 ( .A(n_885), .B(n_937), .Y(n_884) );
XOR2xp5_ASAP7_75t_L g979 ( .A(n_885), .B(n_937), .Y(n_979) );
XNOR2x1_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
AND2x2_ASAP7_75t_L g887 ( .A(n_888), .B(n_924), .Y(n_887) );
AOI21xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B(n_911), .Y(n_888) );
NAND4xp25_ASAP7_75t_L g890 ( .A(n_891), .B(n_894), .C(n_898), .D(n_904), .Y(n_890) );
HB1xp67_ASAP7_75t_L g1064 ( .A(n_910), .Y(n_1064) );
OAI33xp33_ASAP7_75t_L g1347 ( .A1(n_923), .A2(n_1348), .A3(n_1349), .B1(n_1353), .B2(n_1357), .B3(n_1362), .Y(n_1347) );
XNOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_978), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_939), .B(n_952), .Y(n_938) );
NAND4xp25_ASAP7_75t_SL g939 ( .A(n_940), .B(n_943), .C(n_945), .D(n_949), .Y(n_939) );
NAND3xp33_ASAP7_75t_SL g952 ( .A(n_953), .B(n_956), .C(n_958), .Y(n_952) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g982 ( .A1(n_983), .A2(n_1030), .B1(n_1138), .B2(n_1139), .Y(n_982) );
INVx1_ASAP7_75t_L g1138 ( .A(n_983), .Y(n_1138) );
BUFx2_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
O2A1O1Ixp5_ASAP7_75t_L g985 ( .A1(n_986), .A2(n_996), .B(n_1003), .C(n_1004), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g1015 ( .A1(n_998), .A2(n_1016), .B(n_1018), .Y(n_1015) );
NAND3xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1009), .C(n_1027), .Y(n_1004) );
NOR2xp33_ASAP7_75t_L g1005 ( .A(n_1006), .B(n_1008), .Y(n_1005) );
NOR2xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1013), .Y(n_1009) );
OAI22xp5_ASAP7_75t_SL g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1019), .B2(n_1022), .Y(n_1013) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
BUFx2_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1030), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
XNOR2xp5_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1094), .Y(n_1031) );
NAND3xp33_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1066), .C(n_1079), .Y(n_1033) );
NOR2xp33_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1053), .Y(n_1034) );
OAI22xp33_ASAP7_75t_L g1056 ( .A1(n_1037), .A2(n_1049), .B1(n_1057), .B2(n_1059), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1041), .B1(n_1042), .B2(n_1043), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_1042), .A2(n_1047), .B1(n_1057), .B2(n_1059), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1444 ( .A1(n_1043), .A2(n_1445), .B1(n_1446), .B2(n_1447), .Y(n_1444) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1057 ( .A(n_1058), .Y(n_1057) );
INVx2_ASAP7_75t_L g1369 ( .A(n_1058), .Y(n_1369) );
OAI22xp5_ASAP7_75t_L g1377 ( .A1(n_1059), .A2(n_1356), .B1(n_1360), .B2(n_1369), .Y(n_1377) );
BUFx3_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
OAI31xp33_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1071), .A3(n_1076), .B(n_1078), .Y(n_1066) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
OAI31xp33_ASAP7_75t_L g1392 ( .A1(n_1078), .A2(n_1393), .A3(n_1395), .B(n_1401), .Y(n_1392) );
OAI21xp33_ASAP7_75t_L g1454 ( .A1(n_1078), .A2(n_1455), .B(n_1458), .Y(n_1454) );
OAI31xp33_ASAP7_75t_SL g1079 ( .A1(n_1080), .A2(n_1082), .A3(n_1088), .B(n_1093), .Y(n_1079) );
INVx2_ASAP7_75t_L g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_1091), .A2(n_1420), .B1(n_1421), .B2(n_1422), .Y(n_1419) );
INVx2_ASAP7_75t_SL g1091 ( .A(n_1092), .Y(n_1091) );
OAI31xp33_ASAP7_75t_L g1378 ( .A1(n_1093), .A2(n_1379), .A3(n_1381), .B(n_1382), .Y(n_1378) );
XNOR2xp5_ASAP7_75t_L g1094 ( .A(n_1095), .B(n_1137), .Y(n_1094) );
NAND2xp5_ASAP7_75t_SL g1095 ( .A(n_1096), .B(n_1129), .Y(n_1095) );
AOI221xp5_ASAP7_75t_L g1096 ( .A1(n_1097), .A2(n_1098), .B1(n_1099), .B2(n_1112), .C(n_1113), .Y(n_1096) );
NAND3xp33_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1104), .C(n_1109), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1107), .B(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_1122), .Y(n_1121) );
NAND3xp33_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1134), .C(n_1135), .Y(n_1131) );
OAI221xp5_ASAP7_75t_L g1140 ( .A1(n_1141), .A2(n_1341), .B1(n_1344), .B2(n_1405), .C(n_1411), .Y(n_1140) );
NOR2xp67_ASAP7_75t_SL g1141 ( .A(n_1142), .B(n_1292), .Y(n_1141) );
OAI21xp5_ASAP7_75t_L g1142 ( .A1(n_1143), .A2(n_1239), .B(n_1247), .Y(n_1142) );
NOR4xp25_ASAP7_75t_L g1143 ( .A(n_1144), .B(n_1206), .C(n_1218), .D(n_1234), .Y(n_1143) );
OAI211xp5_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1161), .B(n_1179), .C(n_1194), .Y(n_1144) );
CKINVDCx14_ASAP7_75t_R g1145 ( .A(n_1146), .Y(n_1145) );
OAI322xp33_ASAP7_75t_L g1218 ( .A1(n_1146), .A2(n_1163), .A3(n_1219), .B1(n_1220), .B2(n_1225), .C1(n_1230), .C2(n_1232), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1259 ( .A1(n_1146), .A2(n_1172), .B1(n_1260), .B2(n_1261), .Y(n_1259) );
INVx3_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
OR2x2_ASAP7_75t_L g1188 ( .A(n_1147), .B(n_1189), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1147), .B(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1147), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1147), .B(n_1208), .Y(n_1255) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1147), .B(n_1200), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1147), .B(n_1190), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1147), .B(n_1189), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1147), .B(n_1200), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1147), .B(n_1190), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1148), .B(n_1155), .Y(n_1147) );
INVx2_ASAP7_75t_L g1244 ( .A(n_1149), .Y(n_1244) );
AND2x6_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1151), .Y(n_1149) );
AND2x2_ASAP7_75t_L g1153 ( .A(n_1150), .B(n_1154), .Y(n_1153) );
AND2x4_ASAP7_75t_L g1156 ( .A(n_1150), .B(n_1157), .Y(n_1156) );
AND2x6_ASAP7_75t_L g1159 ( .A(n_1150), .B(n_1160), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1150), .B(n_1154), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1150), .B(n_1154), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1152), .B(n_1158), .Y(n_1157) );
INVxp67_ASAP7_75t_L g1246 ( .A(n_1153), .Y(n_1246) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1159), .Y(n_1343) );
HB1xp67_ASAP7_75t_L g1465 ( .A(n_1160), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1167), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1182 ( .A(n_1162), .B(n_1176), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1162), .B(n_1215), .Y(n_1214) );
AND3x1_ASAP7_75t_L g1267 ( .A(n_1162), .B(n_1176), .C(n_1186), .Y(n_1267) );
NAND2xp5_ASAP7_75t_L g1275 ( .A(n_1162), .B(n_1186), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1162), .B(n_1168), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1162), .B(n_1306), .Y(n_1305) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
BUFx2_ASAP7_75t_L g1184 ( .A(n_1163), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1163), .B(n_1215), .Y(n_1231) );
OR2x2_ASAP7_75t_L g1237 ( .A(n_1163), .B(n_1238), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1163), .B(n_1172), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1163), .B(n_1306), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1168), .B(n_1172), .Y(n_1167) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1168), .Y(n_1197) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1168), .B(n_1228), .Y(n_1227) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1168), .B(n_1215), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1168), .B(n_1223), .Y(n_1301) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1169), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1169), .B(n_1181), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1169), .B(n_1200), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1169), .B(n_1200), .Y(n_1208) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1169), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1169), .B(n_1190), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1169), .B(n_1184), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1169), .B(n_1199), .Y(n_1317) );
NOR2xp33_ASAP7_75t_L g1329 ( .A(n_1169), .B(n_1209), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1332 ( .A(n_1169), .B(n_1333), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1172), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1327 ( .A(n_1172), .B(n_1285), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_1173), .B(n_1176), .Y(n_1172) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1173), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1173), .B(n_1216), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1333 ( .A(n_1173), .B(n_1184), .Y(n_1333) );
NAND3xp33_ASAP7_75t_L g1334 ( .A(n_1173), .B(n_1241), .C(n_1296), .Y(n_1334) );
OR2x2_ASAP7_75t_L g1173 ( .A(n_1174), .B(n_1175), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1176), .B(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1176), .Y(n_1216) );
OAI211xp5_ASAP7_75t_L g1258 ( .A1(n_1176), .A2(n_1204), .B(n_1259), .C(n_1263), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1176), .B(n_1317), .Y(n_1316) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1178), .Y(n_1176) );
OAI21xp5_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1183), .B(n_1187), .Y(n_1179) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
NOR2xp33_ASAP7_75t_L g1260 ( .A(n_1182), .B(n_1197), .Y(n_1260) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_1182), .A2(n_1237), .B1(n_1268), .B2(n_1314), .C(n_1315), .Y(n_1313) );
AOI21xp33_ASAP7_75t_L g1318 ( .A1(n_1182), .A2(n_1204), .B(n_1319), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1253 ( .A(n_1183), .B(n_1213), .Y(n_1253) );
NOR2xp33_ASAP7_75t_L g1299 ( .A(n_1183), .B(n_1214), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1185), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1184), .B(n_1186), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_1184), .B(n_1186), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1185), .B(n_1215), .Y(n_1219) );
NAND3xp33_ASAP7_75t_L g1225 ( .A(n_1185), .B(n_1226), .C(n_1229), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1185), .B(n_1285), .Y(n_1284) );
AOI221xp5_ASAP7_75t_L g1254 ( .A1(n_1186), .A2(n_1214), .B1(n_1255), .B2(n_1256), .C(n_1258), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1186), .B(n_1216), .Y(n_1306) );
AOI21xp5_ASAP7_75t_L g1315 ( .A1(n_1187), .A2(n_1316), .B(n_1318), .Y(n_1315) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1187), .B(n_1253), .Y(n_1320) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
NOR2xp33_ASAP7_75t_L g1203 ( .A(n_1189), .B(n_1204), .Y(n_1203) );
NOR2xp33_ASAP7_75t_SL g1221 ( .A(n_1189), .B(n_1222), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1189), .B(n_1199), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1189), .B(n_1241), .Y(n_1249) );
NAND2xp5_ASAP7_75t_L g1272 ( .A(n_1189), .B(n_1261), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1189), .B(n_1223), .Y(n_1325) );
CKINVDCx6p67_ASAP7_75t_R g1189 ( .A(n_1190), .Y(n_1189) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_1190), .Y(n_1217) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1190), .B(n_1236), .Y(n_1235) );
OR2x6_ASAP7_75t_L g1190 ( .A(n_1191), .B(n_1193), .Y(n_1190) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1191), .B(n_1193), .Y(n_1229) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1203), .B(n_1205), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1196 ( .A(n_1197), .B(n_1198), .Y(n_1196) );
CKINVDCx6p67_ASAP7_75t_R g1236 ( .A(n_1198), .Y(n_1236) );
INVx2_ASAP7_75t_L g1228 ( .A(n_1199), .Y(n_1228) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1223 ( .A(n_1200), .B(n_1224), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
CKINVDCx14_ASAP7_75t_R g1281 ( .A(n_1205), .Y(n_1281) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1205), .B(n_1301), .Y(n_1300) );
O2A1O1Ixp33_ASAP7_75t_L g1206 ( .A1(n_1207), .A2(n_1209), .B(n_1210), .C(n_1217), .Y(n_1206) );
AOI21xp33_ASAP7_75t_L g1338 ( .A1(n_1207), .A2(n_1339), .B(n_1340), .Y(n_1338) );
CKINVDCx14_ASAP7_75t_R g1207 ( .A(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1212), .B(n_1214), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1212), .B(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1212), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1212), .B(n_1261), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1212), .B(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1214), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1214), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1215), .B(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1215), .Y(n_1319) );
O2A1O1Ixp33_ASAP7_75t_L g1309 ( .A1(n_1217), .A2(n_1230), .B(n_1310), .C(n_1312), .Y(n_1309) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
AOI21xp33_ASAP7_75t_L g1302 ( .A1(n_1222), .A2(n_1303), .B(n_1304), .Y(n_1302) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_1223), .B(n_1278), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1226), .B(n_1231), .Y(n_1337) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1228), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1228), .B(n_1231), .Y(n_1308) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OAI21xp5_ASAP7_75t_SL g1273 ( .A1(n_1231), .A2(n_1274), .B(n_1276), .Y(n_1273) );
OAI22xp5_ASAP7_75t_L g1326 ( .A1(n_1232), .A2(n_1236), .B1(n_1327), .B2(n_1328), .Y(n_1326) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
NOR2xp33_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1237), .Y(n_1234) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_1236), .A2(n_1331), .B1(n_1332), .B2(n_1334), .Y(n_1330) );
OAI31xp33_ASAP7_75t_SL g1307 ( .A1(n_1239), .A2(n_1308), .A3(n_1309), .B(n_1313), .Y(n_1307) );
INVx3_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx2_ASAP7_75t_SL g1240 ( .A(n_1241), .Y(n_1240) );
INVx2_ASAP7_75t_SL g1282 ( .A(n_1241), .Y(n_1282) );
OAI22xp5_ASAP7_75t_SL g1242 ( .A1(n_1243), .A2(n_1244), .B1(n_1245), .B2(n_1246), .Y(n_1242) );
AOI211xp5_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1250), .B(n_1264), .C(n_1279), .Y(n_1247) );
INVx1_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
OAI21xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1252), .B(n_1254), .Y(n_1250) );
INVx2_ASAP7_75t_L g1257 ( .A(n_1251), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1251), .B(n_1269), .Y(n_1268) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_1251), .B(n_1289), .Y(n_1288) );
INVxp67_ASAP7_75t_L g1252 ( .A(n_1253), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1280 ( .A(n_1255), .Y(n_1280) );
INVx1_ASAP7_75t_L g1256 ( .A(n_1257), .Y(n_1256) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
OAI321xp33_ASAP7_75t_L g1279 ( .A1(n_1262), .A2(n_1280), .A3(n_1281), .B1(n_1282), .B2(n_1283), .C(n_1286), .Y(n_1279) );
OAI221xp5_ASAP7_75t_L g1264 ( .A1(n_1265), .A2(n_1268), .B1(n_1270), .B2(n_1272), .C(n_1273), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1269), .B(n_1296), .Y(n_1314) );
OAI21xp5_ASAP7_75t_L g1335 ( .A1(n_1269), .A2(n_1336), .B(n_1338), .Y(n_1335) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVxp67_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1288), .Y(n_1286) );
AOI211xp5_ASAP7_75t_L g1293 ( .A1(n_1287), .A2(n_1294), .B(n_1297), .C(n_1302), .Y(n_1293) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1287), .Y(n_1303) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1290), .Y(n_1289) );
NAND5xp2_ASAP7_75t_L g1292 ( .A(n_1293), .B(n_1307), .C(n_1320), .D(n_1321), .E(n_1335), .Y(n_1292) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
OAI21xp5_ASAP7_75t_L g1297 ( .A1(n_1298), .A2(n_1299), .B(n_1300), .Y(n_1297) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1305), .Y(n_1312) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NOR3xp33_ASAP7_75t_SL g1321 ( .A(n_1322), .B(n_1326), .C(n_1330), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1325), .Y(n_1323) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1324), .Y(n_1340) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVxp67_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
CKINVDCx20_ASAP7_75t_R g1341 ( .A(n_1342), .Y(n_1341) );
CKINVDCx20_ASAP7_75t_R g1342 ( .A(n_1343), .Y(n_1342) );
XOR2x2_ASAP7_75t_L g1344 ( .A(n_1345), .B(n_1404), .Y(n_1344) );
AND3x1_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1378), .C(n_1392), .Y(n_1345) );
NOR2xp33_ASAP7_75t_SL g1346 ( .A(n_1347), .B(n_1366), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g1368 ( .A1(n_1350), .A2(n_1363), .B1(n_1369), .B2(n_1370), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_1358), .A2(n_1359), .B1(n_1360), .B2(n_1361), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g1436 ( .A1(n_1361), .A2(n_1437), .B1(n_1438), .B2(n_1439), .Y(n_1436) );
OAI33xp33_ASAP7_75t_L g1366 ( .A1(n_1367), .A2(n_1368), .A3(n_1372), .B1(n_1373), .B2(n_1376), .B3(n_1377), .Y(n_1366) );
INVx6_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
AOI22xp33_ASAP7_75t_L g1386 ( .A1(n_1387), .A2(n_1388), .B1(n_1389), .B2(n_1391), .Y(n_1386) );
INVx2_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1390), .Y(n_1427) );
INVxp67_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
CKINVDCx20_ASAP7_75t_R g1405 ( .A(n_1406), .Y(n_1405) );
CKINVDCx20_ASAP7_75t_R g1406 ( .A(n_1407), .Y(n_1406) );
INVx3_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
BUFx3_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVxp33_ASAP7_75t_SL g1412 ( .A(n_1413), .Y(n_1412) );
INVxp67_ASAP7_75t_SL g1415 ( .A(n_1416), .Y(n_1415) );
NAND3x1_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1431), .C(n_1454), .Y(n_1416) );
OAI21xp5_ASAP7_75t_L g1417 ( .A1(n_1418), .A2(n_1428), .B(n_1430), .Y(n_1417) );
NOR2x1_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1448), .Y(n_1431) );
BUFx2_ASAP7_75t_SL g1459 ( .A(n_1460), .Y(n_1459) );
BUFx3_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx2_ASAP7_75t_SL g1462 ( .A(n_1463), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
OAI21xp5_ASAP7_75t_L g1464 ( .A1(n_1465), .A2(n_1466), .B(n_1467), .Y(n_1464) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
endmodule