module fake_aes_5249_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_2), .Y(n_11) );
INVxp67_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
CKINVDCx20_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
BUFx10_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_4), .B(n_5), .Y(n_16) );
OAI22xp5_ASAP7_75t_L g17 ( .A1(n_12), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_17) );
NOR2xp33_ASAP7_75t_R g18 ( .A(n_11), .B(n_10), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_16), .B(n_0), .C(n_1), .Y(n_19) );
OAI221xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_12), .B1(n_14), .B2(n_16), .C(n_15), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_17), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_20), .B(n_15), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_18), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_22), .B(n_15), .Y(n_24) );
AO21x1_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_17), .B(n_14), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
O2A1O1Ixp33_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_13), .B(n_15), .C(n_6), .Y(n_28) );
NAND4xp25_ASAP7_75t_L g29 ( .A(n_26), .B(n_3), .C(n_5), .D(n_7), .Y(n_29) );
CKINVDCx20_ASAP7_75t_R g30 ( .A(n_29), .Y(n_30) );
HB1xp67_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_31), .B(n_27), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_8), .B1(n_9), .B2(n_30), .C1(n_31), .C2(n_26), .Y(n_33) );
endmodule