module real_jpeg_4622_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_1),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_1),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_1),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_1),
.A2(n_112),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_1),
.A2(n_64),
.B1(n_145),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_2),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_2),
.A2(n_51),
.B1(n_66),
.B2(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_5),
.Y(n_69)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_5),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_5),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_5),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_5),
.B(n_9),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_78),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_6),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_7),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_8),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_9),
.A2(n_26),
.B1(n_78),
.B2(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_26),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_26),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_9),
.A2(n_204),
.B(n_205),
.C(n_209),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_29),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_9),
.B(n_242),
.C(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_9),
.B(n_168),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_9),
.B(n_105),
.C(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_9),
.B(n_122),
.Y(n_279)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_10),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_11),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_218),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_216),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_190),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_15),
.B(n_190),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_147),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_82),
.C(n_116),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_17),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_59),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_18),
.A2(n_19),
.B1(n_238),
.B2(n_246),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_18),
.B(n_246),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_18),
.A2(n_19),
.B1(n_166),
.B2(n_176),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_18),
.B(n_166),
.C(n_259),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_18),
.A2(n_19),
.B1(n_59),
.B2(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_19),
.Y(n_18)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_20),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_20),
.B(n_28),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_20),
.A2(n_28),
.B(n_53),
.Y(n_291)
);

INVx5_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_25),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_25),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_26),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_41),
.Y(n_28)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_39),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_53),
.Y(n_183)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_59),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_67),
.B(n_70),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_60),
.A2(n_154),
.B1(n_155),
.B2(n_160),
.Y(n_153)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_63),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_63),
.Y(n_245)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_71),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_71),
.A2(n_77),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_71),
.A2(n_77),
.B1(n_212),
.B2(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_76),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_77),
.B(n_186),
.Y(n_265)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_78),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_82),
.A2(n_116),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_110),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_99),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_84),
.A2(n_99),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B1(n_92),
.B2(n_95),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g262 ( 
.A(n_102),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_104),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_104),
.Y(n_173)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AO22x2_ASAP7_75t_L g166 ( 
.A1(n_110),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_166)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_110),
.Y(n_201)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_116),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_116),
.A2(n_193),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_121),
.B1(n_142),
.B2(n_146),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_117),
.A2(n_121),
.B1(n_142),
.B2(n_146),
.Y(n_165)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_132),
.Y(n_121)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_129),
.Y(n_122)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_124),
.Y(n_204)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_132)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_177),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_164),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_153),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_150),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_150),
.A2(n_197),
.B1(n_272),
.B2(n_273),
.Y(n_271)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_151),
.A2(n_152),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_154),
.B(n_187),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_175),
.B2(n_176),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_199),
.C(n_202),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_165),
.A2(n_175),
.B1(n_199),
.B2(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_166),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_166),
.A2(n_176),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_166),
.B(n_193),
.C(n_291),
.Y(n_309)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_185),
.B2(n_189),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_183),
.B(n_184),
.Y(n_179)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.C(n_198),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_191),
.B(n_195),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_197),
.B(n_211),
.C(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_197),
.B(n_272),
.C(n_274),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_198),
.B(n_301),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_199),
.A2(n_276),
.B1(n_277),
.B2(n_280),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_199),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_202),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_210),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_203),
.A2(n_210),
.B1(n_211),
.B2(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_203),
.Y(n_297)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_211),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_211),
.B(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_233),
.Y(n_234)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_299),
.B(n_315),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_284),
.B(n_298),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_269),
.B(n_283),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_256),
.B(n_268),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_248),
.B(n_255),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_235),
.B(n_247),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B(n_234),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_230),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_236),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_236),
.B(n_278),
.C(n_280),
.Y(n_294)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_249),
.B(n_254),
.Y(n_255)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_258),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_267),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_265),
.B2(n_266),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_266),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_282),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_282),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_274),
.B1(n_275),
.B2(n_281),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_292),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_294),
.C(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_302),
.B(n_310),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_302),
.C(n_316),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_306),
.C(n_308),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_308),
.B1(n_309),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);


endmodule