module real_jpeg_12717_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g90 ( 
.A(n_2),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_4),
.A2(n_66),
.B1(n_68),
.B2(n_73),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_73),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_6),
.A2(n_66),
.B1(n_68),
.B2(n_84),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_84),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_61),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_7),
.A2(n_61),
.B1(n_66),
.B2(n_68),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_61),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_12),
.A2(n_53),
.B1(n_66),
.B2(n_68),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_13),
.A2(n_35),
.B(n_36),
.C(n_41),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_13),
.B(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_13),
.A2(n_38),
.B1(n_41),
.B2(n_42),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_13),
.A2(n_38),
.B1(n_66),
.B2(n_68),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_13),
.A2(n_49),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_13),
.B(n_82),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_14),
.A2(n_66),
.B1(n_68),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_14),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_14),
.A2(n_24),
.B1(n_25),
.B2(n_93),
.Y(n_112)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_96),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_19),
.B(n_96),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_47),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_34),
.B1(n_45),
.B2(n_46),
.Y(n_21)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_23),
.B(n_51),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_23),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_23),
.A2(n_28),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_23),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_24),
.A2(n_25),
.B1(n_88),
.B2(n_89),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_24),
.B(n_38),
.C(n_89),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_24),
.B(n_145),
.Y(n_144)
);

CKINVDCx6p67_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_28),
.B(n_112),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_30),
.A2(n_49),
.B(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_35),
.A2(n_37),
.B1(n_41),
.B2(n_42),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B(n_39),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g109 ( 
.A(n_38),
.B(n_40),
.CON(n_109),
.SN(n_109)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_38),
.B(n_49),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_38),
.B(n_91),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_40),
.B1(n_65),
.B2(n_69),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_L g110 ( 
.A(n_39),
.B(n_66),
.C(n_69),
.Y(n_110)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_54),
.C(n_58),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_48),
.A2(n_54),
.B1(n_55),
.B2(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_49),
.B(n_52),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_49),
.A2(n_139),
.B1(n_147),
.B2(n_148),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_64),
.B2(n_71),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_63),
.B1(n_82),
.B2(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_72),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

OA22x2_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

O2A1O1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_68),
.B(n_108),
.C(n_110),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_68),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_68),
.B(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_80),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_92),
.B(n_94),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_103),
.B1(n_105),
.B2(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_105),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_86),
.A2(n_105),
.B1(n_124),
.B2(n_134),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_105),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_106),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_106),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_104),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_107),
.B(n_111),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_125),
.B(n_170),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_120),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.C(n_123),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_122),
.B(n_123),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_165),
.B(n_169),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_154),
.B(n_164),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_142),
.B(n_153),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_137),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_137),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_129)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_132),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_135),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_148),
.B(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_149),
.B(n_152),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_156),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_160),
.C(n_163),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_168),
.Y(n_169)
);


endmodule