module fake_jpeg_1852_n_211 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_211);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_211;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g67 ( 
.A(n_7),
.B(n_14),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_72),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_61),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_76),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_27),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_58),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_79),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_64),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_74),
.C(n_75),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_55),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_77),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_69),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_73),
.B(n_80),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_60),
.B(n_57),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_66),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_101),
.B(n_107),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_65),
.B1(n_58),
.B2(n_51),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_106),
.Y(n_128)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_81),
.B(n_62),
.CI(n_48),
.CON(n_107),
.SN(n_107)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_70),
.B1(n_53),
.B2(n_69),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_108),
.B1(n_54),
.B2(n_47),
.Y(n_135)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_108),
.A2(n_70),
.B1(n_69),
.B2(n_56),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_114),
.A2(n_121),
.B1(n_135),
.B2(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_116),
.B(n_124),
.Y(n_137)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_96),
.Y(n_136)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_119),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_123),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_50),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_60),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_133),
.Y(n_160)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_1),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_136),
.B(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_53),
.C(n_107),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_146),
.C(n_159),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_139),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_128),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_45),
.B1(n_31),
.B2(n_32),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_130),
.A2(n_52),
.B(n_2),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_12),
.B(n_18),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_29),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_147),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_52),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_126),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_2),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_132),
.B(n_3),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_134),
.B(n_3),
.Y(n_154)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_127),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_9),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_10),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_19),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_118),
.B(n_35),
.C(n_17),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_162),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_164),
.Y(n_180)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_155),
.A2(n_160),
.B(n_139),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_166),
.A2(n_170),
.B(n_41),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_169),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_149),
.B(n_157),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_26),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_20),
.C(n_22),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_174),
.B(n_177),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_23),
.C(n_25),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_178),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_181),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_182),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_170),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_185),
.A2(n_187),
.B1(n_177),
.B2(n_165),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_161),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_193),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_186),
.A2(n_175),
.B(n_168),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_161),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_172),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_184),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_197),
.A2(n_190),
.B1(n_176),
.B2(n_175),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_204),
.A2(n_198),
.B(n_188),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_189),
.B(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_207),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_205),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_189),
.C(n_43),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_42),
.Y(n_211)
);


endmodule