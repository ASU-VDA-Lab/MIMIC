module fake_netlist_6_4721_n_1235 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1235);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1235;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1061;
wire n_783;
wire n_798;
wire n_188;
wire n_509;
wire n_245;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1032;
wire n_893;
wire n_1099;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_836;
wire n_375;
wire n_522;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_224;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_530;
wire n_277;
wire n_618;
wire n_199;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_899;
wire n_189;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_272;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_184;
wire n_552;
wire n_216;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_958;
wire n_292;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_211;
wire n_231;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_217;
wire n_518;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_259;
wire n_177;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_238;
wire n_1095;
wire n_202;
wire n_597;
wire n_280;
wire n_1187;
wire n_610;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_183;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_218;
wire n_1213;
wire n_239;
wire n_782;
wire n_490;
wire n_809;
wire n_220;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_258;
wire n_456;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_273;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_569;
wire n_737;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_502;
wire n_672;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_855;
wire n_591;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_568;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_214;
wire n_246;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_911;
wire n_236;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_709;
wire n_366;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_257;
wire n_730;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_205;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_192;
wire n_649;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_30),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_54),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_83),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_100),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_8),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_8),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_3),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_49),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_162),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_171),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_21),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_141),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_5),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_144),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_156),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_44),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_80),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_76),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_88),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_45),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_97),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_90),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_114),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_94),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_150),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_154),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_11),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_168),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_103),
.Y(n_218)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_85),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_152),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_143),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_79),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_155),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_35),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_27),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_167),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_128),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_135),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_57),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_146),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_93),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_28),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_44),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_66),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_10),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_13),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_161),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_14),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_126),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_158),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_122),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_96),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_34),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_19),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_42),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_37),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_164),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_140),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_2),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_31),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_28),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g262 ( 
.A(n_91),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_33),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_7),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_1),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_15),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_111),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_62),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_70),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_21),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_110),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_78),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_14),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_133),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_47),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_142),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_6),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_92),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_149),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_0),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_48),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_165),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_68),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_65),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_137),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_153),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_29),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_16),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_169),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_151),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_148),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_131),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_184),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_264),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_215),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_226),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_259),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_211),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_187),
.Y(n_305)
);

BUFx6f_ASAP7_75t_SL g306 ( 
.A(n_190),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_228),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_203),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_1),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_191),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_231),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_244),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_254),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_200),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_216),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_223),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_261),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_263),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_173),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_232),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_224),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_267),
.B(n_2),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_275),
.B(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_236),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_235),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_240),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_173),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_237),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_203),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_252),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_174),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_219),
.B(n_4),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_174),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_253),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_270),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_273),
.B(n_4),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_219),
.B(n_5),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_277),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_266),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_257),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_287),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_271),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_258),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_286),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_229),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_178),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_199),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_201),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_205),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_213),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_202),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_206),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_181),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_212),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_222),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_181),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_207),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_275),
.B(n_6),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_208),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_238),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_248),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_182),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_250),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g369 ( 
.A(n_190),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

BUFx2_ASAP7_75t_L g371 ( 
.A(n_182),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_209),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_210),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_177),
.B(n_7),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_276),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_290),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_186),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_177),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_186),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_180),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_196),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_180),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_214),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_295),
.Y(n_384)
);

BUFx8_ASAP7_75t_L g385 ( 
.A(n_306),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_298),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_300),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_356),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_301),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_302),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_175),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_314),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

NAND2xp33_ASAP7_75t_SL g394 ( 
.A(n_343),
.B(n_196),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_305),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_175),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_382),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_353),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_333),
.B(n_241),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_185),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_310),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_316),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_360),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

NOR2x1_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_262),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_303),
.B(n_272),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_323),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_365),
.Y(n_412)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_322),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_368),
.B(n_179),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_370),
.B(n_179),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_329),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_376),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_347),
.B(n_183),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_374),
.A2(n_255),
.B(n_185),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_350),
.B(n_291),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_308),
.B(n_291),
.Y(n_424)
);

NOR2x1_ASAP7_75t_L g425 ( 
.A(n_357),
.B(n_176),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_331),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_334),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_308),
.B(n_176),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_340),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_297),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_381),
.B(n_255),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_336),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_355),
.B(n_190),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_325),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_297),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_326),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_362),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_299),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_294),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_309),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_361),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_299),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_369),
.B(n_183),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_304),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_349),
.A2(n_234),
.B1(n_260),
.B2(n_280),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_304),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_437),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_401),
.B(n_371),
.Y(n_456)
);

NAND3xp33_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_176),
.C(n_217),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_389),
.Y(n_458)
);

INVxp67_ASAP7_75t_SL g459 ( 
.A(n_431),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_390),
.Y(n_461)
);

CKINVDCx6p67_ASAP7_75t_R g462 ( 
.A(n_443),
.Y(n_462)
);

AO22x2_ASAP7_75t_L g463 ( 
.A1(n_437),
.A2(n_204),
.B1(n_265),
.B2(n_12),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_409),
.B(n_439),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_431),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_439),
.B(n_307),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_377),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_439),
.A2(n_371),
.B1(n_377),
.B2(n_176),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_413),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_421),
.A2(n_274),
.B(n_198),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_364),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_439),
.B(n_307),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

BUFx8_ASAP7_75t_SL g477 ( 
.A(n_446),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_418),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_386),
.Y(n_485)
);

AO22x2_ASAP7_75t_L g486 ( 
.A1(n_448),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_409),
.B(n_311),
.Y(n_487)
);

AND3x2_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_274),
.C(n_198),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_425),
.B(n_176),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_418),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_420),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_421),
.A2(n_274),
.B(n_198),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_439),
.A2(n_306),
.B1(n_320),
.B2(n_315),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_424),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_439),
.A2(n_281),
.B1(n_280),
.B2(n_330),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_425),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_431),
.B(n_311),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_388),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_445),
.B(n_312),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_431),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_400),
.Y(n_505)
);

OR2x6_ASAP7_75t_L g506 ( 
.A(n_445),
.B(n_58),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_386),
.Y(n_507)
);

OAI21xp33_ASAP7_75t_L g508 ( 
.A1(n_401),
.A2(n_281),
.B(n_335),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_384),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_384),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_424),
.B(n_312),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_384),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_424),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_386),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_386),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_399),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_423),
.B(n_313),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_445),
.B(n_59),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_400),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_404),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_391),
.B(n_313),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_60),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_386),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_386),
.Y(n_524)
);

INVx8_ASAP7_75t_L g525 ( 
.A(n_489),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_495),
.B(n_391),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_467),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_435),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_454),
.A2(n_422),
.B1(n_434),
.B2(n_433),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_495),
.B(n_513),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_465),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_455),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_513),
.B(n_435),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_459),
.B(n_445),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_465),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_480),
.B(n_435),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_454),
.A2(n_440),
.B1(n_435),
.B2(n_451),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_448),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_465),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_456),
.B(n_436),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_464),
.B(n_445),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_497),
.B(n_445),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_504),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_497),
.B(n_453),
.Y(n_544)
);

O2A1O1Ixp5_ASAP7_75t_L g545 ( 
.A1(n_466),
.A2(n_451),
.B(n_440),
.C(n_417),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_504),
.Y(n_546)
);

BUFx8_ASAP7_75t_L g547 ( 
.A(n_520),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_494),
.B(n_453),
.Y(n_548)
);

AND2x4_ASAP7_75t_SL g549 ( 
.A(n_462),
.B(n_453),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_456),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_504),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_501),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_455),
.Y(n_553)
);

NOR2x1p5_ASAP7_75t_L g554 ( 
.A(n_462),
.B(n_440),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_457),
.A2(n_422),
.B(n_450),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_457),
.A2(n_422),
.B(n_450),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_480),
.B(n_453),
.Y(n_557)
);

INVxp67_ASAP7_75t_SL g558 ( 
.A(n_507),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_480),
.B(n_453),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_511),
.B(n_517),
.Y(n_560)
);

OAI221xp5_ASAP7_75t_L g561 ( 
.A1(n_468),
.A2(n_434),
.B1(n_433),
.B2(n_397),
.C(n_415),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_470),
.B(n_453),
.Y(n_562)
);

BUFx8_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_480),
.B(n_440),
.Y(n_564)
);

INVxp67_ASAP7_75t_SL g565 ( 
.A(n_507),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_511),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_460),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_473),
.B(n_453),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_482),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_489),
.A2(n_422),
.B1(n_423),
.B2(n_436),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_470),
.B(n_441),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_460),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_461),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_474),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_SL g575 ( 
.A(n_474),
.B(n_441),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_482),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_455),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_517),
.B(n_436),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_475),
.B(n_444),
.Y(n_579)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_489),
.A2(n_423),
.B1(n_402),
.B2(n_444),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_475),
.B(n_404),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_476),
.B(n_447),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_461),
.B(n_447),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_516),
.A2(n_415),
.B(n_397),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_487),
.B(n_372),
.Y(n_585)
);

NOR2x1p5_ASAP7_75t_L g586 ( 
.A(n_500),
.B(n_294),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_458),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_476),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_508),
.B(n_423),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_458),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_503),
.A2(n_383),
.B1(n_373),
.B2(n_442),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_479),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_479),
.B(n_399),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_472),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_458),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_481),
.B(n_399),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_481),
.B(n_399),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_484),
.B(n_399),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

OR2x2_ASAP7_75t_SL g600 ( 
.A(n_488),
.B(n_414),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_496),
.B(n_414),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_478),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_478),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_490),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_490),
.B(n_491),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_508),
.B(n_442),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_482),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_399),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_493),
.B(n_399),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_469),
.B(n_320),
.C(n_315),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_493),
.B(n_407),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_498),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_471),
.B(n_335),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_471),
.B(n_296),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_SL g615 ( 
.A(n_498),
.B(n_499),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_471),
.B(n_337),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_499),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_489),
.B(n_407),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_478),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_509),
.B(n_407),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_489),
.B(n_407),
.Y(n_621)
);

A2O1A1Ixp33_ASAP7_75t_L g622 ( 
.A1(n_502),
.A2(n_505),
.B(n_519),
.C(n_408),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_570),
.B(n_509),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_533),
.A2(n_506),
.B1(n_518),
.B2(n_522),
.Y(n_624)
);

INVxp67_ASAP7_75t_SL g625 ( 
.A(n_530),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_555),
.A2(n_510),
.B(n_509),
.Y(n_626)
);

AO21x1_ASAP7_75t_L g627 ( 
.A1(n_548),
.A2(n_438),
.B(n_502),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_541),
.A2(n_514),
.B(n_506),
.Y(n_628)
);

INVx5_ASAP7_75t_L g629 ( 
.A(n_525),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_L g630 ( 
.A1(n_529),
.A2(n_506),
.B1(n_518),
.B2(n_522),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_539),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_534),
.A2(n_514),
.B(n_506),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_528),
.B(n_489),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_556),
.A2(n_512),
.B(n_510),
.Y(n_634)
);

NAND2x1_ASAP7_75t_L g635 ( 
.A(n_569),
.B(n_507),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_560),
.A2(n_348),
.B1(n_346),
.B2(n_293),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_539),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_554),
.B(n_506),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_526),
.B(n_489),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_525),
.A2(n_514),
.B(n_518),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_567),
.B(n_489),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_525),
.A2(n_514),
.B(n_518),
.Y(n_642)
);

AO21x1_ASAP7_75t_L g643 ( 
.A1(n_548),
.A2(n_519),
.B(n_505),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_540),
.B(n_443),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_525),
.A2(n_522),
.B(n_518),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_527),
.B(n_317),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_540),
.B(n_443),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_594),
.B(n_319),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_574),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_572),
.B(n_471),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_584),
.A2(n_522),
.B(n_515),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_562),
.A2(n_522),
.B(n_515),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_566),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_569),
.Y(n_654)
);

A2O1A1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_601),
.A2(n_452),
.B(n_396),
.C(n_430),
.Y(n_655)
);

CKINVDCx8_ASAP7_75t_R g656 ( 
.A(n_566),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_542),
.A2(n_523),
.B(n_515),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_569),
.Y(n_658)
);

OR2x6_ASAP7_75t_L g659 ( 
.A(n_560),
.B(n_463),
.Y(n_659)
);

AND2x2_ASAP7_75t_SL g660 ( 
.A(n_568),
.B(n_486),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_573),
.B(n_492),
.Y(n_661)
);

AOI21xp5_ASAP7_75t_L g662 ( 
.A1(n_542),
.A2(n_524),
.B(n_523),
.Y(n_662)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_537),
.A2(n_344),
.B1(n_332),
.B2(n_324),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_574),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_544),
.A2(n_565),
.B(n_558),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_544),
.A2(n_523),
.B(n_524),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_492),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_576),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_564),
.B(n_492),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_545),
.A2(n_512),
.B(n_510),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_578),
.B(n_492),
.Y(n_671)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_550),
.A2(n_328),
.B1(n_463),
.B2(n_486),
.Y(n_672)
);

OAI22xp5_ASAP7_75t_SL g673 ( 
.A1(n_606),
.A2(n_452),
.B1(n_296),
.B2(n_379),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_622),
.A2(n_512),
.B(n_524),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_588),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_592),
.Y(n_676)
);

AOI21x1_ASAP7_75t_L g677 ( 
.A1(n_615),
.A2(n_417),
.B(n_393),
.Y(n_677)
);

AOI33xp33_ASAP7_75t_L g678 ( 
.A1(n_578),
.A2(n_416),
.A3(n_426),
.B1(n_432),
.B2(n_419),
.B3(n_428),
.Y(n_678)
);

OAI21xp5_ASAP7_75t_L g679 ( 
.A1(n_622),
.A2(n_507),
.B(n_402),
.Y(n_679)
);

O2A1O1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_561),
.A2(n_419),
.B(n_396),
.C(n_432),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_583),
.B(n_321),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_539),
.B(n_407),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_L g683 ( 
.A(n_614),
.B(n_358),
.C(n_337),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_589),
.B(n_463),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_605),
.A2(n_402),
.B(n_406),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_589),
.A2(n_408),
.B(n_411),
.C(n_430),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_585),
.A2(n_407),
.B1(n_463),
.B2(n_402),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_582),
.B(n_463),
.Y(n_688)
);

AO21x1_ASAP7_75t_L g689 ( 
.A1(n_557),
.A2(n_486),
.B(n_393),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_618),
.A2(n_485),
.B(n_483),
.Y(n_690)
);

NOR2xp67_ASAP7_75t_L g691 ( 
.A(n_610),
.B(n_358),
.Y(n_691)
);

BUFx2_ASAP7_75t_L g692 ( 
.A(n_547),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_547),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_571),
.B(n_367),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_579),
.B(n_367),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_613),
.A2(n_411),
.B(n_429),
.C(n_428),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_621),
.A2(n_485),
.B(n_483),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_599),
.B(n_379),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_539),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_557),
.A2(n_486),
.B1(n_283),
.B2(n_282),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_538),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_538),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_576),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_604),
.B(n_407),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_612),
.B(n_406),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_559),
.A2(n_486),
.B1(n_282),
.B2(n_279),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_613),
.B(n_403),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_593),
.A2(n_485),
.B(n_483),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_552),
.B(n_403),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_617),
.B(n_406),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_531),
.B(n_412),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_SL g712 ( 
.A1(n_581),
.A2(n_429),
.B(n_426),
.C(n_416),
.Y(n_712)
);

AO21x1_ASAP7_75t_L g713 ( 
.A1(n_559),
.A2(n_393),
.B(n_392),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_616),
.A2(n_405),
.B1(n_392),
.B2(n_395),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_616),
.B(n_306),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_535),
.B(n_412),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_539),
.B(n_549),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_543),
.B(n_412),
.Y(n_718)
);

OAI21xp5_ASAP7_75t_L g719 ( 
.A1(n_667),
.A2(n_551),
.B(n_546),
.Y(n_719)
);

OAI22xp5_ASAP7_75t_L g720 ( 
.A1(n_630),
.A2(n_625),
.B1(n_624),
.B2(n_669),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_638),
.B(n_549),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_648),
.B(n_581),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_640),
.A2(n_580),
.B(n_596),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_SL g724 ( 
.A(n_655),
.B(n_189),
.C(n_188),
.Y(n_724)
);

AOI221xp5_ASAP7_75t_L g725 ( 
.A1(n_673),
.A2(n_591),
.B1(n_405),
.B2(n_192),
.C(n_194),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_655),
.A2(n_586),
.B(n_620),
.C(n_597),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_627),
.B(n_671),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_SL g728 ( 
.A(n_672),
.B(n_189),
.C(n_188),
.Y(n_728)
);

AOI21xp5_ASAP7_75t_L g729 ( 
.A1(n_642),
.A2(n_608),
.B(n_598),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_625),
.B(n_576),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_709),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_649),
.Y(n_732)
);

OR2x6_ASAP7_75t_L g733 ( 
.A(n_692),
.B(n_547),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_637),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_707),
.B(n_607),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_654),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_664),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_694),
.B(n_607),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_644),
.B(n_427),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_628),
.A2(n_632),
.B(n_651),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_647),
.B(n_427),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_637),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_658),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_629),
.A2(n_611),
.B(n_609),
.Y(n_744)
);

AOI22x1_ASAP7_75t_L g745 ( 
.A1(n_652),
.A2(n_553),
.B1(n_619),
.B2(n_577),
.Y(n_745)
);

OA21x2_ASAP7_75t_L g746 ( 
.A1(n_674),
.A2(n_620),
.B(n_553),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_629),
.A2(n_607),
.B(n_577),
.Y(n_747)
);

NOR2x1_ASAP7_75t_L g748 ( 
.A(n_683),
.B(n_532),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_SL g749 ( 
.A(n_663),
.B(n_194),
.C(n_192),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

INVx6_ASAP7_75t_L g751 ( 
.A(n_637),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_629),
.A2(n_590),
.B(n_587),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_695),
.B(n_575),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_701),
.B(n_427),
.Y(n_754)
);

OAI21xp5_ASAP7_75t_L g755 ( 
.A1(n_639),
.A2(n_590),
.B(n_587),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_615),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_648),
.B(n_600),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_668),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_681),
.B(n_575),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_645),
.B(n_595),
.Y(n_760)
);

INVxp67_ASAP7_75t_L g761 ( 
.A(n_701),
.Y(n_761)
);

INVx3_ASAP7_75t_SL g762 ( 
.A(n_659),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_687),
.A2(n_603),
.B(n_602),
.C(n_595),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_675),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_623),
.A2(n_602),
.B(n_485),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_SL g766 ( 
.A(n_656),
.B(n_477),
.Y(n_766)
);

BUFx2_ASAP7_75t_L g767 ( 
.A(n_653),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_646),
.B(n_600),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_703),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_714),
.B(n_395),
.Y(n_770)
);

BUFx2_ASAP7_75t_L g771 ( 
.A(n_702),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_714),
.B(n_563),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_623),
.A2(n_685),
.B(n_633),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_631),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_646),
.B(n_563),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_665),
.A2(n_483),
.B(n_485),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_676),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_696),
.A2(n_269),
.B(n_218),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_678),
.B(n_385),
.Y(n_779)
);

OAI21xp33_ASAP7_75t_L g780 ( 
.A1(n_702),
.A2(n_195),
.B(n_197),
.Y(n_780)
);

O2A1O1Ixp5_ASAP7_75t_L g781 ( 
.A1(n_643),
.A2(n_256),
.B(n_221),
.C(n_225),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_711),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_SL g783 ( 
.A(n_717),
.B(n_195),
.Y(n_783)
);

CKINVDCx8_ASAP7_75t_R g784 ( 
.A(n_767),
.Y(n_784)
);

OA21x2_ASAP7_75t_L g785 ( 
.A1(n_719),
.A2(n_740),
.B(n_727),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_721),
.B(n_631),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_723),
.A2(n_717),
.B(n_634),
.Y(n_787)
);

O2A1O1Ixp5_ASAP7_75t_SL g788 ( 
.A1(n_727),
.A2(n_700),
.B(n_706),
.C(n_650),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_771),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_722),
.B(n_715),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_722),
.A2(n_680),
.B(n_660),
.C(n_688),
.Y(n_791)
);

OAI21x1_ASAP7_75t_L g792 ( 
.A1(n_745),
.A2(n_670),
.B(n_662),
.Y(n_792)
);

OA21x2_ASAP7_75t_L g793 ( 
.A1(n_763),
.A2(n_626),
.B(n_686),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_731),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_732),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_732),
.Y(n_796)
);

OAI21x1_ASAP7_75t_L g797 ( 
.A1(n_729),
.A2(n_677),
.B(n_666),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_739),
.B(n_741),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_773),
.A2(n_661),
.B(n_641),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_720),
.A2(n_689),
.A3(n_713),
.B(n_686),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_777),
.Y(n_801)
);

CKINVDCx8_ASAP7_75t_R g802 ( 
.A(n_733),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_761),
.B(n_636),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_754),
.B(n_715),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_757),
.B(n_768),
.Y(n_805)
);

AOI221x1_ASAP7_75t_L g806 ( 
.A1(n_763),
.A2(n_768),
.B1(n_757),
.B2(n_778),
.C(n_684),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_775),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_721),
.B(n_638),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_777),
.Y(n_809)
);

AOI22xp5_ASAP7_75t_L g810 ( 
.A1(n_772),
.A2(n_691),
.B1(n_698),
.B2(n_693),
.Y(n_810)
);

O2A1O1Ixp5_ASAP7_75t_L g811 ( 
.A1(n_781),
.A2(n_682),
.B(n_679),
.C(n_657),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_759),
.A2(n_718),
.B(n_716),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_760),
.A2(n_682),
.B(n_704),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_764),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_782),
.B(n_659),
.Y(n_815)
);

NAND2x1_ASAP7_75t_L g816 ( 
.A(n_742),
.B(n_699),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_760),
.A2(n_708),
.B(n_690),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_750),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_750),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_750),
.Y(n_820)
);

AO31x2_ASAP7_75t_L g821 ( 
.A1(n_753),
.A2(n_710),
.A3(n_705),
.B(n_697),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_744),
.A2(n_699),
.B(n_635),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_730),
.A2(n_712),
.B(n_660),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_762),
.A2(n_659),
.B1(n_279),
.B2(n_278),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_737),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_775),
.B(n_197),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_735),
.B(n_712),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_766),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_750),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_738),
.A2(n_485),
.B(n_483),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_743),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_770),
.B(n_385),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_762),
.B(n_385),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_751),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_725),
.A2(n_385),
.B(n_283),
.C(n_284),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_728),
.A2(n_292),
.B(n_289),
.C(n_285),
.Y(n_836)
);

OAI21x1_ASAP7_75t_L g837 ( 
.A1(n_765),
.A2(n_485),
.B(n_483),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_780),
.B(n_724),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_743),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_790),
.B(n_749),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_SL g841 ( 
.A1(n_805),
.A2(n_733),
.B1(n_728),
.B2(n_724),
.Y(n_841)
);

CKINVDCx6p67_ASAP7_75t_R g842 ( 
.A(n_789),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_818),
.Y(n_843)
);

INVx6_ASAP7_75t_L g844 ( 
.A(n_807),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_806),
.A2(n_733),
.B1(n_779),
.B2(n_758),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_SL g846 ( 
.A1(n_826),
.A2(n_749),
.B1(n_278),
.B2(n_284),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_801),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_801),
.Y(n_848)
);

OAI22xp33_ASAP7_75t_L g849 ( 
.A1(n_798),
.A2(n_758),
.B1(n_736),
.B2(n_769),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_SL g850 ( 
.A1(n_803),
.A2(n_289),
.B1(n_285),
.B2(n_292),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_814),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_825),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_803),
.A2(n_838),
.B1(n_804),
.B2(n_832),
.Y(n_853)
);

BUFx8_ASAP7_75t_L g854 ( 
.A(n_789),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_809),
.Y(n_855)
);

INVx4_ASAP7_75t_L g856 ( 
.A(n_818),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_810),
.A2(n_748),
.B1(n_726),
.B2(n_756),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_794),
.A2(n_783),
.B1(n_774),
.B2(n_734),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_SL g859 ( 
.A1(n_807),
.A2(n_746),
.B1(n_756),
.B2(n_755),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_SL g860 ( 
.A1(n_807),
.A2(n_746),
.B1(n_230),
.B2(n_233),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_824),
.A2(n_746),
.B1(n_239),
.B2(n_242),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_791),
.A2(n_751),
.B1(n_742),
.B2(n_734),
.Y(n_862)
);

CKINVDCx11_ASAP7_75t_R g863 ( 
.A(n_784),
.Y(n_863)
);

INVx4_ASAP7_75t_L g864 ( 
.A(n_818),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_808),
.A2(n_774),
.B1(n_751),
.B2(n_220),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_828),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_818),
.Y(n_867)
);

AND2x4_ASAP7_75t_L g868 ( 
.A(n_808),
.B(n_774),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_834),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_SL g870 ( 
.A1(n_808),
.A2(n_833),
.B1(n_815),
.B2(n_796),
.Y(n_870)
);

BUFx4f_ASAP7_75t_L g871 ( 
.A(n_819),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_833),
.A2(n_245),
.B1(n_247),
.B2(n_249),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_795),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_819),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_819),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_795),
.B(n_774),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_831),
.Y(n_877)
);

OAI22x1_ASAP7_75t_SL g878 ( 
.A1(n_802),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_823),
.A2(n_752),
.B1(n_747),
.B2(n_776),
.Y(n_879)
);

BUFx8_ASAP7_75t_L g880 ( 
.A(n_834),
.Y(n_880)
);

AOI22xp33_ASAP7_75t_SL g881 ( 
.A1(n_793),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_820),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_820),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_819),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_839),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_829),
.Y(n_886)
);

INVx4_ASAP7_75t_L g887 ( 
.A(n_829),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_793),
.A2(n_20),
.B1(n_22),
.B2(n_23),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_829),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_SL g890 ( 
.A1(n_793),
.A2(n_785),
.B1(n_787),
.B2(n_827),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_829),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_836),
.B(n_23),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_786),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_786),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_816),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_812),
.A2(n_398),
.B1(n_387),
.B2(n_26),
.Y(n_896)
);

OAI21x1_ASAP7_75t_L g897 ( 
.A1(n_879),
.A2(n_817),
.B(n_797),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_853),
.B(n_785),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_883),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_873),
.Y(n_900)
);

OAI22xp33_ASAP7_75t_L g901 ( 
.A1(n_840),
.A2(n_785),
.B1(n_799),
.B2(n_813),
.Y(n_901)
);

OAI22xp33_ASAP7_75t_L g902 ( 
.A1(n_892),
.A2(n_836),
.B1(n_835),
.B2(n_788),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_844),
.Y(n_903)
);

INVx2_ASAP7_75t_SL g904 ( 
.A(n_844),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_863),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_855),
.Y(n_906)
);

OR2x2_ASAP7_75t_L g907 ( 
.A(n_890),
.B(n_800),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_885),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_844),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_851),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_852),
.Y(n_911)
);

OR2x6_ASAP7_75t_L g912 ( 
.A(n_857),
.B(n_797),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_870),
.B(n_821),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_877),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_847),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_890),
.B(n_800),
.Y(n_916)
);

OR2x2_ASAP7_75t_L g917 ( 
.A(n_845),
.B(n_800),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_848),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_L g919 ( 
.A1(n_850),
.A2(n_398),
.B1(n_792),
.B2(n_822),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_849),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_876),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_886),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_895),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_849),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_895),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_893),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_894),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_845),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_850),
.A2(n_398),
.B1(n_817),
.B2(n_387),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_859),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_859),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_875),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_862),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_930),
.B(n_881),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_929),
.A2(n_846),
.B1(n_841),
.B2(n_872),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_901),
.A2(n_830),
.B(n_837),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_902),
.A2(n_872),
.B(n_846),
.Y(n_937)
);

INVxp67_ASAP7_75t_L g938 ( 
.A(n_899),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_929),
.A2(n_860),
.B(n_896),
.Y(n_939)
);

NOR2x1_ASAP7_75t_SL g940 ( 
.A(n_912),
.B(n_875),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_908),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_921),
.B(n_882),
.Y(n_942)
);

OR2x2_ASAP7_75t_L g943 ( 
.A(n_907),
.B(n_821),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_930),
.B(n_931),
.Y(n_944)
);

OA21x2_ASAP7_75t_L g945 ( 
.A1(n_897),
.A2(n_811),
.B(n_858),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_907),
.B(n_869),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_931),
.B(n_881),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_902),
.A2(n_841),
.B1(n_878),
.B2(n_866),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_912),
.B(n_893),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_908),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_897),
.A2(n_843),
.B(n_867),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_913),
.B(n_888),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_928),
.A2(n_888),
.B1(n_861),
.B2(n_842),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_928),
.A2(n_861),
.B1(n_860),
.B2(n_865),
.Y(n_954)
);

OAI21x1_ASAP7_75t_L g955 ( 
.A1(n_897),
.A2(n_889),
.B(n_843),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_908),
.B(n_868),
.Y(n_956)
);

INVx3_ASAP7_75t_L g957 ( 
.A(n_923),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_913),
.B(n_868),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_913),
.B(n_867),
.Y(n_959)
);

NOR2x1_ASAP7_75t_SL g960 ( 
.A(n_912),
.B(n_875),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_905),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_913),
.B(n_874),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_899),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_910),
.B(n_874),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_900),
.B(n_889),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_906),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_900),
.Y(n_967)
);

OA21x2_ASAP7_75t_L g968 ( 
.A1(n_898),
.A2(n_875),
.B(n_891),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_912),
.B(n_894),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_910),
.B(n_894),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_933),
.A2(n_854),
.B1(n_880),
.B2(n_884),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_906),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_900),
.B(n_856),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_SL g974 ( 
.A(n_934),
.B(n_904),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_966),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_943),
.B(n_941),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_943),
.B(n_916),
.Y(n_977)
);

OR2x6_ASAP7_75t_SL g978 ( 
.A(n_953),
.B(n_917),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_967),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_966),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_941),
.B(n_912),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_950),
.B(n_912),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_968),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_946),
.B(n_916),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_972),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_967),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_972),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_946),
.B(n_917),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_968),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_950),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_963),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_963),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_957),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_957),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_957),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_951),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_968),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_952),
.B(n_919),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_964),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_991),
.Y(n_1000)
);

OAI222xp33_ASAP7_75t_L g1001 ( 
.A1(n_978),
.A2(n_948),
.B1(n_935),
.B2(n_954),
.C1(n_939),
.C2(n_934),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_976),
.B(n_940),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_990),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_976),
.B(n_938),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_986),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_986),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_976),
.B(n_940),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_991),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_992),
.B(n_944),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_990),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_986),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_977),
.B(n_968),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_992),
.B(n_944),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_R g1014 ( 
.A(n_978),
.B(n_961),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_989),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_SL g1016 ( 
.A1(n_978),
.A2(n_937),
.B(n_971),
.Y(n_1016)
);

AOI33xp33_ASAP7_75t_L g1017 ( 
.A1(n_999),
.A2(n_947),
.A3(n_952),
.B1(n_970),
.B2(n_964),
.B3(n_911),
.Y(n_1017)
);

OAI31xp33_ASAP7_75t_L g1018 ( 
.A1(n_998),
.A2(n_947),
.A3(n_933),
.B(n_942),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_986),
.Y(n_1019)
);

OR2x2_ASAP7_75t_L g1020 ( 
.A(n_977),
.B(n_949),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_990),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1002),
.B(n_981),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_1003),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1002),
.B(n_981),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1003),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_1007),
.B(n_1015),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1007),
.B(n_981),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_1015),
.B(n_982),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_1012),
.B(n_977),
.Y(n_1029)
);

NOR2x1_ASAP7_75t_L g1030 ( 
.A(n_1016),
.B(n_989),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_1010),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1015),
.B(n_982),
.Y(n_1032)
);

INVx3_ASAP7_75t_R g1033 ( 
.A(n_1014),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1030),
.B(n_989),
.Y(n_1034)
);

AND2x2_ASAP7_75t_SL g1035 ( 
.A(n_1033),
.B(n_998),
.Y(n_1035)
);

OR2x2_ASAP7_75t_L g1036 ( 
.A(n_1029),
.B(n_1012),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_1026),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1023),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1022),
.B(n_1024),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_1029),
.B(n_1009),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1023),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1035),
.B(n_1016),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1038),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_1037),
.B(n_1026),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1037),
.B(n_1026),
.Y(n_1045)
);

OR2x2_ASAP7_75t_L g1046 ( 
.A(n_1040),
.B(n_1020),
.Y(n_1046)
);

OAI211xp5_ASAP7_75t_L g1047 ( 
.A1(n_1042),
.A2(n_1018),
.B(n_1035),
.C(n_1037),
.Y(n_1047)
);

AOI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_1044),
.A2(n_1034),
.B1(n_998),
.B2(n_1039),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1044),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_SL g1050 ( 
.A(n_1045),
.B(n_1014),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1045),
.B(n_1039),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_1022),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1043),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_1046),
.B(n_1033),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1043),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1043),
.Y(n_1056)
);

OAI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_1042),
.A2(n_1001),
.B1(n_1018),
.B2(n_1034),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1053),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_1054),
.B(n_1034),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1049),
.B(n_1024),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1057),
.A2(n_1001),
.B(n_1038),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1057),
.B(n_961),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1053),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1056),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_1049),
.B(n_1027),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1048),
.A2(n_998),
.B1(n_1040),
.B2(n_1020),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1054),
.B(n_1027),
.Y(n_1067)
);

AOI222xp33_ASAP7_75t_L g1068 ( 
.A1(n_1047),
.A2(n_983),
.B1(n_989),
.B2(n_1000),
.C1(n_1008),
.C2(n_1015),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_1050),
.A2(n_1041),
.B(n_1008),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1051),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1055),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_1052),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1057),
.A2(n_949),
.B1(n_1041),
.B2(n_969),
.Y(n_1073)
);

NAND4xp25_ASAP7_75t_L g1074 ( 
.A(n_1062),
.B(n_1017),
.C(n_1036),
.D(n_1028),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1061),
.A2(n_1036),
.B(n_1000),
.C(n_997),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1068),
.A2(n_983),
.B1(n_997),
.B2(n_854),
.Y(n_1076)
);

AOI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1066),
.A2(n_983),
.B(n_1032),
.C(n_1028),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_L g1078 ( 
.A1(n_1067),
.A2(n_1032),
.B(n_1004),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_1069),
.B(n_1009),
.Y(n_1079)
);

INVx3_ASAP7_75t_SL g1080 ( 
.A(n_1059),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1070),
.B(n_1025),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1059),
.Y(n_1082)
);

O2A1O1Ixp33_ASAP7_75t_L g1083 ( 
.A1(n_1064),
.A2(n_1013),
.B(n_1004),
.C(n_1025),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_1059),
.B(n_1031),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1058),
.Y(n_1085)
);

XNOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1072),
.B(n_24),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1063),
.Y(n_1087)
);

O2A1O1Ixp5_ASAP7_75t_SL g1088 ( 
.A1(n_1071),
.A2(n_1031),
.B(n_1021),
.C(n_1010),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_1060),
.B(n_903),
.C(n_909),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_1073),
.A2(n_1013),
.B(n_919),
.C(n_901),
.Y(n_1090)
);

AOI211xp5_ASAP7_75t_L g1091 ( 
.A1(n_1065),
.A2(n_904),
.B(n_903),
.C(n_984),
.Y(n_1091)
);

AOI222xp33_ASAP7_75t_L g1092 ( 
.A1(n_1062),
.A2(n_960),
.B1(n_898),
.B2(n_982),
.C1(n_970),
.C2(n_924),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1085),
.Y(n_1093)
);

NOR3xp33_ASAP7_75t_L g1094 ( 
.A(n_1082),
.B(n_1075),
.C(n_1087),
.Y(n_1094)
);

OAI221xp5_ASAP7_75t_L g1095 ( 
.A1(n_1080),
.A2(n_904),
.B1(n_903),
.B2(n_949),
.C(n_984),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1086),
.B(n_880),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1084),
.B(n_1005),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1081),
.B(n_1005),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1078),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1083),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_SL g1101 ( 
.A(n_1076),
.B(n_24),
.C(n_25),
.Y(n_1101)
);

NAND3xp33_ASAP7_75t_SL g1102 ( 
.A(n_1076),
.B(n_984),
.C(n_909),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1079),
.B(n_1005),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1077),
.B(n_1006),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_1074),
.B(n_1006),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1091),
.Y(n_1106)
);

NAND4xp75_ASAP7_75t_L g1107 ( 
.A(n_1089),
.B(n_25),
.C(n_26),
.D(n_27),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1090),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1092),
.Y(n_1109)
);

AOI211xp5_ASAP7_75t_L g1110 ( 
.A1(n_1101),
.A2(n_1088),
.B(n_30),
.C(n_31),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1096),
.B(n_29),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1099),
.A2(n_903),
.B1(n_909),
.B2(n_949),
.Y(n_1112)
);

NAND4xp75_ASAP7_75t_L g1113 ( 
.A(n_1093),
.B(n_32),
.C(n_35),
.D(n_36),
.Y(n_1113)
);

OAI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1101),
.A2(n_909),
.B(n_37),
.C(n_38),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1094),
.B(n_1006),
.Y(n_1115)
);

OAI32xp33_ASAP7_75t_L g1116 ( 
.A1(n_1100),
.A2(n_1019),
.A3(n_1011),
.B1(n_988),
.B2(n_996),
.Y(n_1116)
);

NAND2xp33_ASAP7_75t_R g1117 ( 
.A(n_1108),
.B(n_32),
.Y(n_1117)
);

NAND4xp25_ASAP7_75t_L g1118 ( 
.A(n_1109),
.B(n_988),
.C(n_959),
.D(n_962),
.Y(n_1118)
);

NAND4xp75_ASAP7_75t_L g1119 ( 
.A(n_1106),
.B(n_38),
.C(n_39),
.D(n_40),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_1105),
.B(n_927),
.C(n_864),
.Y(n_1120)
);

OAI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_1095),
.A2(n_949),
.B1(n_969),
.B2(n_1021),
.C(n_988),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1097),
.Y(n_1122)
);

OAI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1102),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_1107),
.B(n_41),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1098),
.Y(n_1125)
);

NOR2x1_ASAP7_75t_L g1126 ( 
.A(n_1103),
.B(n_42),
.Y(n_1126)
);

OAI221xp5_ASAP7_75t_L g1127 ( 
.A1(n_1104),
.A2(n_969),
.B1(n_1011),
.B2(n_1019),
.C(n_996),
.Y(n_1127)
);

OAI211xp5_ASAP7_75t_L g1128 ( 
.A1(n_1101),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1096),
.B(n_46),
.Y(n_1129)
);

NAND4xp25_ASAP7_75t_L g1130 ( 
.A(n_1099),
.B(n_959),
.C(n_962),
.D(n_911),
.Y(n_1130)
);

INVx2_ASAP7_75t_SL g1131 ( 
.A(n_1093),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1094),
.B(n_1019),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_L g1133 ( 
.A(n_1094),
.B(n_927),
.C(n_864),
.Y(n_1133)
);

NAND4xp25_ASAP7_75t_SL g1134 ( 
.A(n_1110),
.B(n_1011),
.C(n_932),
.D(n_974),
.Y(n_1134)
);

OAI211xp5_ASAP7_75t_L g1135 ( 
.A1(n_1114),
.A2(n_1128),
.B(n_1123),
.C(n_1124),
.Y(n_1135)
);

NAND2x1p5_ASAP7_75t_L g1136 ( 
.A(n_1126),
.B(n_871),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1133),
.A2(n_996),
.B1(n_969),
.B2(n_999),
.Y(n_1137)
);

AOI221xp5_ASAP7_75t_L g1138 ( 
.A1(n_1120),
.A2(n_974),
.B1(n_927),
.B2(n_922),
.C(n_987),
.Y(n_1138)
);

OAI221xp5_ASAP7_75t_SL g1139 ( 
.A1(n_1112),
.A2(n_1132),
.B1(n_1115),
.B2(n_1118),
.C(n_1131),
.Y(n_1139)
);

AOI31xp33_ASAP7_75t_L g1140 ( 
.A1(n_1117),
.A2(n_932),
.A3(n_974),
.B(n_49),
.Y(n_1140)
);

AOI221xp5_ASAP7_75t_L g1141 ( 
.A1(n_1122),
.A2(n_974),
.B1(n_927),
.B2(n_922),
.C(n_987),
.Y(n_1141)
);

AOI211xp5_ASAP7_75t_L g1142 ( 
.A1(n_1111),
.A2(n_47),
.B(n_48),
.C(n_50),
.Y(n_1142)
);

AOI321xp33_ASAP7_75t_L g1143 ( 
.A1(n_1125),
.A2(n_51),
.A3(n_52),
.B1(n_53),
.B2(n_54),
.C(n_55),
.Y(n_1143)
);

NAND2x1p5_ASAP7_75t_L g1144 ( 
.A(n_1129),
.B(n_871),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1121),
.A2(n_1127),
.B1(n_1130),
.B2(n_1119),
.Y(n_1145)
);

NAND4xp75_ASAP7_75t_L g1146 ( 
.A(n_1113),
.B(n_51),
.C(n_52),
.D(n_53),
.Y(n_1146)
);

NOR3xp33_ASAP7_75t_L g1147 ( 
.A(n_1116),
.B(n_856),
.C(n_884),
.Y(n_1147)
);

OAI211xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1110),
.A2(n_55),
.B(n_56),
.C(n_914),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_L g1149 ( 
.A(n_1114),
.B(n_887),
.C(n_926),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1126),
.Y(n_1150)
);

NAND5xp2_ASAP7_75t_L g1151 ( 
.A(n_1110),
.B(n_56),
.C(n_924),
.D(n_920),
.E(n_914),
.Y(n_1151)
);

AO22x1_ASAP7_75t_L g1152 ( 
.A1(n_1126),
.A2(n_887),
.B1(n_932),
.B2(n_926),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_L g1153 ( 
.A(n_1114),
.B(n_926),
.C(n_922),
.Y(n_1153)
);

AOI222xp33_ASAP7_75t_L g1154 ( 
.A1(n_1115),
.A2(n_960),
.B1(n_920),
.B2(n_975),
.C1(n_980),
.C2(n_985),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1117),
.A2(n_969),
.B1(n_927),
.B2(n_962),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1126),
.Y(n_1156)
);

OAI211xp5_ASAP7_75t_L g1157 ( 
.A1(n_1114),
.A2(n_926),
.B(n_927),
.C(n_975),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1134),
.A2(n_927),
.B1(n_962),
.B2(n_993),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1136),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1150),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1155),
.A2(n_1139),
.B1(n_1156),
.B2(n_1140),
.Y(n_1161)
);

AO22x2_ASAP7_75t_L g1162 ( 
.A1(n_1146),
.A2(n_995),
.B1(n_994),
.B2(n_993),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1135),
.B(n_921),
.Y(n_1163)
);

NOR2x1_ASAP7_75t_L g1164 ( 
.A(n_1148),
.B(n_980),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1143),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1151),
.B(n_985),
.Y(n_1166)
);

NOR2x1p5_ASAP7_75t_L g1167 ( 
.A(n_1149),
.B(n_986),
.Y(n_1167)
);

XNOR2xp5_ASAP7_75t_L g1168 ( 
.A(n_1142),
.B(n_61),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_1157),
.B(n_979),
.Y(n_1169)
);

XNOR2xp5_ASAP7_75t_L g1170 ( 
.A(n_1144),
.B(n_63),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1145),
.A2(n_923),
.B(n_925),
.C(n_995),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_1153),
.B(n_958),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_1137),
.B(n_398),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1152),
.Y(n_1174)
);

NOR3xp33_ASAP7_75t_L g1175 ( 
.A(n_1147),
.B(n_921),
.C(n_918),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1154),
.Y(n_1176)
);

NOR3xp33_ASAP7_75t_L g1177 ( 
.A(n_1138),
.B(n_918),
.C(n_923),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1141),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1150),
.B(n_958),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1162),
.Y(n_1180)
);

AND3x1_ASAP7_75t_L g1181 ( 
.A(n_1165),
.B(n_994),
.C(n_979),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1160),
.B(n_979),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_1179),
.B(n_891),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1159),
.B(n_965),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1161),
.B(n_398),
.C(n_925),
.Y(n_1185)
);

AND2x4_ASAP7_75t_L g1186 ( 
.A(n_1167),
.B(n_958),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1166),
.B(n_64),
.Y(n_1187)
);

NOR3xp33_ASAP7_75t_L g1188 ( 
.A(n_1171),
.B(n_955),
.C(n_951),
.Y(n_1188)
);

AND2x2_ASAP7_75t_SL g1189 ( 
.A(n_1174),
.B(n_973),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1176),
.A2(n_973),
.B1(n_965),
.B2(n_925),
.C(n_958),
.Y(n_1190)
);

OAI211xp5_ASAP7_75t_L g1191 ( 
.A1(n_1163),
.A2(n_945),
.B(n_69),
.C(n_71),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1164),
.B(n_973),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_L g1193 ( 
.A(n_1168),
.B(n_398),
.C(n_973),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_1170),
.B(n_67),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1180),
.Y(n_1195)
);

XNOR2x1_ASAP7_75t_L g1196 ( 
.A(n_1193),
.B(n_1162),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1189),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1187),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_SL g1199 ( 
.A1(n_1185),
.A2(n_1178),
.B1(n_1173),
.B2(n_1172),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1194),
.B(n_1175),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1182),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1181),
.Y(n_1202)
);

AOI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1190),
.A2(n_1177),
.B1(n_1169),
.B2(n_1158),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1184),
.A2(n_965),
.B1(n_956),
.B2(n_945),
.Y(n_1204)
);

NAND4xp25_ASAP7_75t_L g1205 ( 
.A(n_1183),
.B(n_956),
.C(n_965),
.D(n_74),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1192),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1186),
.B(n_956),
.Y(n_1207)
);

BUFx2_ASAP7_75t_L g1208 ( 
.A(n_1191),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1188),
.B(n_956),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1206),
.A2(n_945),
.B1(n_936),
.B2(n_955),
.Y(n_1210)
);

NAND4xp25_ASAP7_75t_L g1211 ( 
.A(n_1208),
.B(n_72),
.C(n_73),
.D(n_75),
.Y(n_1211)
);

NAND4xp25_ASAP7_75t_L g1212 ( 
.A(n_1200),
.B(n_77),
.C(n_81),
.D(n_82),
.Y(n_1212)
);

HB1xp67_ASAP7_75t_L g1213 ( 
.A(n_1202),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1197),
.Y(n_1214)
);

XNOR2x1_ASAP7_75t_L g1215 ( 
.A(n_1196),
.B(n_86),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1195),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1198),
.A2(n_945),
.B1(n_936),
.B2(n_915),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1199),
.A2(n_936),
.B1(n_915),
.B2(n_387),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_1201),
.A2(n_915),
.B1(n_95),
.B2(n_101),
.Y(n_1219)
);

AOI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1214),
.A2(n_1205),
.B1(n_1203),
.B2(n_1209),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1216),
.A2(n_1207),
.B1(n_1209),
.B2(n_1204),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1213),
.Y(n_1222)
);

NAND4xp25_ASAP7_75t_L g1223 ( 
.A(n_1211),
.B(n_89),
.C(n_102),
.D(n_104),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1215),
.Y(n_1224)
);

NAND4xp25_ASAP7_75t_SL g1225 ( 
.A(n_1218),
.B(n_107),
.C(n_108),
.D(n_109),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_1220),
.A2(n_1219),
.B1(n_1212),
.B2(n_1217),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1222),
.A2(n_1210),
.B1(n_113),
.B2(n_117),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1224),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1221),
.A2(n_387),
.B1(n_118),
.B2(n_119),
.Y(n_1229)
);

OAI22x1_ASAP7_75t_L g1230 ( 
.A1(n_1228),
.A2(n_1225),
.B1(n_1223),
.B2(n_123),
.Y(n_1230)
);

OAI221xp5_ASAP7_75t_R g1231 ( 
.A1(n_1230),
.A2(n_1229),
.B1(n_1226),
.B2(n_1227),
.C(n_127),
.Y(n_1231)
);

OR2x6_ASAP7_75t_L g1232 ( 
.A(n_1231),
.B(n_387),
.Y(n_1232)
);

AOI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1232),
.A2(n_112),
.B1(n_120),
.B2(n_125),
.Y(n_1233)
);

AOI221xp5_ASAP7_75t_L g1234 ( 
.A1(n_1233),
.A2(n_387),
.B1(n_130),
.B2(n_132),
.C(n_136),
.Y(n_1234)
);

AOI211xp5_ASAP7_75t_L g1235 ( 
.A1(n_1234),
.A2(n_129),
.B(n_138),
.C(n_139),
.Y(n_1235)
);


endmodule