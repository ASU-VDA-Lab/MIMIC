module fake_jpeg_9430_n_145 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_26),
.Y(n_33)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_16),
.B1(n_14),
.B2(n_22),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_29),
.B1(n_39),
.B2(n_35),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_14),
.Y(n_37)
);

XNOR2x1_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_25),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_26),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_43),
.A2(n_42),
.B1(n_31),
.B2(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_49),
.B1(n_28),
.B2(n_35),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_25),
.C(n_23),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_26),
.B(n_20),
.C(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_51),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_12),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_25),
.C(n_23),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_42),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_37),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_62),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_28),
.B(n_13),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_13),
.B(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_64),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_67),
.B(n_69),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_68),
.A2(n_70),
.B1(n_18),
.B2(n_15),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_42),
.B1(n_31),
.B2(n_30),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_50),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_74),
.Y(n_86)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_64),
.A2(n_54),
.B1(n_51),
.B2(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_85),
.B1(n_17),
.B2(n_21),
.Y(n_93)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_44),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_12),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_21),
.B1(n_19),
.B2(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_63),
.B1(n_58),
.B2(n_30),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_19),
.C(n_9),
.Y(n_84)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_17),
.A3(n_68),
.B1(n_58),
.B2(n_59),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_61),
.C(n_57),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_57),
.B(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_19),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_97),
.Y(n_104)
);

OAI32xp33_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_79),
.A3(n_77),
.B1(n_83),
.B2(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_93),
.A2(n_77),
.B1(n_73),
.B2(n_81),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_96),
.B(n_94),
.Y(n_113)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_106),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_22),
.B(n_12),
.C(n_74),
.D(n_4),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_98),
.B(n_87),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_95),
.Y(n_115)
);

AO21x1_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_113),
.B(n_104),
.Y(n_120)
);

BUFx12f_ASAP7_75t_SL g111 ( 
.A(n_103),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_117),
.B(n_118),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_107),
.B(n_74),
.C(n_12),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_12),
.C(n_2),
.Y(n_124)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_107),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_100),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_111),
.A2(n_109),
.B1(n_105),
.B2(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_117),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_3),
.C(n_5),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_0),
.B(n_2),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_121),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_123),
.B(n_110),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_131),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_122),
.B(n_9),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_130),
.Y(n_136)
);

NOR3xp33_ASAP7_75t_SL g131 ( 
.A(n_120),
.B(n_117),
.C(n_10),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_134),
.B(n_6),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_127),
.B(n_3),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_3),
.C(n_5),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_137),
.A2(n_138),
.B(n_140),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_6),
.C(n_7),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_134),
.B(n_6),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_133),
.B(n_8),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_143),
.B(n_142),
.CI(n_8),
.CON(n_144),
.SN(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_139),
.Y(n_145)
);


endmodule