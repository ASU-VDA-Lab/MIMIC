module fake_aes_1395_n_1505 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1505);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1505;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_822;
wire n_706;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1270;
wire n_1474;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_1489;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_345;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1291;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1442;
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_186), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_168), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_198), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_42), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_79), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_194), .Y(n_340) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_252), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_309), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_333), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_300), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_263), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_249), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_118), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_184), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_0), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_72), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_193), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g352 ( .A(n_271), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_240), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_77), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_32), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_76), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_290), .Y(n_358) );
NOR2xp67_ASAP7_75t_L g359 ( .A(n_86), .B(n_304), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_294), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_135), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_215), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_72), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_306), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_292), .Y(n_365) );
BUFx5_ASAP7_75t_L g366 ( .A(n_317), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_282), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_124), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_245), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_13), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_307), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_89), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_108), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_310), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_11), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_196), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_8), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_202), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_233), .Y(n_380) );
CKINVDCx20_ASAP7_75t_R g381 ( .A(n_185), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_241), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_295), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_164), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_137), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_272), .Y(n_386) );
INVxp33_ASAP7_75t_SL g387 ( .A(n_70), .Y(n_387) );
CKINVDCx14_ASAP7_75t_R g388 ( .A(n_64), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_86), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_236), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_12), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_42), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_180), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_264), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_182), .Y(n_395) );
BUFx5_ASAP7_75t_L g396 ( .A(n_320), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_160), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_321), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_66), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_325), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_175), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_75), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_330), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_24), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_187), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_146), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_77), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_139), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_132), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_68), .Y(n_411) );
INVxp33_ASAP7_75t_SL g412 ( .A(n_289), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_178), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_281), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_254), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_80), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_291), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_85), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_270), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_229), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_268), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_159), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g423 ( .A(n_152), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_214), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_92), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
BUFx10_ASAP7_75t_L g427 ( .A(n_130), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_68), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_280), .Y(n_429) );
INVx1_ASAP7_75t_SL g430 ( .A(n_213), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_297), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_9), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_172), .B(n_326), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_90), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_31), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_24), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_16), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_299), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_3), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_209), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_71), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_127), .B(n_191), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_181), .Y(n_443) );
CKINVDCx16_ASAP7_75t_R g444 ( .A(n_27), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_157), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_259), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_207), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_173), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_155), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_276), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_98), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_158), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_296), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_176), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_85), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g456 ( .A(n_89), .Y(n_456) );
INVxp67_ASAP7_75t_SL g457 ( .A(n_232), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_5), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_278), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_239), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_312), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_141), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_273), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_243), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_150), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_65), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_228), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_274), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_43), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_14), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_217), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_4), .Y(n_472) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_54), .Y(n_473) );
CKINVDCx5p33_ASAP7_75t_R g474 ( .A(n_9), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_50), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_109), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_119), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_112), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_143), .Y(n_479) );
INVxp33_ASAP7_75t_SL g480 ( .A(n_0), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_122), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_199), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_177), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_286), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_46), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_50), .Y(n_486) );
BUFx3_ASAP7_75t_L g487 ( .A(n_246), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_165), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_20), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_163), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_303), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_174), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_115), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_219), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_190), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_222), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_46), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_78), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_43), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_113), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_31), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_45), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_197), .Y(n_503) );
BUFx3_ASAP7_75t_L g504 ( .A(n_94), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_63), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_262), .Y(n_506) );
BUFx2_ASAP7_75t_L g507 ( .A(n_48), .Y(n_507) );
BUFx3_ASAP7_75t_L g508 ( .A(n_195), .Y(n_508) );
CKINVDCx16_ASAP7_75t_R g509 ( .A(n_51), .Y(n_509) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_129), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_301), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_17), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_386), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_366), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_376), .B(n_1), .Y(n_515) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_374), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_425), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_366), .B(n_1), .Y(n_518) );
INVx5_ASAP7_75t_L g519 ( .A(n_374), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_388), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_520) );
BUFx2_ASAP7_75t_L g521 ( .A(n_388), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_422), .B(n_2), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_366), .Y(n_523) );
AND2x4_ASAP7_75t_L g524 ( .A(n_431), .B(n_5), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_366), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_440), .B(n_6), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_374), .Y(n_527) );
BUFx3_ASAP7_75t_L g528 ( .A(n_386), .Y(n_528) );
INVx3_ASAP7_75t_L g529 ( .A(n_427), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g530 ( .A(n_361), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_427), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_425), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_427), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_490), .B(n_6), .Y(n_534) );
INVx3_ASAP7_75t_L g535 ( .A(n_373), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_366), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_469), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_371), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_469), .B(n_7), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_373), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_366), .Y(n_541) );
INVx2_ASAP7_75t_L g542 ( .A(n_366), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_507), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_374), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_504), .B(n_7), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_396), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_343), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_338), .B(n_10), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_336), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_437), .B(n_10), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_349), .B(n_11), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_396), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g554 ( .A1(n_520), .A2(n_470), .B1(n_509), .B2(n_444), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_521), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_514), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_529), .B(n_380), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_529), .B(n_356), .Y(n_558) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_516), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_514), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_514), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_521), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_521), .Y(n_563) );
BUFx4f_ASAP7_75t_L g564 ( .A(n_546), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_529), .B(n_357), .Y(n_565) );
BUFx8_ASAP7_75t_SL g566 ( .A(n_530), .Y(n_566) );
INVx1_ASAP7_75t_SL g567 ( .A(n_544), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_514), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_523), .Y(n_569) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_546), .B(n_471), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_539), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_529), .B(n_339), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_529), .B(n_419), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_523), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_523), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_525), .Y(n_577) );
OAI22x1_ASAP7_75t_L g578 ( .A1(n_520), .A2(n_339), .B1(n_474), .B2(n_378), .Y(n_578) );
INVx5_ASAP7_75t_L g579 ( .A(n_535), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g580 ( .A1(n_544), .A2(n_505), .B1(n_497), .B2(n_473), .C(n_392), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_538), .A2(n_474), .B1(n_498), .B2(n_378), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_525), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_525), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_525), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_531), .B(n_363), .Y(n_585) );
INVxp67_ASAP7_75t_L g586 ( .A(n_515), .Y(n_586) );
INVxp67_ASAP7_75t_SL g587 ( .A(n_515), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_541), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_531), .B(n_498), .Y(n_589) );
INVx3_ASAP7_75t_L g590 ( .A(n_539), .Y(n_590) );
CKINVDCx8_ASAP7_75t_R g591 ( .A(n_524), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_541), .Y(n_592) );
INVx4_ASAP7_75t_L g593 ( .A(n_546), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_531), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_539), .Y(n_595) );
BUFx2_ASAP7_75t_L g596 ( .A(n_531), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_541), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_541), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_531), .Y(n_599) );
AND2x4_ASAP7_75t_L g600 ( .A(n_562), .B(n_533), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_571), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_587), .B(n_533), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_596), .B(n_573), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_558), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_572), .A2(n_539), .B1(n_546), .B2(n_550), .Y(n_605) );
INVx3_ASAP7_75t_L g606 ( .A(n_593), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_571), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_567), .B(n_551), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_581), .B(n_551), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_558), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_596), .B(n_533), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_589), .B(n_562), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_563), .B(n_533), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_563), .B(n_533), .Y(n_614) );
NOR3xp33_ASAP7_75t_SL g615 ( .A(n_554), .B(n_512), .C(n_391), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_558), .B(n_524), .Y(n_616) );
OR2x6_ASAP7_75t_L g617 ( .A(n_578), .B(n_551), .Y(n_617) );
BUFx4f_ASAP7_75t_L g618 ( .A(n_570), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_571), .Y(n_619) );
NOR2xp33_ASAP7_75t_R g620 ( .A(n_591), .B(n_341), .Y(n_620) );
NOR3xp33_ASAP7_75t_SL g621 ( .A(n_580), .B(n_512), .C(n_399), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_565), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_565), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_565), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_575), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_575), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_575), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_555), .B(n_524), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_564), .B(n_524), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_585), .B(n_524), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_585), .B(n_550), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_585), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_585), .B(n_522), .Y(n_634) );
BUFx12f_ASAP7_75t_L g635 ( .A(n_570), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_572), .Y(n_636) );
O2A1O1Ixp33_ASAP7_75t_L g637 ( .A1(n_586), .A2(n_534), .B(n_526), .C(n_522), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_593), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_557), .B(n_526), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_591), .A2(n_341), .B1(n_381), .B2(n_372), .Y(n_640) );
INVx5_ASAP7_75t_L g641 ( .A(n_593), .Y(n_641) );
OR2x6_ASAP7_75t_L g642 ( .A(n_578), .B(n_534), .Y(n_642) );
BUFx3_ASAP7_75t_L g643 ( .A(n_564), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_572), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_572), .A2(n_590), .B1(n_595), .B2(n_564), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_593), .Y(n_646) );
INVx2_ASAP7_75t_SL g647 ( .A(n_570), .Y(n_647) );
INVxp67_ASAP7_75t_L g648 ( .A(n_566), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_590), .A2(n_381), .B1(n_385), .B2(n_372), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_574), .B(n_549), .Y(n_650) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_590), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_590), .B(n_546), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_595), .Y(n_653) );
INVx8_ASAP7_75t_L g654 ( .A(n_595), .Y(n_654) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_595), .B(n_539), .Y(n_655) );
AND2x4_ASAP7_75t_L g656 ( .A(n_594), .B(n_599), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
AND2x6_ASAP7_75t_SL g658 ( .A(n_556), .B(n_549), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_556), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_561), .A2(n_548), .B1(n_553), .B2(n_542), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_561), .B(n_553), .Y(n_661) );
OR2x6_ASAP7_75t_L g662 ( .A(n_568), .B(n_552), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_588), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_579), .Y(n_664) );
BUFx6f_ASAP7_75t_L g665 ( .A(n_588), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_579), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_598), .B(n_552), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_598), .Y(n_668) );
INVx5_ASAP7_75t_L g669 ( .A(n_579), .Y(n_669) );
INVx5_ASAP7_75t_L g670 ( .A(n_579), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_568), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_569), .A2(n_548), .B1(n_553), .B2(n_542), .Y(n_672) );
INVx3_ASAP7_75t_L g673 ( .A(n_579), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_597), .B(n_350), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_569), .B(n_412), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_577), .B(n_553), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_577), .B(n_536), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_582), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_582), .B(n_412), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_592), .B(n_540), .Y(n_680) );
OAI21xp33_ASAP7_75t_SL g681 ( .A1(n_592), .A2(n_518), .B(n_540), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_579), .Y(n_682) );
AND2x4_ASAP7_75t_L g683 ( .A(n_597), .B(n_385), .Y(n_683) );
AND2x6_ASAP7_75t_SL g684 ( .A(n_560), .B(n_389), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_560), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_576), .Y(n_686) );
AND2x4_ASAP7_75t_L g687 ( .A(n_576), .B(n_401), .Y(n_687) );
INVxp67_ASAP7_75t_L g688 ( .A(n_583), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_583), .A2(n_480), .B1(n_387), .B2(n_532), .C(n_517), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_584), .B(n_513), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_584), .Y(n_691) );
OR2x6_ASAP7_75t_L g692 ( .A(n_648), .B(n_518), .Y(n_692) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_663), .Y(n_693) );
INVx2_ASAP7_75t_SL g694 ( .A(n_608), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_667), .B(n_387), .Y(n_695) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_663), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_683), .B(n_405), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_604), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g699 ( .A1(n_662), .A2(n_462), .B1(n_478), .B2(n_401), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_634), .B(n_480), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_610), .Y(n_701) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_617), .B(n_462), .Y(n_702) );
BUFx12f_ASAP7_75t_L g703 ( .A(n_684), .Y(n_703) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_662), .A2(n_492), .B1(n_478), .B2(n_365), .Y(n_704) );
AOI222xp33_ASAP7_75t_L g705 ( .A1(n_635), .A2(n_532), .B1(n_537), .B2(n_517), .C1(n_402), .C2(n_408), .Y(n_705) );
INVx3_ASAP7_75t_L g706 ( .A(n_646), .Y(n_706) );
INVx4_ASAP7_75t_L g707 ( .A(n_641), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_649), .B(n_456), .Y(n_708) );
NOR2x1_ASAP7_75t_SL g709 ( .A(n_662), .B(n_442), .Y(n_709) );
INVx2_ASAP7_75t_SL g710 ( .A(n_600), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_618), .A2(n_535), .B1(n_513), .B2(n_528), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_620), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_647), .A2(n_492), .B1(n_365), .B2(n_398), .Y(n_713) );
BUFx2_ASAP7_75t_L g714 ( .A(n_620), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_650), .B(n_535), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_652), .A2(n_547), .B(n_536), .Y(n_716) );
OAI22xp5_ASAP7_75t_SL g717 ( .A1(n_617), .A2(n_398), .B1(n_407), .B2(n_335), .Y(n_717) );
AND2x4_ASAP7_75t_L g718 ( .A(n_674), .B(n_411), .Y(n_718) );
INVxp67_ASAP7_75t_L g719 ( .A(n_640), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_687), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_622), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_650), .B(n_535), .Y(n_722) );
INVx3_ASAP7_75t_L g723 ( .A(n_646), .Y(n_723) );
INVx6_ASAP7_75t_L g724 ( .A(n_658), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_637), .A2(n_535), .B(n_547), .C(n_543), .Y(n_725) );
HB1xp67_ASAP7_75t_L g726 ( .A(n_687), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_630), .A2(n_547), .B(n_433), .Y(n_727) );
OR2x2_ASAP7_75t_L g728 ( .A(n_609), .B(n_537), .Y(n_728) );
INVx4_ASAP7_75t_L g729 ( .A(n_641), .Y(n_729) );
BUFx2_ASAP7_75t_L g730 ( .A(n_629), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_612), .B(n_416), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_639), .B(n_513), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_618), .B(n_418), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_668), .Y(n_734) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_641), .Y(n_735) );
INVx3_ASAP7_75t_L g736 ( .A(n_641), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_643), .B(n_428), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_643), .B(n_432), .Y(n_738) );
BUFx6f_ASAP7_75t_L g739 ( .A(n_665), .Y(n_739) );
OR2x2_ASAP7_75t_L g740 ( .A(n_617), .B(n_543), .Y(n_740) );
BUFx6f_ASAP7_75t_L g741 ( .A(n_665), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_642), .Y(n_742) );
BUFx2_ASAP7_75t_L g743 ( .A(n_686), .Y(n_743) );
OAI21x1_ASAP7_75t_L g744 ( .A1(n_661), .A2(n_360), .B(n_343), .Y(n_744) );
BUFx3_ASAP7_75t_L g745 ( .A(n_669), .Y(n_745) );
OAI22xp5_ASAP7_75t_L g746 ( .A1(n_668), .A2(n_407), .B1(n_410), .B2(n_335), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_600), .B(n_434), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_623), .Y(n_748) );
BUFx2_ASAP7_75t_L g749 ( .A(n_656), .Y(n_749) );
AND2x4_ASAP7_75t_L g750 ( .A(n_624), .B(n_435), .Y(n_750) );
O2A1O1Ixp5_ASAP7_75t_L g751 ( .A1(n_630), .A2(n_457), .B(n_400), .C(n_364), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_638), .Y(n_752) );
INVx3_ASAP7_75t_L g753 ( .A(n_606), .Y(n_753) );
OAI33xp33_ASAP7_75t_L g754 ( .A1(n_602), .A2(n_451), .A3(n_439), .B1(n_455), .B2(n_441), .B3(n_436), .Y(n_754) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_671), .A2(n_410), .B1(n_465), .B2(n_423), .Y(n_755) );
O2A1O1Ixp33_ASAP7_75t_L g756 ( .A1(n_655), .A2(n_466), .B(n_472), .C(n_458), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_642), .A2(n_528), .B1(n_513), .B2(n_475), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_671), .A2(n_423), .B1(n_477), .B2(n_465), .Y(n_758) );
INVx1_ASAP7_75t_SL g759 ( .A(n_613), .Y(n_759) );
NOR2xp67_ASAP7_75t_L g760 ( .A(n_681), .B(n_477), .Y(n_760) );
AO32x2_ASAP7_75t_L g761 ( .A1(n_642), .A2(n_548), .A3(n_528), .B1(n_359), .B2(n_396), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g762 ( .A1(n_616), .A2(n_631), .B(n_614), .Y(n_762) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_689), .A2(n_511), .B1(n_510), .B2(n_486), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_626), .B(n_485), .Y(n_764) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_633), .B(n_489), .Y(n_765) );
BUFx6f_ASAP7_75t_L g766 ( .A(n_665), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_632), .B(n_499), .Y(n_767) );
BUFx2_ASAP7_75t_L g768 ( .A(n_654), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_632), .B(n_501), .Y(n_769) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_665), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_636), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_603), .A2(n_340), .B(n_337), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g773 ( .A(n_675), .B(n_502), .Y(n_773) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_605), .A2(n_352), .B(n_346), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_675), .B(n_500), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_621), .B(n_548), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_606), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_644), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_651), .Y(n_779) );
INVxp67_ASAP7_75t_L g780 ( .A(n_679), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_601), .Y(n_781) );
INVx2_ASAP7_75t_SL g782 ( .A(n_654), .Y(n_782) );
O2A1O1Ixp33_ASAP7_75t_L g783 ( .A1(n_621), .A2(n_548), .B(n_344), .C(n_345), .Y(n_783) );
BUFx6f_ASAP7_75t_L g784 ( .A(n_654), .Y(n_784) );
AND2x4_ASAP7_75t_L g785 ( .A(n_645), .B(n_342), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_653), .A2(n_348), .B(n_347), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_651), .B(n_351), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_615), .B(n_355), .Y(n_788) );
CKINVDCx16_ASAP7_75t_R g789 ( .A(n_679), .Y(n_789) );
INVx4_ASAP7_75t_L g790 ( .A(n_669), .Y(n_790) );
INVx2_ASAP7_75t_L g791 ( .A(n_601), .Y(n_791) );
BUFx12f_ASAP7_75t_L g792 ( .A(n_669), .Y(n_792) );
OR2x2_ASAP7_75t_L g793 ( .A(n_611), .B(n_12), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_607), .Y(n_794) );
AOI21xp5_ASAP7_75t_L g795 ( .A1(n_690), .A2(n_354), .B(n_353), .Y(n_795) );
O2A1O1Ixp33_ASAP7_75t_L g796 ( .A1(n_659), .A2(n_358), .B(n_367), .C(n_362), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_680), .A2(n_369), .B(n_375), .C(n_368), .Y(n_797) );
BUFx2_ASAP7_75t_L g798 ( .A(n_688), .Y(n_798) );
INVx3_ASAP7_75t_L g799 ( .A(n_673), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_678), .Y(n_800) );
CKINVDCx11_ASAP7_75t_R g801 ( .A(n_664), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_680), .A2(n_355), .B1(n_379), .B2(n_377), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_607), .B(n_393), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_619), .A2(n_355), .B1(n_383), .B2(n_382), .Y(n_804) );
INVx3_ASAP7_75t_L g805 ( .A(n_673), .Y(n_805) );
OR2x2_ASAP7_75t_L g806 ( .A(n_619), .B(n_13), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_661), .A2(n_394), .B(n_390), .Y(n_807) );
CKINVDCx11_ASAP7_75t_R g808 ( .A(n_666), .Y(n_808) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_670), .Y(n_809) );
A2O1A1Ixp33_ASAP7_75t_L g810 ( .A1(n_660), .A2(n_397), .B(n_404), .C(n_395), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_625), .Y(n_811) );
OR2x6_ASAP7_75t_L g812 ( .A(n_615), .B(n_355), .Y(n_812) );
INVx4_ASAP7_75t_L g813 ( .A(n_670), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_625), .Y(n_814) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_670), .Y(n_815) );
AND2x2_ASAP7_75t_L g816 ( .A(n_627), .B(n_14), .Y(n_816) );
OR2x6_ASAP7_75t_L g817 ( .A(n_682), .B(n_406), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_627), .Y(n_818) );
AND2x4_ASAP7_75t_L g819 ( .A(n_682), .B(n_409), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_628), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_628), .B(n_420), .Y(n_821) );
BUFx4f_ASAP7_75t_L g822 ( .A(n_657), .Y(n_822) );
INVx4_ASAP7_75t_L g823 ( .A(n_657), .Y(n_823) );
BUFx3_ASAP7_75t_L g824 ( .A(n_685), .Y(n_824) );
A2O1A1Ixp33_ASAP7_75t_L g825 ( .A1(n_660), .A2(n_414), .B(n_415), .C(n_413), .Y(n_825) );
OAI21x1_ASAP7_75t_L g826 ( .A1(n_744), .A2(n_676), .B(n_677), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g827 ( .A(n_789), .B(n_685), .Y(n_827) );
INVx6_ASAP7_75t_L g828 ( .A(n_792), .Y(n_828) );
OA21x2_ASAP7_75t_L g829 ( .A1(n_725), .A2(n_364), .B(n_360), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_798), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_716), .A2(n_672), .B(n_691), .Y(n_831) );
OA21x2_ASAP7_75t_L g832 ( .A1(n_760), .A2(n_426), .B(n_384), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_694), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_719), .A2(n_672), .B1(n_421), .B2(n_445), .Y(n_834) );
AO31x2_ASAP7_75t_L g835 ( .A1(n_797), .A2(n_810), .A3(n_825), .B(n_709), .Y(n_835) );
OAI21x1_ASAP7_75t_L g836 ( .A1(n_762), .A2(n_426), .B(n_384), .Y(n_836) );
AND2x4_ASAP7_75t_L g837 ( .A(n_784), .B(n_438), .Y(n_837) );
INVx2_ASAP7_75t_L g838 ( .A(n_818), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_750), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_818), .Y(n_840) );
CKINVDCx11_ASAP7_75t_R g841 ( .A(n_801), .Y(n_841) );
INVx3_ASAP7_75t_L g842 ( .A(n_707), .Y(n_842) );
OAI21xp5_ASAP7_75t_L g843 ( .A1(n_780), .A2(n_448), .B(n_447), .Y(n_843) );
BUFx3_ASAP7_75t_L g844 ( .A(n_808), .Y(n_844) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_734), .A2(n_454), .B1(n_459), .B2(n_450), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_750), .Y(n_846) );
NOR2x1_ASAP7_75t_SL g847 ( .A(n_784), .B(n_403), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g848 ( .A1(n_734), .A2(n_461), .B1(n_463), .B2(n_460), .Y(n_848) );
AO21x2_ASAP7_75t_L g849 ( .A1(n_715), .A2(n_468), .B(n_467), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_727), .A2(n_449), .B(n_446), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_800), .B(n_476), .Y(n_851) );
A2O1A1Ixp33_ASAP7_75t_L g852 ( .A1(n_783), .A2(n_479), .B(n_482), .C(n_481), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_699), .B(n_370), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_695), .B(n_483), .Y(n_854) );
AOI21x1_ASAP7_75t_SL g855 ( .A1(n_776), .A2(n_396), .B(n_403), .Y(n_855) );
INVx6_ASAP7_75t_SL g856 ( .A(n_692), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_730), .B(n_484), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_703), .Y(n_858) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_712), .Y(n_859) );
OAI21x1_ASAP7_75t_SL g860 ( .A1(n_709), .A2(n_503), .B(n_453), .Y(n_860) );
AO31x2_ASAP7_75t_L g861 ( .A1(n_773), .A2(n_453), .A3(n_503), .B(n_491), .Y(n_861) );
OAI21x1_ASAP7_75t_L g862 ( .A1(n_800), .A2(n_493), .B(n_488), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_720), .Y(n_863) );
AO21x2_ASAP7_75t_L g864 ( .A1(n_722), .A2(n_495), .B(n_494), .Y(n_864) );
INVx2_ASAP7_75t_SL g865 ( .A(n_743), .Y(n_865) );
OR2x6_ASAP7_75t_L g866 ( .A(n_704), .B(n_496), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_726), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g868 ( .A1(n_708), .A2(n_424), .B1(n_429), .B2(n_452), .Y(n_868) );
INVx3_ASAP7_75t_L g869 ( .A(n_707), .Y(n_869) );
INVx4_ASAP7_75t_L g870 ( .A(n_784), .Y(n_870) );
OAI21xp5_ASAP7_75t_L g871 ( .A1(n_771), .A2(n_506), .B(n_430), .Y(n_871) );
OAI21x1_ASAP7_75t_L g872 ( .A1(n_771), .A2(n_396), .B(n_516), .Y(n_872) );
NAND3xp33_ASAP7_75t_L g873 ( .A(n_788), .B(n_527), .C(n_516), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_724), .A2(n_452), .B1(n_487), .B2(n_464), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_698), .B(n_396), .Y(n_875) );
OR2x6_ASAP7_75t_L g876 ( .A(n_768), .B(n_464), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_728), .B(n_15), .Y(n_877) );
INVx2_ASAP7_75t_SL g878 ( .A(n_817), .Y(n_878) );
CKINVDCx11_ASAP7_75t_R g879 ( .A(n_742), .Y(n_879) );
A2O1A1Ixp33_ASAP7_75t_L g880 ( .A1(n_756), .A2(n_508), .B(n_443), .C(n_417), .Y(n_880) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_778), .A2(n_508), .B(n_519), .Y(n_881) );
OR2x6_ASAP7_75t_L g882 ( .A(n_782), .B(n_16), .Y(n_882) );
INVx2_ASAP7_75t_L g883 ( .A(n_823), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_823), .Y(n_884) );
BUFx5_ASAP7_75t_L g885 ( .A(n_811), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_806), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_824), .Y(n_887) );
OAI21xp5_ASAP7_75t_L g888 ( .A1(n_778), .A2(n_519), .B(n_516), .Y(n_888) );
CKINVDCx20_ASAP7_75t_R g889 ( .A(n_717), .Y(n_889) );
INVx2_ASAP7_75t_L g890 ( .A(n_781), .Y(n_890) );
AND2x4_ASAP7_75t_L g891 ( .A(n_729), .B(n_17), .Y(n_891) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_785), .A2(n_822), .B1(n_793), .B2(n_817), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_697), .B(n_18), .Y(n_893) );
INVx1_ASAP7_75t_L g894 ( .A(n_718), .Y(n_894) );
AOI21xp33_ASAP7_75t_L g895 ( .A1(n_796), .A2(n_527), .B(n_516), .Y(n_895) );
NOR2x1_ASAP7_75t_R g896 ( .A(n_714), .B(n_519), .Y(n_896) );
AO21x2_ASAP7_75t_L g897 ( .A1(n_795), .A2(n_527), .B(n_516), .Y(n_897) );
OAI22xp5_ASAP7_75t_SL g898 ( .A1(n_812), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_718), .Y(n_899) );
BUFx2_ASAP7_75t_L g900 ( .A(n_749), .Y(n_900) );
OAI21x1_ASAP7_75t_L g901 ( .A1(n_791), .A2(n_527), .B(n_516), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_794), .Y(n_902) );
OAI21x1_ASAP7_75t_L g903 ( .A1(n_820), .A2(n_527), .B(n_516), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_754), .A2(n_527), .B1(n_545), .B2(n_519), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_701), .Y(n_905) );
INVxp67_ASAP7_75t_L g906 ( .A(n_746), .Y(n_906) );
OAI21x1_ASAP7_75t_L g907 ( .A1(n_814), .A2(n_711), .B(n_751), .Y(n_907) );
OA21x2_ASAP7_75t_L g908 ( .A1(n_757), .A2(n_545), .B(n_527), .Y(n_908) );
AO31x2_ASAP7_75t_L g909 ( .A1(n_769), .A2(n_527), .A3(n_545), .B(n_519), .Y(n_909) );
OAI21x1_ASAP7_75t_L g910 ( .A1(n_807), .A2(n_545), .B(n_559), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_759), .B(n_19), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_752), .Y(n_912) );
CKINVDCx5p33_ASAP7_75t_R g913 ( .A(n_692), .Y(n_913) );
OAI21x1_ASAP7_75t_L g914 ( .A1(n_799), .A2(n_545), .B(n_559), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_721), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_748), .Y(n_916) );
NAND3xp33_ASAP7_75t_L g917 ( .A(n_705), .B(n_545), .C(n_519), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_785), .A2(n_545), .B1(n_519), .B2(n_23), .Y(n_918) );
INVx6_ASAP7_75t_L g919 ( .A(n_735), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_816), .Y(n_920) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_822), .A2(n_519), .B1(n_545), .B2(n_23), .Y(n_921) );
INVx1_ASAP7_75t_L g922 ( .A(n_740), .Y(n_922) );
INVxp67_ASAP7_75t_SL g923 ( .A(n_693), .Y(n_923) );
AO21x2_ASAP7_75t_L g924 ( .A1(n_772), .A2(n_559), .B(n_100), .Y(n_924) );
CKINVDCx6p67_ASAP7_75t_R g925 ( .A(n_812), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_731), .A2(n_559), .B1(n_22), .B2(n_25), .C(n_26), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_787), .Y(n_927) );
O2A1O1Ixp33_ASAP7_75t_L g928 ( .A1(n_767), .A2(n_25), .B(n_21), .C(n_22), .Y(n_928) );
INVx4_ASAP7_75t_L g929 ( .A(n_735), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_787), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_779), .B(n_21), .Y(n_931) );
OA21x2_ASAP7_75t_L g932 ( .A1(n_732), .A2(n_559), .B(n_101), .Y(n_932) );
AOI21xp5_ASAP7_75t_L g933 ( .A1(n_803), .A2(n_559), .B(n_102), .Y(n_933) );
INVx3_ASAP7_75t_L g934 ( .A(n_729), .Y(n_934) );
INVx5_ASAP7_75t_L g935 ( .A(n_735), .Y(n_935) );
AOI21xp5_ASAP7_75t_L g936 ( .A1(n_821), .A2(n_103), .B(n_99), .Y(n_936) );
NAND2xp5_ASAP7_75t_SL g937 ( .A(n_693), .B(n_26), .Y(n_937) );
OA21x2_ASAP7_75t_L g938 ( .A1(n_786), .A2(n_105), .B(n_104), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_700), .A2(n_107), .B(n_106), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_739), .A2(n_111), .B(n_110), .Y(n_940) );
OAI21x1_ASAP7_75t_L g941 ( .A1(n_799), .A2(n_116), .B(n_114), .Y(n_941) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_713), .B(n_27), .Y(n_942) );
OAI21xp5_ASAP7_75t_L g943 ( .A1(n_733), .A2(n_28), .B(n_29), .Y(n_943) );
OAI21x1_ASAP7_75t_SL g944 ( .A1(n_790), .A2(n_28), .B(n_29), .Y(n_944) );
AOI21xp5_ASAP7_75t_L g945 ( .A1(n_739), .A2(n_120), .B(n_117), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_755), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_819), .Y(n_947) );
AO21x2_ASAP7_75t_L g948 ( .A1(n_761), .A2(n_123), .B(n_121), .Y(n_948) );
INVx1_ASAP7_75t_SL g949 ( .A(n_693), .Y(n_949) );
OAI21x1_ASAP7_75t_L g950 ( .A1(n_805), .A2(n_126), .B(n_125), .Y(n_950) );
OAI21x1_ASAP7_75t_L g951 ( .A1(n_805), .A2(n_131), .B(n_128), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_764), .B(n_30), .Y(n_952) );
OAI21x1_ASAP7_75t_L g953 ( .A1(n_706), .A2(n_134), .B(n_133), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_819), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g955 ( .A(n_702), .B(n_30), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_737), .Y(n_956) );
NAND2x1p5_ASAP7_75t_L g957 ( .A(n_696), .B(n_33), .Y(n_957) );
AOI21xp33_ASAP7_75t_L g958 ( .A1(n_775), .A2(n_33), .B(n_34), .Y(n_958) );
INVx8_ASAP7_75t_L g959 ( .A(n_809), .Y(n_959) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_696), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_738), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_747), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_765), .Y(n_963) );
NAND4xp25_ASAP7_75t_L g964 ( .A(n_763), .B(n_35), .C(n_36), .D(n_37), .Y(n_964) );
INVx2_ASAP7_75t_L g965 ( .A(n_706), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_710), .Y(n_966) );
BUFx4f_ASAP7_75t_L g967 ( .A(n_809), .Y(n_967) );
OAI21x1_ASAP7_75t_L g968 ( .A1(n_723), .A2(n_138), .B(n_136), .Y(n_968) );
AO21x2_ASAP7_75t_L g969 ( .A1(n_761), .A2(n_142), .B(n_140), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_723), .A2(n_145), .B(n_144), .Y(n_970) );
INVx3_ASAP7_75t_L g971 ( .A(n_790), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_777), .Y(n_972) );
NOR2xp33_ASAP7_75t_L g973 ( .A(n_758), .B(n_37), .Y(n_973) );
AO21x2_ASAP7_75t_L g974 ( .A1(n_761), .A2(n_148), .B(n_147), .Y(n_974) );
OAI21xp5_ASAP7_75t_L g975 ( .A1(n_802), .A2(n_38), .B(n_39), .Y(n_975) );
OAI21x1_ASAP7_75t_L g976 ( .A1(n_736), .A2(n_151), .B(n_149), .Y(n_976) );
NAND3xp33_ASAP7_75t_L g977 ( .A(n_804), .B(n_39), .C(n_40), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_774), .A2(n_40), .B1(n_41), .B2(n_44), .Y(n_978) );
OAI21xp5_ASAP7_75t_L g979 ( .A1(n_753), .A2(n_41), .B(n_44), .Y(n_979) );
AO21x2_ASAP7_75t_L g980 ( .A1(n_739), .A2(n_154), .B(n_153), .Y(n_980) );
INVxp67_ASAP7_75t_SL g981 ( .A(n_696), .Y(n_981) );
AND2x2_ASAP7_75t_L g982 ( .A(n_813), .B(n_45), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_753), .Y(n_983) );
OA21x2_ASAP7_75t_L g984 ( .A1(n_836), .A2(n_872), .B(n_850), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_866), .B(n_745), .Y(n_985) );
AOI21xp5_ASAP7_75t_L g986 ( .A1(n_933), .A2(n_766), .B(n_741), .Y(n_986) );
BUFx12f_ASAP7_75t_L g987 ( .A(n_841), .Y(n_987) );
OAI21x1_ASAP7_75t_L g988 ( .A1(n_914), .A2(n_736), .B(n_741), .Y(n_988) );
NAND2x1p5_ASAP7_75t_L g989 ( .A(n_935), .B(n_813), .Y(n_989) );
NAND2x1p5_ASAP7_75t_L g990 ( .A(n_935), .B(n_809), .Y(n_990) );
INVx4_ASAP7_75t_SL g991 ( .A(n_882), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g992 ( .A1(n_866), .A2(n_946), .B1(n_917), .B2(n_962), .Y(n_992) );
OAI22xp33_ASAP7_75t_L g993 ( .A1(n_882), .A2(n_815), .B1(n_770), .B2(n_766), .Y(n_993) );
AO21x2_ASAP7_75t_L g994 ( .A1(n_881), .A2(n_766), .B(n_741), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_892), .A2(n_770), .B1(n_815), .B2(n_49), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_882), .A2(n_770), .B1(n_48), .B2(n_49), .Y(n_996) );
AOI21xp5_ASAP7_75t_L g997 ( .A1(n_892), .A2(n_161), .B(n_156), .Y(n_997) );
BUFx6f_ASAP7_75t_L g998 ( .A(n_967), .Y(n_998) );
A2O1A1Ixp33_ASAP7_75t_L g999 ( .A1(n_963), .A2(n_47), .B(n_52), .C(n_53), .Y(n_999) );
INVxp67_ASAP7_75t_L g1000 ( .A(n_827), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g1001 ( .A1(n_898), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_918), .A2(n_55), .B1(n_56), .B2(n_57), .Y(n_1002) );
BUFx12f_ASAP7_75t_L g1003 ( .A(n_858), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1004 ( .A(n_877), .B(n_56), .Y(n_1004) );
OR2x6_ASAP7_75t_L g1005 ( .A(n_828), .B(n_57), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1006 ( .A(n_926), .B(n_928), .C(n_977), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_918), .A2(n_58), .B1(n_59), .B2(n_60), .Y(n_1007) );
OAI221xp5_ASAP7_75t_L g1008 ( .A1(n_853), .A2(n_58), .B1(n_59), .B2(n_60), .C(n_61), .Y(n_1008) );
OAI211xp5_ASAP7_75t_L g1009 ( .A1(n_964), .A2(n_61), .B(n_62), .C(n_63), .Y(n_1009) );
OAI21xp5_ASAP7_75t_L g1010 ( .A1(n_852), .A2(n_62), .B(n_64), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_942), .A2(n_65), .B1(n_66), .B2(n_67), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_906), .B(n_922), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_878), .B(n_67), .Y(n_1013) );
AO21x2_ASAP7_75t_L g1014 ( .A1(n_881), .A2(n_166), .B(n_162), .Y(n_1014) );
OAI221xp5_ASAP7_75t_L g1015 ( .A1(n_956), .A2(n_69), .B1(n_70), .B2(n_71), .C(n_73), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_830), .B(n_69), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_931), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_961), .B(n_73), .Y(n_1018) );
AOI21xp5_ASAP7_75t_L g1019 ( .A1(n_875), .A2(n_169), .B(n_167), .Y(n_1019) );
OAI221xp5_ASAP7_75t_L g1020 ( .A1(n_854), .A2(n_74), .B1(n_75), .B2(n_76), .C(n_78), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_931), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_875), .A2(n_226), .B(n_332), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_964), .A2(n_74), .B1(n_79), .B2(n_80), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1024 ( .A1(n_876), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_1024) );
AOI222xp33_ASAP7_75t_L g1025 ( .A1(n_894), .A2(n_899), .B1(n_889), .B2(n_898), .C1(n_973), .C2(n_905), .Y(n_1025) );
INVx1_ASAP7_75t_SL g1026 ( .A(n_935), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1027 ( .A1(n_856), .A2(n_82), .B1(n_83), .B2(n_84), .Y(n_1027) );
OAI22xp5_ASAP7_75t_L g1028 ( .A1(n_886), .A2(n_84), .B1(n_87), .B2(n_88), .Y(n_1028) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_843), .A2(n_955), .B1(n_871), .B2(n_839), .C(n_846), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_845), .A2(n_87), .B1(n_88), .B2(n_90), .C(n_91), .Y(n_1030) );
OA21x2_ASAP7_75t_L g1031 ( .A1(n_901), .A2(n_234), .B(n_331), .Y(n_1031) );
INVx1_ASAP7_75t_L g1032 ( .A(n_863), .Y(n_1032) );
O2A1O1Ixp33_ASAP7_75t_L g1033 ( .A1(n_880), .A2(n_91), .B(n_92), .C(n_93), .Y(n_1033) );
OA21x2_ASAP7_75t_L g1034 ( .A1(n_903), .A2(n_235), .B(n_328), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_856), .A2(n_93), .B1(n_94), .B2(n_95), .Y(n_1035) );
AOI21xp33_ASAP7_75t_L g1036 ( .A1(n_896), .A2(n_95), .B(n_96), .Y(n_1036) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_843), .B(n_96), .Y(n_1037) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_910), .A2(n_238), .B(n_327), .Y(n_1038) );
AOI21xp5_ASAP7_75t_L g1039 ( .A1(n_888), .A2(n_237), .B(n_324), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_893), .B(n_97), .Y(n_1040) );
OAI22xp33_ASAP7_75t_L g1041 ( .A1(n_876), .A2(n_97), .B1(n_98), .B2(n_170), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_915), .B(n_171), .Y(n_1042) );
INVxp67_ASAP7_75t_L g1043 ( .A(n_865), .Y(n_1043) );
OAI21xp33_ASAP7_75t_L g1044 ( .A1(n_952), .A2(n_179), .B(n_183), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g1045 ( .A1(n_913), .A2(n_188), .B1(n_189), .B2(n_192), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_867), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_838), .Y(n_1047) );
INVx1_ASAP7_75t_SL g1048 ( .A(n_949), .Y(n_1048) );
BUFx6f_ASAP7_75t_L g1049 ( .A(n_967), .Y(n_1049) );
OAI21xp5_ASAP7_75t_L g1050 ( .A1(n_831), .A2(n_200), .B(n_201), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g1051 ( .A1(n_876), .A2(n_203), .B1(n_204), .B2(n_205), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_916), .Y(n_1052) );
AOI211xp5_ASAP7_75t_L g1053 ( .A1(n_868), .A2(n_206), .B(n_208), .C(n_210), .Y(n_1053) );
CKINVDCx16_ASAP7_75t_R g1054 ( .A(n_844), .Y(n_1054) );
BUFx2_ASAP7_75t_L g1055 ( .A(n_870), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_891), .Y(n_1056) );
OAI211xp5_ASAP7_75t_L g1057 ( .A1(n_943), .A2(n_211), .B(n_212), .C(n_216), .Y(n_1057) );
NAND2xp5_ASAP7_75t_L g1058 ( .A(n_927), .B(n_323), .Y(n_1058) );
INVx1_ASAP7_75t_L g1059 ( .A(n_833), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_840), .Y(n_1060) );
OAI22xp5_ASAP7_75t_L g1061 ( .A1(n_920), .A2(n_218), .B1(n_220), .B2(n_221), .Y(n_1061) );
CKINVDCx11_ASAP7_75t_R g1062 ( .A(n_879), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_871), .B(n_223), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_911), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_851), .Y(n_1065) );
INVxp67_ASAP7_75t_L g1066 ( .A(n_900), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_930), .B(n_224), .Y(n_1067) );
INVx2_ASAP7_75t_L g1068 ( .A(n_890), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_837), .B(n_225), .Y(n_1069) );
OAI211xp5_ASAP7_75t_L g1070 ( .A1(n_943), .A2(n_227), .B(n_230), .C(n_231), .Y(n_1070) );
OR2x2_ASAP7_75t_L g1071 ( .A(n_857), .B(n_242), .Y(n_1071) );
AOI22xp5_ASAP7_75t_L g1072 ( .A1(n_947), .A2(n_244), .B1(n_247), .B2(n_248), .Y(n_1072) );
INVx2_ASAP7_75t_L g1073 ( .A(n_902), .Y(n_1073) );
AOI21xp5_ASAP7_75t_L g1074 ( .A1(n_888), .A2(n_250), .B(n_251), .Y(n_1074) );
OAI22xp5_ASAP7_75t_L g1075 ( .A1(n_851), .A2(n_253), .B1(n_255), .B2(n_256), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_925), .A2(n_257), .B1(n_258), .B2(n_260), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1077 ( .A(n_954), .B(n_261), .Y(n_1077) );
NAND3xp33_ASAP7_75t_L g1078 ( .A(n_977), .B(n_265), .C(n_266), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_912), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_834), .B(n_322), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_957), .Y(n_1081) );
AO21x2_ASAP7_75t_L g1082 ( .A1(n_948), .A2(n_267), .B(n_269), .Y(n_1082) );
INVx2_ASAP7_75t_L g1083 ( .A(n_957), .Y(n_1083) );
AO21x2_ASAP7_75t_L g1084 ( .A1(n_948), .A2(n_275), .B(n_277), .Y(n_1084) );
INVx2_ASAP7_75t_L g1085 ( .A(n_885), .Y(n_1085) );
INVx3_ASAP7_75t_L g1086 ( .A(n_959), .Y(n_1086) );
NAND2xp5_ASAP7_75t_L g1087 ( .A(n_845), .B(n_316), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_979), .Y(n_1088) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_848), .B(n_870), .Y(n_1089) );
CKINVDCx16_ASAP7_75t_R g1090 ( .A(n_929), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_885), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_848), .B(n_279), .Y(n_1092) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_828), .Y(n_1093) );
AND2x2_ASAP7_75t_L g1094 ( .A(n_982), .B(n_979), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1095 ( .A1(n_975), .A2(n_283), .B1(n_284), .B2(n_285), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_966), .B(n_287), .Y(n_1096) );
OAI22xp5_ASAP7_75t_L g1097 ( .A1(n_975), .A2(n_288), .B1(n_293), .B2(n_298), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g1098 ( .A1(n_921), .A2(n_302), .B1(n_305), .B2(n_308), .Y(n_1098) );
NOR3xp33_ASAP7_75t_L g1099 ( .A(n_958), .B(n_311), .C(n_313), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_932), .A2(n_314), .B(n_315), .Y(n_1100) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_921), .A2(n_960), .B1(n_978), .B2(n_934), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_972), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_944), .Y(n_1103) );
NOR2xp33_ASAP7_75t_L g1104 ( .A(n_859), .B(n_869), .Y(n_1104) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_958), .A2(n_895), .B1(n_860), .B2(n_887), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_959), .Y(n_1106) );
OA21x2_ASAP7_75t_L g1107 ( .A1(n_941), .A2(n_951), .B(n_950), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_874), .A2(n_884), .B1(n_883), .B2(n_934), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_861), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_861), .Y(n_1110) );
CKINVDCx20_ASAP7_75t_R g1111 ( .A(n_959), .Y(n_1111) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_929), .B(n_971), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g1113 ( .A(n_919), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_842), .A2(n_971), .B1(n_919), .B2(n_949), .Y(n_1114) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_849), .A2(n_864), .B1(n_937), .B2(n_885), .Y(n_1115) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_885), .Y(n_1116) );
INVx1_ASAP7_75t_SL g1117 ( .A(n_885), .Y(n_1117) );
OAI211xp5_ASAP7_75t_L g1118 ( .A1(n_904), .A2(n_939), .B(n_832), .C(n_983), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_862), .B(n_835), .Y(n_1119) );
A2O1A1Ixp33_ASAP7_75t_L g1120 ( .A1(n_907), .A2(n_936), .B(n_904), .C(n_873), .Y(n_1120) );
NAND2xp5_ASAP7_75t_L g1121 ( .A(n_835), .B(n_861), .Y(n_1121) );
BUFx2_ASAP7_75t_L g1122 ( .A(n_923), .Y(n_1122) );
INVx1_ASAP7_75t_L g1123 ( .A(n_965), .Y(n_1123) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_835), .B(n_981), .Y(n_1124) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_909), .B(n_829), .Y(n_1125) );
OR2x2_ASAP7_75t_L g1126 ( .A(n_1012), .B(n_829), .Y(n_1126) );
BUFx4f_ASAP7_75t_SL g1127 ( .A(n_987), .Y(n_1127) );
HB1xp67_ASAP7_75t_L g1128 ( .A(n_1090), .Y(n_1128) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_989), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1130 ( .A(n_991), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1131 ( .A(n_1025), .B(n_847), .Y(n_1131) );
INVxp67_ASAP7_75t_L g1132 ( .A(n_1005), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1047), .B(n_974), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1109), .Y(n_1134) );
BUFx2_ASAP7_75t_L g1135 ( .A(n_1117), .Y(n_1135) );
HB1xp67_ASAP7_75t_L g1136 ( .A(n_991), .Y(n_1136) );
AND2x2_ASAP7_75t_L g1137 ( .A(n_1060), .B(n_974), .Y(n_1137) );
INVx3_ASAP7_75t_L g1138 ( .A(n_1117), .Y(n_1138) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_1037), .B(n_1068), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1110), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1073), .B(n_969), .Y(n_1141) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1116), .B(n_969), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1143 ( .A(n_991), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1121), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1052), .Y(n_1145) );
INVx2_ASAP7_75t_L g1146 ( .A(n_988), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1147 ( .A(n_1065), .B(n_909), .Y(n_1147) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_1085), .B(n_976), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1079), .B(n_909), .Y(n_1149) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1125), .Y(n_1150) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1119), .Y(n_1151) );
HB1xp67_ASAP7_75t_L g1152 ( .A(n_1026), .Y(n_1152) );
HB1xp67_ASAP7_75t_L g1153 ( .A(n_1026), .Y(n_1153) );
OR2x6_ASAP7_75t_L g1154 ( .A(n_995), .B(n_970), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_1089), .B(n_908), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1000), .B(n_897), .Y(n_1156) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1124), .Y(n_1157) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_1055), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1017), .Y(n_1159) );
BUFx3_ASAP7_75t_L g1160 ( .A(n_989), .Y(n_1160) );
OAI22xp5_ASAP7_75t_L g1161 ( .A1(n_992), .A2(n_873), .B1(n_908), .B2(n_938), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1043), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1021), .Y(n_1163) );
OR2x2_ASAP7_75t_L g1164 ( .A(n_1094), .B(n_924), .Y(n_1164) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1103), .Y(n_1165) );
INVx2_ASAP7_75t_L g1166 ( .A(n_1031), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1167 ( .A(n_1032), .B(n_897), .Y(n_1167) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1056), .B(n_932), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1088), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1102), .Y(n_1170) );
INVx1_ASAP7_75t_L g1171 ( .A(n_1091), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1123), .Y(n_1172) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1034), .Y(n_1173) );
NAND2xp5_ASAP7_75t_L g1174 ( .A(n_1046), .B(n_826), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1092), .B(n_980), .Y(n_1175) );
HB1xp67_ASAP7_75t_L g1176 ( .A(n_1066), .Y(n_1176) );
INVx2_ASAP7_75t_L g1177 ( .A(n_1034), .Y(n_1177) );
INVx2_ASAP7_75t_L g1178 ( .A(n_984), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1081), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1083), .Y(n_1180) );
INVx1_ASAP7_75t_L g1181 ( .A(n_994), .Y(n_1181) );
BUFx2_ASAP7_75t_L g1182 ( .A(n_994), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1063), .B(n_980), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1082), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_985), .B(n_953), .Y(n_1185) );
HB1xp67_ASAP7_75t_L g1186 ( .A(n_1005), .Y(n_1186) );
INVx2_ASAP7_75t_L g1187 ( .A(n_984), .Y(n_1187) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_990), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1082), .Y(n_1189) );
INVxp67_ASAP7_75t_SL g1190 ( .A(n_995), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1112), .B(n_1064), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1084), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1004), .B(n_1040), .Y(n_1193) );
INVx1_ASAP7_75t_SL g1194 ( .A(n_1111), .Y(n_1194) );
NAND2xp5_ASAP7_75t_L g1195 ( .A(n_1059), .B(n_940), .Y(n_1195) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1084), .Y(n_1196) );
BUFx3_ASAP7_75t_L g1197 ( .A(n_990), .Y(n_1197) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1107), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1107), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1112), .B(n_968), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1001), .B(n_945), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1042), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1010), .B(n_855), .Y(n_1203) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_1122), .Y(n_1204) );
BUFx3_ASAP7_75t_L g1205 ( .A(n_998), .Y(n_1205) );
HB1xp67_ASAP7_75t_L g1206 ( .A(n_1005), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1028), .Y(n_1207) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1014), .Y(n_1208) );
AOI222xp33_ASAP7_75t_L g1209 ( .A1(n_1028), .A2(n_1030), .B1(n_1029), .B2(n_1023), .C1(n_1007), .C2(n_1002), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1010), .B(n_1069), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1016), .B(n_1048), .Y(n_1211) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1014), .Y(n_1212) );
INVx3_ASAP7_75t_L g1213 ( .A(n_998), .Y(n_1213) );
INVxp67_ASAP7_75t_L g1214 ( .A(n_1013), .Y(n_1214) );
BUFx3_ASAP7_75t_L g1215 ( .A(n_998), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1048), .B(n_999), .Y(n_1216) );
INVx3_ASAP7_75t_L g1217 ( .A(n_1049), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1108), .Y(n_1218) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1050), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1077), .B(n_1018), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1106), .B(n_1104), .Y(n_1221) );
OAI332xp33_ASAP7_75t_L g1222 ( .A1(n_1008), .A2(n_1054), .A3(n_1015), .B1(n_1024), .B2(n_1020), .B3(n_1041), .C1(n_996), .C2(n_1093), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1050), .Y(n_1223) );
AND2x4_ASAP7_75t_L g1224 ( .A(n_1120), .B(n_1113), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1108), .Y(n_1225) );
INVx2_ASAP7_75t_L g1226 ( .A(n_1078), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1009), .Y(n_1227) );
BUFx2_ASAP7_75t_L g1228 ( .A(n_993), .Y(n_1228) );
NOR2xp67_ASAP7_75t_L g1229 ( .A(n_1057), .B(n_1070), .Y(n_1229) );
AND2x2_ASAP7_75t_L g1230 ( .A(n_1011), .B(n_1053), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1053), .B(n_1096), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1058), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1086), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1086), .B(n_1105), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1067), .Y(n_1235) );
HB1xp67_ASAP7_75t_L g1236 ( .A(n_1049), .Y(n_1236) );
INVx2_ASAP7_75t_L g1237 ( .A(n_1078), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1087), .B(n_1115), .Y(n_1238) );
AOI21xp5_ASAP7_75t_L g1239 ( .A1(n_986), .A2(n_1118), .B(n_1100), .Y(n_1239) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1113), .Y(n_1240) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1113), .B(n_997), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1027), .B(n_1035), .Y(n_1242) );
BUFx3_ASAP7_75t_L g1243 ( .A(n_1114), .Y(n_1243) );
INVx4_ASAP7_75t_L g1244 ( .A(n_1129), .Y(n_1244) );
HB1xp67_ASAP7_75t_L g1245 ( .A(n_1204), .Y(n_1245) );
AOI22xp33_ASAP7_75t_L g1246 ( .A1(n_1230), .A2(n_1006), .B1(n_1101), .B2(n_1036), .Y(n_1246) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1145), .Y(n_1247) );
AND2x4_ASAP7_75t_L g1248 ( .A(n_1151), .B(n_1045), .Y(n_1248) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1159), .B(n_1006), .Y(n_1249) );
INVxp67_ASAP7_75t_SL g1250 ( .A(n_1204), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1151), .B(n_1099), .Y(n_1251) );
OAI221xp5_ASAP7_75t_L g1252 ( .A1(n_1131), .A2(n_1033), .B1(n_1071), .B2(n_1051), .C(n_1076), .Y(n_1252) );
INVx2_ASAP7_75t_L g1253 ( .A(n_1187), .Y(n_1253) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1187), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1158), .B(n_1075), .Y(n_1255) );
INVxp67_ASAP7_75t_SL g1256 ( .A(n_1135), .Y(n_1256) );
NOR2x1_ASAP7_75t_SL g1257 ( .A(n_1129), .B(n_1075), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1163), .B(n_1145), .Y(n_1258) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_1152), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1150), .B(n_1061), .Y(n_1260) );
INVx3_ASAP7_75t_L g1261 ( .A(n_1138), .Y(n_1261) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1170), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1263 ( .A(n_1153), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_1230), .A2(n_1097), .B1(n_1095), .B2(n_1098), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1150), .B(n_1061), .Y(n_1265) );
INVxp67_ASAP7_75t_SL g1266 ( .A(n_1135), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1170), .Y(n_1267) );
AND2x4_ASAP7_75t_L g1268 ( .A(n_1185), .B(n_1072), .Y(n_1268) );
AND2x4_ASAP7_75t_L g1269 ( .A(n_1185), .B(n_1039), .Y(n_1269) );
BUFx3_ASAP7_75t_L g1270 ( .A(n_1160), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1271 ( .A(n_1211), .B(n_1139), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1172), .Y(n_1272) );
AO21x2_ASAP7_75t_L g1273 ( .A1(n_1239), .A2(n_1038), .B(n_1044), .Y(n_1273) );
OAI221xp5_ASAP7_75t_L g1274 ( .A1(n_1132), .A2(n_1080), .B1(n_1019), .B2(n_1022), .C(n_1074), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1193), .B(n_1062), .Y(n_1275) );
AND2x4_ASAP7_75t_L g1276 ( .A(n_1134), .B(n_1003), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1128), .B(n_1172), .Y(n_1277) );
INVx4_ASAP7_75t_L g1278 ( .A(n_1160), .Y(n_1278) );
HB1xp67_ASAP7_75t_L g1279 ( .A(n_1191), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1147), .B(n_1149), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1149), .B(n_1134), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_1209), .A2(n_1242), .B1(n_1227), .B2(n_1207), .Y(n_1282) );
NAND2xp33_ASAP7_75t_L g1283 ( .A(n_1231), .B(n_1210), .Y(n_1283) );
INVx2_ASAP7_75t_L g1284 ( .A(n_1187), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1285 ( .A(n_1191), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1176), .B(n_1186), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1198), .Y(n_1287) );
BUFx3_ASAP7_75t_L g1288 ( .A(n_1188), .Y(n_1288) );
OR2x2_ASAP7_75t_L g1289 ( .A(n_1194), .B(n_1162), .Y(n_1289) );
AND2x4_ASAP7_75t_L g1290 ( .A(n_1140), .B(n_1224), .Y(n_1290) );
AO21x2_ASAP7_75t_L g1291 ( .A1(n_1184), .A2(n_1196), .B(n_1192), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1169), .B(n_1144), .Y(n_1292) );
AND2x4_ASAP7_75t_L g1293 ( .A(n_1224), .B(n_1234), .Y(n_1293) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1165), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1144), .B(n_1165), .Y(n_1295) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1198), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1179), .B(n_1180), .Y(n_1297) );
AOI322xp5_ASAP7_75t_L g1298 ( .A1(n_1206), .A2(n_1190), .A3(n_1231), .B1(n_1130), .B2(n_1136), .C1(n_1143), .C2(n_1214), .Y(n_1298) );
AND2x4_ASAP7_75t_SL g1299 ( .A(n_1233), .B(n_1236), .Y(n_1299) );
INVx2_ASAP7_75t_SL g1300 ( .A(n_1188), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1157), .B(n_1218), .Y(n_1301) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1174), .Y(n_1302) );
INVx2_ASAP7_75t_L g1303 ( .A(n_1199), .Y(n_1303) );
INVx2_ASAP7_75t_L g1304 ( .A(n_1199), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1167), .Y(n_1305) );
BUFx6f_ASAP7_75t_L g1306 ( .A(n_1188), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1171), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1218), .B(n_1133), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1171), .Y(n_1309) );
AND2x4_ASAP7_75t_L g1310 ( .A(n_1224), .B(n_1200), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1311 ( .A1(n_1220), .A2(n_1201), .B1(n_1228), .B2(n_1238), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1156), .Y(n_1312) );
HB1xp67_ASAP7_75t_L g1313 ( .A(n_1197), .Y(n_1313) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1222), .B(n_1202), .Y(n_1314) );
AND2x2_ASAP7_75t_L g1315 ( .A(n_1137), .B(n_1175), .Y(n_1315) );
BUFx2_ASAP7_75t_L g1316 ( .A(n_1197), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1126), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1175), .B(n_1141), .Y(n_1318) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1141), .B(n_1238), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1126), .B(n_1155), .Y(n_1320) );
OR2x2_ASAP7_75t_L g1321 ( .A(n_1155), .B(n_1221), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1322 ( .A1(n_1202), .A2(n_1201), .B1(n_1216), .B2(n_1195), .C(n_1203), .Y(n_1322) );
AND2x4_ASAP7_75t_L g1323 ( .A(n_1224), .B(n_1200), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1247), .Y(n_1324) );
OAI21x1_ASAP7_75t_L g1325 ( .A1(n_1253), .A2(n_1166), .B(n_1173), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1282), .B(n_1225), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1327 ( .A1(n_1283), .A2(n_1203), .B1(n_1243), .B2(n_1216), .Y(n_1327) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1253), .Y(n_1328) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1262), .Y(n_1329) );
NAND2xp5_ASAP7_75t_SL g1330 ( .A(n_1244), .B(n_1243), .Y(n_1330) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1280), .B(n_1164), .Y(n_1331) );
OAI221xp5_ASAP7_75t_L g1332 ( .A1(n_1314), .A2(n_1154), .B1(n_1235), .B2(n_1232), .C(n_1229), .Y(n_1332) );
NOR2x1_ASAP7_75t_L g1333 ( .A(n_1244), .B(n_1154), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1334 ( .A(n_1282), .B(n_1225), .Y(n_1334) );
HB1xp67_ASAP7_75t_L g1335 ( .A(n_1245), .Y(n_1335) );
HB1xp67_ASAP7_75t_L g1336 ( .A(n_1259), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1267), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1280), .B(n_1181), .Y(n_1338) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1315), .B(n_1181), .Y(n_1339) );
INVx2_ASAP7_75t_SL g1340 ( .A(n_1299), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1315), .B(n_1164), .Y(n_1341) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1271), .B(n_1232), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1279), .B(n_1240), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1318), .B(n_1182), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1318), .B(n_1182), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1319), .B(n_1142), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1285), .B(n_1240), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1272), .Y(n_1348) );
OR2x2_ASAP7_75t_SL g1349 ( .A(n_1289), .B(n_1127), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1277), .Y(n_1350) );
HB1xp67_ASAP7_75t_L g1351 ( .A(n_1263), .Y(n_1351) );
OR2x2_ASAP7_75t_L g1352 ( .A(n_1320), .B(n_1168), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1319), .B(n_1142), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1321), .B(n_1168), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1258), .Y(n_1355) );
INVx2_ASAP7_75t_L g1356 ( .A(n_1254), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1281), .B(n_1178), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1286), .Y(n_1358) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1281), .B(n_1183), .Y(n_1359) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1294), .Y(n_1360) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1254), .Y(n_1361) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1284), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1308), .B(n_1183), .Y(n_1363) );
INVx1_ASAP7_75t_SL g1364 ( .A(n_1275), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1308), .B(n_1189), .Y(n_1365) );
NOR2x1_ASAP7_75t_L g1366 ( .A(n_1244), .B(n_1154), .Y(n_1366) );
AND2x4_ASAP7_75t_L g1367 ( .A(n_1310), .B(n_1138), .Y(n_1367) );
NAND3xp33_ASAP7_75t_L g1368 ( .A(n_1246), .B(n_1154), .C(n_1161), .Y(n_1368) );
INVx2_ASAP7_75t_SL g1369 ( .A(n_1278), .Y(n_1369) );
OR2x2_ASAP7_75t_L g1370 ( .A(n_1250), .B(n_1138), .Y(n_1370) );
AO21x2_ASAP7_75t_L g1371 ( .A1(n_1273), .A2(n_1177), .B(n_1173), .Y(n_1371) );
NOR3xp33_ASAP7_75t_SL g1372 ( .A(n_1252), .B(n_1205), .C(n_1215), .Y(n_1372) );
INVx1_ASAP7_75t_SL g1373 ( .A(n_1276), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1307), .Y(n_1374) );
AOI221xp5_ASAP7_75t_L g1375 ( .A1(n_1311), .A2(n_1213), .B1(n_1217), .B2(n_1205), .C(n_1215), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1295), .B(n_1213), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1309), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1378 ( .A(n_1295), .B(n_1213), .Y(n_1378) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1284), .Y(n_1379) );
BUFx2_ASAP7_75t_L g1380 ( .A(n_1270), .Y(n_1380) );
INVx1_ASAP7_75t_SL g1381 ( .A(n_1276), .Y(n_1381) );
OR2x2_ASAP7_75t_L g1382 ( .A(n_1331), .B(n_1312), .Y(n_1382) );
INVx2_ASAP7_75t_L g1383 ( .A(n_1328), .Y(n_1383) );
OR2x6_ASAP7_75t_L g1384 ( .A(n_1333), .B(n_1290), .Y(n_1384) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_1340), .Y(n_1385) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1336), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1363), .B(n_1293), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1351), .Y(n_1388) );
NAND2x1p5_ASAP7_75t_L g1389 ( .A(n_1369), .B(n_1270), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1324), .Y(n_1390) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1329), .Y(n_1391) );
NAND2x1p5_ASAP7_75t_L g1392 ( .A(n_1369), .B(n_1288), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1359), .B(n_1293), .Y(n_1393) );
INVx1_ASAP7_75t_SL g1394 ( .A(n_1340), .Y(n_1394) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1331), .B(n_1305), .Y(n_1395) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1337), .Y(n_1396) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1358), .B(n_1292), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1350), .B(n_1292), .Y(n_1398) );
NAND4xp25_ASAP7_75t_SL g1399 ( .A(n_1373), .B(n_1381), .C(n_1349), .D(n_1327), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1359), .B(n_1293), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1341), .B(n_1323), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_1326), .A2(n_1322), .B1(n_1248), .B2(n_1276), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1341), .B(n_1323), .Y(n_1403) );
INVxp67_ASAP7_75t_L g1404 ( .A(n_1335), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1363), .B(n_1323), .Y(n_1405) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1338), .B(n_1310), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1348), .Y(n_1407) );
OR2x2_ASAP7_75t_L g1408 ( .A(n_1338), .B(n_1317), .Y(n_1408) );
OR2x2_ASAP7_75t_L g1409 ( .A(n_1339), .B(n_1297), .Y(n_1409) );
OR2x6_ASAP7_75t_L g1410 ( .A(n_1366), .B(n_1290), .Y(n_1410) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1360), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1412 ( .A(n_1344), .B(n_1310), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1413 ( .A(n_1364), .B(n_1249), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1355), .B(n_1301), .Y(n_1414) );
INVx3_ASAP7_75t_L g1415 ( .A(n_1367), .Y(n_1415) );
INVx2_ASAP7_75t_L g1416 ( .A(n_1328), .Y(n_1416) );
AND2x4_ASAP7_75t_L g1417 ( .A(n_1367), .B(n_1290), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1344), .B(n_1266), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1374), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1377), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1342), .B(n_1298), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1422 ( .A(n_1345), .B(n_1256), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g1423 ( .A(n_1356), .Y(n_1423) );
OR2x2_ASAP7_75t_L g1424 ( .A(n_1354), .B(n_1345), .Y(n_1424) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_1399), .A2(n_1368), .B1(n_1332), .B2(n_1334), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1390), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1421), .B(n_1365), .Y(n_1427) );
OR2x2_ASAP7_75t_L g1428 ( .A(n_1424), .B(n_1352), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1386), .B(n_1365), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1388), .B(n_1357), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1391), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1396), .Y(n_1432) );
NAND2xp5_ASAP7_75t_SL g1433 ( .A(n_1385), .B(n_1380), .Y(n_1433) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1407), .Y(n_1434) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_1402), .A2(n_1372), .B1(n_1248), .B2(n_1375), .Y(n_1435) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1411), .Y(n_1436) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1419), .Y(n_1437) );
OAI22xp33_ASAP7_75t_L g1438 ( .A1(n_1385), .A2(n_1255), .B1(n_1330), .B2(n_1316), .Y(n_1438) );
NAND3xp33_ASAP7_75t_SL g1439 ( .A(n_1394), .B(n_1264), .C(n_1313), .Y(n_1439) );
OAI22xp5_ASAP7_75t_L g1440 ( .A1(n_1402), .A2(n_1264), .B1(n_1300), .B2(n_1376), .Y(n_1440) );
NOR2xp33_ASAP7_75t_L g1441 ( .A(n_1413), .B(n_1378), .Y(n_1441) );
OAI22x1_ASAP7_75t_L g1442 ( .A1(n_1404), .A2(n_1367), .B1(n_1346), .B2(n_1353), .Y(n_1442) );
OA21x2_ASAP7_75t_L g1443 ( .A1(n_1423), .A2(n_1325), .B(n_1379), .Y(n_1443) );
INVx2_ASAP7_75t_L g1444 ( .A(n_1383), .Y(n_1444) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1409), .B(n_1352), .Y(n_1445) );
O2A1O1Ixp33_ASAP7_75t_SL g1446 ( .A1(n_1397), .A2(n_1347), .B(n_1343), .C(n_1370), .Y(n_1446) );
AOI221x1_ASAP7_75t_L g1447 ( .A1(n_1413), .A2(n_1306), .B1(n_1302), .B2(n_1251), .C(n_1241), .Y(n_1447) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1414), .B(n_1353), .Y(n_1448) );
O2A1O1Ixp33_ASAP7_75t_L g1449 ( .A1(n_1389), .A2(n_1274), .B(n_1251), .C(n_1217), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1426), .Y(n_1450) );
OAI221xp5_ASAP7_75t_L g1451 ( .A1(n_1425), .A2(n_1382), .B1(n_1395), .B2(n_1398), .C(n_1389), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1442), .B(n_1387), .Y(n_1452) );
INVxp33_ASAP7_75t_L g1453 ( .A(n_1433), .Y(n_1453) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1431), .Y(n_1454) );
NOR2x1_ASAP7_75t_L g1455 ( .A(n_1439), .B(n_1410), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1456 ( .A(n_1445), .B(n_1408), .Y(n_1456) );
INVx2_ASAP7_75t_SL g1457 ( .A(n_1444), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1432), .Y(n_1458) );
INVx2_ASAP7_75t_SL g1459 ( .A(n_1428), .Y(n_1459) );
OAI322xp33_ASAP7_75t_SL g1460 ( .A1(n_1427), .A2(n_1420), .A3(n_1416), .B1(n_1383), .B2(n_1379), .C1(n_1362), .C2(n_1361), .Y(n_1460) );
AOI221xp5_ASAP7_75t_L g1461 ( .A1(n_1440), .A2(n_1405), .B1(n_1400), .B2(n_1393), .C(n_1406), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1441), .B(n_1405), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1463 ( .A(n_1446), .B(n_1422), .Y(n_1463) );
AOI211xp5_ASAP7_75t_L g1464 ( .A1(n_1438), .A2(n_1417), .B(n_1415), .C(n_1418), .Y(n_1464) );
OAI211xp5_ASAP7_75t_L g1465 ( .A1(n_1435), .A2(n_1415), .B(n_1412), .C(n_1401), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1434), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1436), .Y(n_1467) );
XNOR2x2_ASAP7_75t_L g1468 ( .A(n_1439), .B(n_1403), .Y(n_1468) );
NOR2xp33_ASAP7_75t_L g1469 ( .A(n_1453), .B(n_1437), .Y(n_1469) );
AOI22xp5_ASAP7_75t_L g1470 ( .A1(n_1465), .A2(n_1429), .B1(n_1430), .B2(n_1448), .Y(n_1470) );
INVx2_ASAP7_75t_L g1471 ( .A(n_1457), .Y(n_1471) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1450), .Y(n_1472) );
AOI21xp5_ASAP7_75t_L g1473 ( .A1(n_1460), .A2(n_1449), .B(n_1447), .Y(n_1473) );
AOI211xp5_ASAP7_75t_L g1474 ( .A1(n_1453), .A2(n_1449), .B(n_1417), .C(n_1268), .Y(n_1474) );
AOI21xp5_ASAP7_75t_L g1475 ( .A1(n_1455), .A2(n_1392), .B(n_1384), .Y(n_1475) );
AOI22xp5_ASAP7_75t_L g1476 ( .A1(n_1451), .A2(n_1417), .B1(n_1384), .B2(n_1410), .Y(n_1476) );
INVxp67_ASAP7_75t_L g1477 ( .A(n_1463), .Y(n_1477) );
INVxp33_ASAP7_75t_L g1478 ( .A(n_1452), .Y(n_1478) );
AOI21xp5_ASAP7_75t_L g1479 ( .A1(n_1464), .A2(n_1257), .B(n_1443), .Y(n_1479) );
OAI211xp5_ASAP7_75t_SL g1480 ( .A1(n_1477), .A2(n_1461), .B(n_1468), .C(n_1466), .Y(n_1480) );
OAI211xp5_ASAP7_75t_SL g1481 ( .A1(n_1474), .A2(n_1473), .B(n_1476), .C(n_1475), .Y(n_1481) );
NAND3xp33_ASAP7_75t_L g1482 ( .A(n_1479), .B(n_1458), .C(n_1454), .Y(n_1482) );
OAI211xp5_ASAP7_75t_SL g1483 ( .A1(n_1470), .A2(n_1468), .B(n_1467), .C(n_1459), .Y(n_1483) );
AOI211xp5_ASAP7_75t_L g1484 ( .A1(n_1478), .A2(n_1452), .B(n_1462), .C(n_1456), .Y(n_1484) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_1469), .A2(n_1443), .B1(n_1217), .B2(n_1306), .C(n_1261), .Y(n_1485) );
AOI221xp5_ASAP7_75t_L g1486 ( .A1(n_1472), .A2(n_1269), .B1(n_1265), .B2(n_1260), .C(n_1361), .Y(n_1486) );
NOR2x1_ASAP7_75t_L g1487 ( .A(n_1483), .B(n_1471), .Y(n_1487) );
NOR2xp67_ASAP7_75t_L g1488 ( .A(n_1482), .B(n_1356), .Y(n_1488) );
OAI211xp5_ASAP7_75t_SL g1489 ( .A1(n_1484), .A2(n_1261), .B(n_1237), .C(n_1226), .Y(n_1489) );
NOR2xp33_ASAP7_75t_L g1490 ( .A(n_1481), .B(n_1261), .Y(n_1490) );
NOR2xp33_ASAP7_75t_L g1491 ( .A(n_1480), .B(n_1362), .Y(n_1491) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1485), .Y(n_1492) );
INVxp67_ASAP7_75t_SL g1493 ( .A(n_1492), .Y(n_1493) );
OAI222xp33_ASAP7_75t_L g1494 ( .A1(n_1487), .A2(n_1486), .B1(n_1241), .B2(n_1304), .C1(n_1303), .C2(n_1296), .Y(n_1494) );
NAND3xp33_ASAP7_75t_SL g1495 ( .A(n_1490), .B(n_1208), .C(n_1212), .Y(n_1495) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1491), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1493), .Y(n_1497) );
OR2x2_ASAP7_75t_SL g1498 ( .A(n_1496), .B(n_1489), .Y(n_1498) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1495), .Y(n_1499) );
AO22x2_ASAP7_75t_L g1500 ( .A1(n_1497), .A2(n_1495), .B1(n_1494), .B2(n_1488), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g1501 ( .A1(n_1499), .A2(n_1291), .B1(n_1371), .B2(n_1273), .Y(n_1501) );
INVx2_ASAP7_75t_L g1502 ( .A(n_1500), .Y(n_1502) );
AOI21xp5_ASAP7_75t_L g1503 ( .A1(n_1502), .A2(n_1501), .B(n_1498), .Y(n_1503) );
AOI22x1_ASAP7_75t_L g1504 ( .A1(n_1503), .A2(n_1148), .B1(n_1219), .B2(n_1223), .Y(n_1504) );
AOI222xp33_ASAP7_75t_L g1505 ( .A1(n_1504), .A2(n_1146), .B1(n_1296), .B2(n_1287), .C1(n_1303), .C2(n_1304), .Y(n_1505) );
endmodule